-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jan 3 2025 14:09:01

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MAIN" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MAIN
entity MAIN is
port (
    rgb_g : out std_logic;
    T01 : out std_logic;
    start_stop : in std_logic;
    s2_phy : out std_logic;
    T23 : out std_logic;
    s3_phy : out std_logic;
    il_min_comp2 : in std_logic;
    il_max_comp1 : in std_logic;
    clock_output : out std_logic;
    s1_phy : out std_logic;
    reset : in std_logic;
    il_min_comp1 : in std_logic;
    delay_tr_input : in std_logic;
    T45 : out std_logic;
    T12 : out std_logic;
    s4_phy : out std_logic;
    rgb_r : out std_logic;
    rgb_b : out std_logic;
    pwm_output : out std_logic;
    il_max_comp2 : in std_logic;
    delay_hc_input : in std_logic);
end MAIN;

-- Architecture of MAIN
-- View name is \INTERFACE\
architecture \INTERFACE\ of MAIN is

signal \N__50564\ : std_logic;
signal \N__50563\ : std_logic;
signal \N__50562\ : std_logic;
signal \N__50553\ : std_logic;
signal \N__50552\ : std_logic;
signal \N__50551\ : std_logic;
signal \N__50544\ : std_logic;
signal \N__50543\ : std_logic;
signal \N__50542\ : std_logic;
signal \N__50535\ : std_logic;
signal \N__50534\ : std_logic;
signal \N__50533\ : std_logic;
signal \N__50526\ : std_logic;
signal \N__50525\ : std_logic;
signal \N__50524\ : std_logic;
signal \N__50517\ : std_logic;
signal \N__50516\ : std_logic;
signal \N__50515\ : std_logic;
signal \N__50508\ : std_logic;
signal \N__50507\ : std_logic;
signal \N__50506\ : std_logic;
signal \N__50499\ : std_logic;
signal \N__50498\ : std_logic;
signal \N__50497\ : std_logic;
signal \N__50490\ : std_logic;
signal \N__50489\ : std_logic;
signal \N__50488\ : std_logic;
signal \N__50481\ : std_logic;
signal \N__50480\ : std_logic;
signal \N__50479\ : std_logic;
signal \N__50472\ : std_logic;
signal \N__50471\ : std_logic;
signal \N__50470\ : std_logic;
signal \N__50463\ : std_logic;
signal \N__50462\ : std_logic;
signal \N__50461\ : std_logic;
signal \N__50454\ : std_logic;
signal \N__50453\ : std_logic;
signal \N__50452\ : std_logic;
signal \N__50445\ : std_logic;
signal \N__50444\ : std_logic;
signal \N__50443\ : std_logic;
signal \N__50436\ : std_logic;
signal \N__50435\ : std_logic;
signal \N__50434\ : std_logic;
signal \N__50427\ : std_logic;
signal \N__50426\ : std_logic;
signal \N__50425\ : std_logic;
signal \N__50418\ : std_logic;
signal \N__50417\ : std_logic;
signal \N__50416\ : std_logic;
signal \N__50409\ : std_logic;
signal \N__50408\ : std_logic;
signal \N__50407\ : std_logic;
signal \N__50390\ : std_logic;
signal \N__50387\ : std_logic;
signal \N__50386\ : std_logic;
signal \N__50385\ : std_logic;
signal \N__50382\ : std_logic;
signal \N__50379\ : std_logic;
signal \N__50376\ : std_logic;
signal \N__50371\ : std_logic;
signal \N__50366\ : std_logic;
signal \N__50363\ : std_logic;
signal \N__50362\ : std_logic;
signal \N__50359\ : std_logic;
signal \N__50356\ : std_logic;
signal \N__50355\ : std_logic;
signal \N__50354\ : std_logic;
signal \N__50349\ : std_logic;
signal \N__50346\ : std_logic;
signal \N__50343\ : std_logic;
signal \N__50338\ : std_logic;
signal \N__50335\ : std_logic;
signal \N__50332\ : std_logic;
signal \N__50329\ : std_logic;
signal \N__50324\ : std_logic;
signal \N__50321\ : std_logic;
signal \N__50320\ : std_logic;
signal \N__50319\ : std_logic;
signal \N__50318\ : std_logic;
signal \N__50317\ : std_logic;
signal \N__50316\ : std_logic;
signal \N__50315\ : std_logic;
signal \N__50314\ : std_logic;
signal \N__50313\ : std_logic;
signal \N__50312\ : std_logic;
signal \N__50311\ : std_logic;
signal \N__50310\ : std_logic;
signal \N__50309\ : std_logic;
signal \N__50308\ : std_logic;
signal \N__50307\ : std_logic;
signal \N__50306\ : std_logic;
signal \N__50305\ : std_logic;
signal \N__50304\ : std_logic;
signal \N__50303\ : std_logic;
signal \N__50302\ : std_logic;
signal \N__50301\ : std_logic;
signal \N__50300\ : std_logic;
signal \N__50299\ : std_logic;
signal \N__50298\ : std_logic;
signal \N__50297\ : std_logic;
signal \N__50296\ : std_logic;
signal \N__50295\ : std_logic;
signal \N__50294\ : std_logic;
signal \N__50293\ : std_logic;
signal \N__50292\ : std_logic;
signal \N__50291\ : std_logic;
signal \N__50290\ : std_logic;
signal \N__50289\ : std_logic;
signal \N__50288\ : std_logic;
signal \N__50287\ : std_logic;
signal \N__50286\ : std_logic;
signal \N__50285\ : std_logic;
signal \N__50284\ : std_logic;
signal \N__50283\ : std_logic;
signal \N__50282\ : std_logic;
signal \N__50281\ : std_logic;
signal \N__50280\ : std_logic;
signal \N__50279\ : std_logic;
signal \N__50278\ : std_logic;
signal \N__50277\ : std_logic;
signal \N__50276\ : std_logic;
signal \N__50275\ : std_logic;
signal \N__50274\ : std_logic;
signal \N__50273\ : std_logic;
signal \N__50272\ : std_logic;
signal \N__50271\ : std_logic;
signal \N__50270\ : std_logic;
signal \N__50269\ : std_logic;
signal \N__50268\ : std_logic;
signal \N__50267\ : std_logic;
signal \N__50266\ : std_logic;
signal \N__50265\ : std_logic;
signal \N__50264\ : std_logic;
signal \N__50263\ : std_logic;
signal \N__50262\ : std_logic;
signal \N__50261\ : std_logic;
signal \N__50260\ : std_logic;
signal \N__50259\ : std_logic;
signal \N__50258\ : std_logic;
signal \N__50257\ : std_logic;
signal \N__50256\ : std_logic;
signal \N__50255\ : std_logic;
signal \N__50254\ : std_logic;
signal \N__50253\ : std_logic;
signal \N__50252\ : std_logic;
signal \N__50251\ : std_logic;
signal \N__50250\ : std_logic;
signal \N__50249\ : std_logic;
signal \N__50248\ : std_logic;
signal \N__50247\ : std_logic;
signal \N__50246\ : std_logic;
signal \N__50245\ : std_logic;
signal \N__50244\ : std_logic;
signal \N__50243\ : std_logic;
signal \N__50242\ : std_logic;
signal \N__50241\ : std_logic;
signal \N__50240\ : std_logic;
signal \N__50239\ : std_logic;
signal \N__50238\ : std_logic;
signal \N__50237\ : std_logic;
signal \N__50236\ : std_logic;
signal \N__50235\ : std_logic;
signal \N__50234\ : std_logic;
signal \N__50233\ : std_logic;
signal \N__50232\ : std_logic;
signal \N__50231\ : std_logic;
signal \N__50230\ : std_logic;
signal \N__50229\ : std_logic;
signal \N__50228\ : std_logic;
signal \N__50227\ : std_logic;
signal \N__50226\ : std_logic;
signal \N__50225\ : std_logic;
signal \N__50224\ : std_logic;
signal \N__50223\ : std_logic;
signal \N__50222\ : std_logic;
signal \N__50221\ : std_logic;
signal \N__50220\ : std_logic;
signal \N__50219\ : std_logic;
signal \N__50218\ : std_logic;
signal \N__50217\ : std_logic;
signal \N__50216\ : std_logic;
signal \N__50215\ : std_logic;
signal \N__50214\ : std_logic;
signal \N__50213\ : std_logic;
signal \N__50212\ : std_logic;
signal \N__50211\ : std_logic;
signal \N__50210\ : std_logic;
signal \N__50209\ : std_logic;
signal \N__50208\ : std_logic;
signal \N__50207\ : std_logic;
signal \N__50206\ : std_logic;
signal \N__50205\ : std_logic;
signal \N__50204\ : std_logic;
signal \N__50203\ : std_logic;
signal \N__50202\ : std_logic;
signal \N__50201\ : std_logic;
signal \N__50200\ : std_logic;
signal \N__50199\ : std_logic;
signal \N__50198\ : std_logic;
signal \N__50197\ : std_logic;
signal \N__50196\ : std_logic;
signal \N__50195\ : std_logic;
signal \N__50194\ : std_logic;
signal \N__50193\ : std_logic;
signal \N__50192\ : std_logic;
signal \N__50191\ : std_logic;
signal \N__50190\ : std_logic;
signal \N__50189\ : std_logic;
signal \N__50188\ : std_logic;
signal \N__50187\ : std_logic;
signal \N__50186\ : std_logic;
signal \N__50185\ : std_logic;
signal \N__50184\ : std_logic;
signal \N__50183\ : std_logic;
signal \N__50182\ : std_logic;
signal \N__50181\ : std_logic;
signal \N__50180\ : std_logic;
signal \N__50179\ : std_logic;
signal \N__50178\ : std_logic;
signal \N__50177\ : std_logic;
signal \N__50176\ : std_logic;
signal \N__50175\ : std_logic;
signal \N__50174\ : std_logic;
signal \N__50173\ : std_logic;
signal \N__50172\ : std_logic;
signal \N__50171\ : std_logic;
signal \N__50170\ : std_logic;
signal \N__50169\ : std_logic;
signal \N__50166\ : std_logic;
signal \N__50165\ : std_logic;
signal \N__49856\ : std_logic;
signal \N__49853\ : std_logic;
signal \N__49852\ : std_logic;
signal \N__49851\ : std_logic;
signal \N__49850\ : std_logic;
signal \N__49849\ : std_logic;
signal \N__49848\ : std_logic;
signal \N__49847\ : std_logic;
signal \N__49840\ : std_logic;
signal \N__49839\ : std_logic;
signal \N__49838\ : std_logic;
signal \N__49837\ : std_logic;
signal \N__49836\ : std_logic;
signal \N__49835\ : std_logic;
signal \N__49834\ : std_logic;
signal \N__49833\ : std_logic;
signal \N__49832\ : std_logic;
signal \N__49823\ : std_logic;
signal \N__49820\ : std_logic;
signal \N__49811\ : std_logic;
signal \N__49808\ : std_logic;
signal \N__49807\ : std_logic;
signal \N__49806\ : std_logic;
signal \N__49805\ : std_logic;
signal \N__49804\ : std_logic;
signal \N__49803\ : std_logic;
signal \N__49800\ : std_logic;
signal \N__49799\ : std_logic;
signal \N__49796\ : std_logic;
signal \N__49793\ : std_logic;
signal \N__49792\ : std_logic;
signal \N__49791\ : std_logic;
signal \N__49790\ : std_logic;
signal \N__49789\ : std_logic;
signal \N__49788\ : std_logic;
signal \N__49781\ : std_logic;
signal \N__49778\ : std_logic;
signal \N__49777\ : std_logic;
signal \N__49776\ : std_logic;
signal \N__49775\ : std_logic;
signal \N__49774\ : std_logic;
signal \N__49773\ : std_logic;
signal \N__49772\ : std_logic;
signal \N__49771\ : std_logic;
signal \N__49770\ : std_logic;
signal \N__49769\ : std_logic;
signal \N__49768\ : std_logic;
signal \N__49767\ : std_logic;
signal \N__49766\ : std_logic;
signal \N__49763\ : std_logic;
signal \N__49760\ : std_logic;
signal \N__49757\ : std_logic;
signal \N__49754\ : std_logic;
signal \N__49751\ : std_logic;
signal \N__49748\ : std_logic;
signal \N__49747\ : std_logic;
signal \N__49746\ : std_logic;
signal \N__49745\ : std_logic;
signal \N__49744\ : std_logic;
signal \N__49741\ : std_logic;
signal \N__49736\ : std_logic;
signal \N__49735\ : std_logic;
signal \N__49734\ : std_logic;
signal \N__49733\ : std_logic;
signal \N__49730\ : std_logic;
signal \N__49727\ : std_logic;
signal \N__49720\ : std_logic;
signal \N__49715\ : std_logic;
signal \N__49706\ : std_logic;
signal \N__49697\ : std_logic;
signal \N__49688\ : std_logic;
signal \N__49685\ : std_logic;
signal \N__49680\ : std_logic;
signal \N__49677\ : std_logic;
signal \N__49672\ : std_logic;
signal \N__49663\ : std_logic;
signal \N__49660\ : std_logic;
signal \N__49657\ : std_logic;
signal \N__49654\ : std_logic;
signal \N__49651\ : std_logic;
signal \N__49648\ : std_logic;
signal \N__49645\ : std_logic;
signal \N__49642\ : std_logic;
signal \N__49631\ : std_logic;
signal \N__49628\ : std_logic;
signal \N__49625\ : std_logic;
signal \N__49614\ : std_logic;
signal \N__49611\ : std_logic;
signal \N__49608\ : std_logic;
signal \N__49603\ : std_logic;
signal \N__49598\ : std_logic;
signal \N__49595\ : std_logic;
signal \N__49592\ : std_logic;
signal \N__49589\ : std_logic;
signal \N__49574\ : std_logic;
signal \N__49573\ : std_logic;
signal \N__49572\ : std_logic;
signal \N__49571\ : std_logic;
signal \N__49568\ : std_logic;
signal \N__49565\ : std_logic;
signal \N__49562\ : std_logic;
signal \N__49559\ : std_logic;
signal \N__49556\ : std_logic;
signal \N__49553\ : std_logic;
signal \N__49552\ : std_logic;
signal \N__49551\ : std_logic;
signal \N__49550\ : std_logic;
signal \N__49549\ : std_logic;
signal \N__49548\ : std_logic;
signal \N__49545\ : std_logic;
signal \N__49544\ : std_logic;
signal \N__49541\ : std_logic;
signal \N__49540\ : std_logic;
signal \N__49539\ : std_logic;
signal \N__49538\ : std_logic;
signal \N__49537\ : std_logic;
signal \N__49536\ : std_logic;
signal \N__49535\ : std_logic;
signal \N__49534\ : std_logic;
signal \N__49533\ : std_logic;
signal \N__49532\ : std_logic;
signal \N__49531\ : std_logic;
signal \N__49530\ : std_logic;
signal \N__49529\ : std_logic;
signal \N__49528\ : std_logic;
signal \N__49527\ : std_logic;
signal \N__49526\ : std_logic;
signal \N__49525\ : std_logic;
signal \N__49524\ : std_logic;
signal \N__49523\ : std_logic;
signal \N__49522\ : std_logic;
signal \N__49521\ : std_logic;
signal \N__49520\ : std_logic;
signal \N__49519\ : std_logic;
signal \N__49518\ : std_logic;
signal \N__49517\ : std_logic;
signal \N__49516\ : std_logic;
signal \N__49515\ : std_logic;
signal \N__49514\ : std_logic;
signal \N__49513\ : std_logic;
signal \N__49512\ : std_logic;
signal \N__49511\ : std_logic;
signal \N__49510\ : std_logic;
signal \N__49509\ : std_logic;
signal \N__49508\ : std_logic;
signal \N__49507\ : std_logic;
signal \N__49506\ : std_logic;
signal \N__49505\ : std_logic;
signal \N__49504\ : std_logic;
signal \N__49503\ : std_logic;
signal \N__49502\ : std_logic;
signal \N__49501\ : std_logic;
signal \N__49500\ : std_logic;
signal \N__49499\ : std_logic;
signal \N__49498\ : std_logic;
signal \N__49497\ : std_logic;
signal \N__49496\ : std_logic;
signal \N__49495\ : std_logic;
signal \N__49494\ : std_logic;
signal \N__49493\ : std_logic;
signal \N__49492\ : std_logic;
signal \N__49491\ : std_logic;
signal \N__49490\ : std_logic;
signal \N__49489\ : std_logic;
signal \N__49488\ : std_logic;
signal \N__49487\ : std_logic;
signal \N__49486\ : std_logic;
signal \N__49485\ : std_logic;
signal \N__49484\ : std_logic;
signal \N__49483\ : std_logic;
signal \N__49482\ : std_logic;
signal \N__49481\ : std_logic;
signal \N__49480\ : std_logic;
signal \N__49479\ : std_logic;
signal \N__49478\ : std_logic;
signal \N__49477\ : std_logic;
signal \N__49476\ : std_logic;
signal \N__49475\ : std_logic;
signal \N__49474\ : std_logic;
signal \N__49473\ : std_logic;
signal \N__49472\ : std_logic;
signal \N__49471\ : std_logic;
signal \N__49470\ : std_logic;
signal \N__49469\ : std_logic;
signal \N__49468\ : std_logic;
signal \N__49467\ : std_logic;
signal \N__49466\ : std_logic;
signal \N__49465\ : std_logic;
signal \N__49464\ : std_logic;
signal \N__49463\ : std_logic;
signal \N__49462\ : std_logic;
signal \N__49461\ : std_logic;
signal \N__49460\ : std_logic;
signal \N__49459\ : std_logic;
signal \N__49458\ : std_logic;
signal \N__49457\ : std_logic;
signal \N__49456\ : std_logic;
signal \N__49455\ : std_logic;
signal \N__49454\ : std_logic;
signal \N__49453\ : std_logic;
signal \N__49452\ : std_logic;
signal \N__49451\ : std_logic;
signal \N__49450\ : std_logic;
signal \N__49449\ : std_logic;
signal \N__49448\ : std_logic;
signal \N__49447\ : std_logic;
signal \N__49446\ : std_logic;
signal \N__49445\ : std_logic;
signal \N__49444\ : std_logic;
signal \N__49443\ : std_logic;
signal \N__49442\ : std_logic;
signal \N__49441\ : std_logic;
signal \N__49440\ : std_logic;
signal \N__49439\ : std_logic;
signal \N__49438\ : std_logic;
signal \N__49437\ : std_logic;
signal \N__49436\ : std_logic;
signal \N__49435\ : std_logic;
signal \N__49434\ : std_logic;
signal \N__49433\ : std_logic;
signal \N__49432\ : std_logic;
signal \N__49431\ : std_logic;
signal \N__49430\ : std_logic;
signal \N__49429\ : std_logic;
signal \N__49428\ : std_logic;
signal \N__49427\ : std_logic;
signal \N__49426\ : std_logic;
signal \N__49425\ : std_logic;
signal \N__49424\ : std_logic;
signal \N__49423\ : std_logic;
signal \N__49422\ : std_logic;
signal \N__49421\ : std_logic;
signal \N__49420\ : std_logic;
signal \N__49419\ : std_logic;
signal \N__49418\ : std_logic;
signal \N__49417\ : std_logic;
signal \N__49416\ : std_logic;
signal \N__49415\ : std_logic;
signal \N__49414\ : std_logic;
signal \N__49413\ : std_logic;
signal \N__49412\ : std_logic;
signal \N__49411\ : std_logic;
signal \N__49410\ : std_logic;
signal \N__49409\ : std_logic;
signal \N__49408\ : std_logic;
signal \N__49407\ : std_logic;
signal \N__49406\ : std_logic;
signal \N__49405\ : std_logic;
signal \N__49404\ : std_logic;
signal \N__49403\ : std_logic;
signal \N__49402\ : std_logic;
signal \N__49401\ : std_logic;
signal \N__49400\ : std_logic;
signal \N__49399\ : std_logic;
signal \N__49398\ : std_logic;
signal \N__49397\ : std_logic;
signal \N__49396\ : std_logic;
signal \N__49395\ : std_logic;
signal \N__49394\ : std_logic;
signal \N__49393\ : std_logic;
signal \N__49076\ : std_logic;
signal \N__49073\ : std_logic;
signal \N__49070\ : std_logic;
signal \N__49067\ : std_logic;
signal \N__49064\ : std_logic;
signal \N__49061\ : std_logic;
signal \N__49058\ : std_logic;
signal \N__49055\ : std_logic;
signal \N__49054\ : std_logic;
signal \N__49049\ : std_logic;
signal \N__49046\ : std_logic;
signal \N__49045\ : std_logic;
signal \N__49044\ : std_logic;
signal \N__49039\ : std_logic;
signal \N__49036\ : std_logic;
signal \N__49033\ : std_logic;
signal \N__49028\ : std_logic;
signal \N__49027\ : std_logic;
signal \N__49024\ : std_logic;
signal \N__49021\ : std_logic;
signal \N__49020\ : std_logic;
signal \N__49015\ : std_logic;
signal \N__49012\ : std_logic;
signal \N__49009\ : std_logic;
signal \N__49004\ : std_logic;
signal \N__49003\ : std_logic;
signal \N__48998\ : std_logic;
signal \N__48995\ : std_logic;
signal \N__48992\ : std_logic;
signal \N__48989\ : std_logic;
signal \N__48986\ : std_logic;
signal \N__48983\ : std_logic;
signal \N__48982\ : std_logic;
signal \N__48979\ : std_logic;
signal \N__48978\ : std_logic;
signal \N__48975\ : std_logic;
signal \N__48972\ : std_logic;
signal \N__48969\ : std_logic;
signal \N__48968\ : std_logic;
signal \N__48965\ : std_logic;
signal \N__48960\ : std_logic;
signal \N__48957\ : std_logic;
signal \N__48954\ : std_logic;
signal \N__48949\ : std_logic;
signal \N__48946\ : std_logic;
signal \N__48943\ : std_logic;
signal \N__48938\ : std_logic;
signal \N__48937\ : std_logic;
signal \N__48936\ : std_logic;
signal \N__48935\ : std_logic;
signal \N__48932\ : std_logic;
signal \N__48931\ : std_logic;
signal \N__48930\ : std_logic;
signal \N__48927\ : std_logic;
signal \N__48926\ : std_logic;
signal \N__48925\ : std_logic;
signal \N__48924\ : std_logic;
signal \N__48923\ : std_logic;
signal \N__48922\ : std_logic;
signal \N__48921\ : std_logic;
signal \N__48920\ : std_logic;
signal \N__48911\ : std_logic;
signal \N__48910\ : std_logic;
signal \N__48909\ : std_logic;
signal \N__48908\ : std_logic;
signal \N__48907\ : std_logic;
signal \N__48906\ : std_logic;
signal \N__48905\ : std_logic;
signal \N__48904\ : std_logic;
signal \N__48903\ : std_logic;
signal \N__48902\ : std_logic;
signal \N__48901\ : std_logic;
signal \N__48894\ : std_logic;
signal \N__48893\ : std_logic;
signal \N__48892\ : std_logic;
signal \N__48891\ : std_logic;
signal \N__48890\ : std_logic;
signal \N__48889\ : std_logic;
signal \N__48888\ : std_logic;
signal \N__48887\ : std_logic;
signal \N__48886\ : std_logic;
signal \N__48885\ : std_logic;
signal \N__48884\ : std_logic;
signal \N__48881\ : std_logic;
signal \N__48880\ : std_logic;
signal \N__48879\ : std_logic;
signal \N__48878\ : std_logic;
signal \N__48877\ : std_logic;
signal \N__48876\ : std_logic;
signal \N__48875\ : std_logic;
signal \N__48874\ : std_logic;
signal \N__48873\ : std_logic;
signal \N__48872\ : std_logic;
signal \N__48871\ : std_logic;
signal \N__48870\ : std_logic;
signal \N__48869\ : std_logic;
signal \N__48864\ : std_logic;
signal \N__48863\ : std_logic;
signal \N__48862\ : std_logic;
signal \N__48861\ : std_logic;
signal \N__48860\ : std_logic;
signal \N__48859\ : std_logic;
signal \N__48858\ : std_logic;
signal \N__48857\ : std_logic;
signal \N__48856\ : std_logic;
signal \N__48855\ : std_logic;
signal \N__48854\ : std_logic;
signal \N__48851\ : std_logic;
signal \N__48846\ : std_logic;
signal \N__48843\ : std_logic;
signal \N__48840\ : std_logic;
signal \N__48839\ : std_logic;
signal \N__48836\ : std_logic;
signal \N__48835\ : std_logic;
signal \N__48834\ : std_logic;
signal \N__48833\ : std_logic;
signal \N__48832\ : std_logic;
signal \N__48831\ : std_logic;
signal \N__48830\ : std_logic;
signal \N__48829\ : std_logic;
signal \N__48828\ : std_logic;
signal \N__48827\ : std_logic;
signal \N__48826\ : std_logic;
signal \N__48823\ : std_logic;
signal \N__48820\ : std_logic;
signal \N__48817\ : std_logic;
signal \N__48814\ : std_logic;
signal \N__48805\ : std_logic;
signal \N__48802\ : std_logic;
signal \N__48795\ : std_logic;
signal \N__48788\ : std_logic;
signal \N__48779\ : std_logic;
signal \N__48778\ : std_logic;
signal \N__48777\ : std_logic;
signal \N__48776\ : std_logic;
signal \N__48773\ : std_logic;
signal \N__48770\ : std_logic;
signal \N__48765\ : std_logic;
signal \N__48760\ : std_logic;
signal \N__48759\ : std_logic;
signal \N__48758\ : std_logic;
signal \N__48757\ : std_logic;
signal \N__48752\ : std_logic;
signal \N__48749\ : std_logic;
signal \N__48744\ : std_logic;
signal \N__48739\ : std_logic;
signal \N__48736\ : std_logic;
signal \N__48727\ : std_logic;
signal \N__48724\ : std_logic;
signal \N__48719\ : std_logic;
signal \N__48716\ : std_logic;
signal \N__48711\ : std_logic;
signal \N__48702\ : std_logic;
signal \N__48699\ : std_logic;
signal \N__48696\ : std_logic;
signal \N__48693\ : std_logic;
signal \N__48692\ : std_logic;
signal \N__48691\ : std_logic;
signal \N__48690\ : std_logic;
signal \N__48689\ : std_logic;
signal \N__48678\ : std_logic;
signal \N__48677\ : std_logic;
signal \N__48676\ : std_logic;
signal \N__48675\ : std_logic;
signal \N__48674\ : std_logic;
signal \N__48673\ : std_logic;
signal \N__48672\ : std_logic;
signal \N__48671\ : std_logic;
signal \N__48670\ : std_logic;
signal \N__48669\ : std_logic;
signal \N__48668\ : std_logic;
signal \N__48667\ : std_logic;
signal \N__48666\ : std_logic;
signal \N__48665\ : std_logic;
signal \N__48662\ : std_logic;
signal \N__48657\ : std_logic;
signal \N__48654\ : std_logic;
signal \N__48653\ : std_logic;
signal \N__48652\ : std_logic;
signal \N__48651\ : std_logic;
signal \N__48644\ : std_logic;
signal \N__48631\ : std_logic;
signal \N__48624\ : std_logic;
signal \N__48619\ : std_logic;
signal \N__48614\ : std_logic;
signal \N__48607\ : std_logic;
signal \N__48590\ : std_logic;
signal \N__48583\ : std_logic;
signal \N__48580\ : std_logic;
signal \N__48575\ : std_logic;
signal \N__48568\ : std_logic;
signal \N__48565\ : std_logic;
signal \N__48562\ : std_logic;
signal \N__48549\ : std_logic;
signal \N__48540\ : std_logic;
signal \N__48533\ : std_logic;
signal \N__48526\ : std_logic;
signal \N__48519\ : std_logic;
signal \N__48512\ : std_logic;
signal \N__48507\ : std_logic;
signal \N__48500\ : std_logic;
signal \N__48495\ : std_logic;
signal \N__48488\ : std_logic;
signal \N__48467\ : std_logic;
signal \N__48464\ : std_logic;
signal \N__48463\ : std_logic;
signal \N__48462\ : std_logic;
signal \N__48459\ : std_logic;
signal \N__48456\ : std_logic;
signal \N__48453\ : std_logic;
signal \N__48450\ : std_logic;
signal \N__48447\ : std_logic;
signal \N__48440\ : std_logic;
signal \N__48439\ : std_logic;
signal \N__48438\ : std_logic;
signal \N__48437\ : std_logic;
signal \N__48436\ : std_logic;
signal \N__48435\ : std_logic;
signal \N__48432\ : std_logic;
signal \N__48431\ : std_logic;
signal \N__48428\ : std_logic;
signal \N__48425\ : std_logic;
signal \N__48422\ : std_logic;
signal \N__48419\ : std_logic;
signal \N__48418\ : std_logic;
signal \N__48417\ : std_logic;
signal \N__48416\ : std_logic;
signal \N__48415\ : std_logic;
signal \N__48414\ : std_logic;
signal \N__48413\ : std_logic;
signal \N__48412\ : std_logic;
signal \N__48411\ : std_logic;
signal \N__48410\ : std_logic;
signal \N__48409\ : std_logic;
signal \N__48408\ : std_logic;
signal \N__48407\ : std_logic;
signal \N__48406\ : std_logic;
signal \N__48405\ : std_logic;
signal \N__48404\ : std_logic;
signal \N__48397\ : std_logic;
signal \N__48388\ : std_logic;
signal \N__48381\ : std_logic;
signal \N__48372\ : std_logic;
signal \N__48371\ : std_logic;
signal \N__48368\ : std_logic;
signal \N__48363\ : std_logic;
signal \N__48360\ : std_logic;
signal \N__48355\ : std_logic;
signal \N__48352\ : std_logic;
signal \N__48349\ : std_logic;
signal \N__48348\ : std_logic;
signal \N__48345\ : std_logic;
signal \N__48344\ : std_logic;
signal \N__48343\ : std_logic;
signal \N__48342\ : std_logic;
signal \N__48341\ : std_logic;
signal \N__48340\ : std_logic;
signal \N__48339\ : std_logic;
signal \N__48338\ : std_logic;
signal \N__48337\ : std_logic;
signal \N__48336\ : std_logic;
signal \N__48335\ : std_logic;
signal \N__48334\ : std_logic;
signal \N__48333\ : std_logic;
signal \N__48326\ : std_logic;
signal \N__48323\ : std_logic;
signal \N__48312\ : std_logic;
signal \N__48309\ : std_logic;
signal \N__48306\ : std_logic;
signal \N__48305\ : std_logic;
signal \N__48304\ : std_logic;
signal \N__48303\ : std_logic;
signal \N__48302\ : std_logic;
signal \N__48301\ : std_logic;
signal \N__48300\ : std_logic;
signal \N__48299\ : std_logic;
signal \N__48296\ : std_logic;
signal \N__48295\ : std_logic;
signal \N__48292\ : std_logic;
signal \N__48291\ : std_logic;
signal \N__48288\ : std_logic;
signal \N__48287\ : std_logic;
signal \N__48284\ : std_logic;
signal \N__48283\ : std_logic;
signal \N__48280\ : std_logic;
signal \N__48279\ : std_logic;
signal \N__48276\ : std_logic;
signal \N__48275\ : std_logic;
signal \N__48272\ : std_logic;
signal \N__48271\ : std_logic;
signal \N__48268\ : std_logic;
signal \N__48267\ : std_logic;
signal \N__48264\ : std_logic;
signal \N__48263\ : std_logic;
signal \N__48260\ : std_logic;
signal \N__48259\ : std_logic;
signal \N__48256\ : std_logic;
signal \N__48255\ : std_logic;
signal \N__48252\ : std_logic;
signal \N__48251\ : std_logic;
signal \N__48250\ : std_logic;
signal \N__48249\ : std_logic;
signal \N__48248\ : std_logic;
signal \N__48245\ : std_logic;
signal \N__48238\ : std_logic;
signal \N__48235\ : std_logic;
signal \N__48232\ : std_logic;
signal \N__48225\ : std_logic;
signal \N__48216\ : std_logic;
signal \N__48213\ : std_logic;
signal \N__48198\ : std_logic;
signal \N__48181\ : std_logic;
signal \N__48164\ : std_logic;
signal \N__48163\ : std_logic;
signal \N__48160\ : std_logic;
signal \N__48159\ : std_logic;
signal \N__48156\ : std_logic;
signal \N__48155\ : std_logic;
signal \N__48152\ : std_logic;
signal \N__48151\ : std_logic;
signal \N__48150\ : std_logic;
signal \N__48147\ : std_logic;
signal \N__48144\ : std_logic;
signal \N__48139\ : std_logic;
signal \N__48134\ : std_logic;
signal \N__48129\ : std_logic;
signal \N__48126\ : std_logic;
signal \N__48123\ : std_logic;
signal \N__48108\ : std_logic;
signal \N__48105\ : std_logic;
signal \N__48102\ : std_logic;
signal \N__48095\ : std_logic;
signal \N__48084\ : std_logic;
signal \N__48081\ : std_logic;
signal \N__48078\ : std_logic;
signal \N__48075\ : std_logic;
signal \N__48072\ : std_logic;
signal \N__48065\ : std_logic;
signal \N__48064\ : std_logic;
signal \N__48063\ : std_logic;
signal \N__48060\ : std_logic;
signal \N__48057\ : std_logic;
signal \N__48054\ : std_logic;
signal \N__48051\ : std_logic;
signal \N__48048\ : std_logic;
signal \N__48047\ : std_logic;
signal \N__48044\ : std_logic;
signal \N__48041\ : std_logic;
signal \N__48038\ : std_logic;
signal \N__48035\ : std_logic;
signal \N__48032\ : std_logic;
signal \N__48027\ : std_logic;
signal \N__48020\ : std_logic;
signal \N__48017\ : std_logic;
signal \N__48014\ : std_logic;
signal \N__48013\ : std_logic;
signal \N__48010\ : std_logic;
signal \N__48007\ : std_logic;
signal \N__48004\ : std_logic;
signal \N__48001\ : std_logic;
signal \N__48000\ : std_logic;
signal \N__47997\ : std_logic;
signal \N__47996\ : std_logic;
signal \N__47993\ : std_logic;
signal \N__47990\ : std_logic;
signal \N__47987\ : std_logic;
signal \N__47984\ : std_logic;
signal \N__47981\ : std_logic;
signal \N__47978\ : std_logic;
signal \N__47969\ : std_logic;
signal \N__47966\ : std_logic;
signal \N__47963\ : std_logic;
signal \N__47962\ : std_logic;
signal \N__47959\ : std_logic;
signal \N__47956\ : std_logic;
signal \N__47953\ : std_logic;
signal \N__47950\ : std_logic;
signal \N__47945\ : std_logic;
signal \N__47944\ : std_logic;
signal \N__47943\ : std_logic;
signal \N__47940\ : std_logic;
signal \N__47937\ : std_logic;
signal \N__47934\ : std_logic;
signal \N__47931\ : std_logic;
signal \N__47924\ : std_logic;
signal \N__47923\ : std_logic;
signal \N__47922\ : std_logic;
signal \N__47919\ : std_logic;
signal \N__47916\ : std_logic;
signal \N__47913\ : std_logic;
signal \N__47908\ : std_logic;
signal \N__47907\ : std_logic;
signal \N__47904\ : std_logic;
signal \N__47901\ : std_logic;
signal \N__47898\ : std_logic;
signal \N__47891\ : std_logic;
signal \N__47890\ : std_logic;
signal \N__47885\ : std_logic;
signal \N__47882\ : std_logic;
signal \N__47879\ : std_logic;
signal \N__47876\ : std_logic;
signal \N__47873\ : std_logic;
signal \N__47872\ : std_logic;
signal \N__47871\ : std_logic;
signal \N__47870\ : std_logic;
signal \N__47869\ : std_logic;
signal \N__47868\ : std_logic;
signal \N__47867\ : std_logic;
signal \N__47866\ : std_logic;
signal \N__47865\ : std_logic;
signal \N__47864\ : std_logic;
signal \N__47863\ : std_logic;
signal \N__47862\ : std_logic;
signal \N__47861\ : std_logic;
signal \N__47860\ : std_logic;
signal \N__47831\ : std_logic;
signal \N__47828\ : std_logic;
signal \N__47825\ : std_logic;
signal \N__47824\ : std_logic;
signal \N__47823\ : std_logic;
signal \N__47820\ : std_logic;
signal \N__47817\ : std_logic;
signal \N__47814\ : std_logic;
signal \N__47807\ : std_logic;
signal \N__47804\ : std_logic;
signal \N__47803\ : std_logic;
signal \N__47802\ : std_logic;
signal \N__47799\ : std_logic;
signal \N__47796\ : std_logic;
signal \N__47793\ : std_logic;
signal \N__47792\ : std_logic;
signal \N__47789\ : std_logic;
signal \N__47784\ : std_logic;
signal \N__47781\ : std_logic;
signal \N__47778\ : std_logic;
signal \N__47775\ : std_logic;
signal \N__47772\ : std_logic;
signal \N__47765\ : std_logic;
signal \N__47764\ : std_logic;
signal \N__47759\ : std_logic;
signal \N__47756\ : std_logic;
signal \N__47753\ : std_logic;
signal \N__47750\ : std_logic;
signal \N__47749\ : std_logic;
signal \N__47748\ : std_logic;
signal \N__47745\ : std_logic;
signal \N__47742\ : std_logic;
signal \N__47739\ : std_logic;
signal \N__47734\ : std_logic;
signal \N__47729\ : std_logic;
signal \N__47728\ : std_logic;
signal \N__47727\ : std_logic;
signal \N__47724\ : std_logic;
signal \N__47721\ : std_logic;
signal \N__47720\ : std_logic;
signal \N__47717\ : std_logic;
signal \N__47714\ : std_logic;
signal \N__47711\ : std_logic;
signal \N__47708\ : std_logic;
signal \N__47705\ : std_logic;
signal \N__47700\ : std_logic;
signal \N__47697\ : std_logic;
signal \N__47690\ : std_logic;
signal \N__47687\ : std_logic;
signal \N__47684\ : std_logic;
signal \N__47681\ : std_logic;
signal \N__47678\ : std_logic;
signal \N__47675\ : std_logic;
signal \N__47672\ : std_logic;
signal \N__47669\ : std_logic;
signal \N__47668\ : std_logic;
signal \N__47665\ : std_logic;
signal \N__47662\ : std_logic;
signal \N__47657\ : std_logic;
signal \N__47656\ : std_logic;
signal \N__47655\ : std_logic;
signal \N__47650\ : std_logic;
signal \N__47647\ : std_logic;
signal \N__47644\ : std_logic;
signal \N__47643\ : std_logic;
signal \N__47640\ : std_logic;
signal \N__47637\ : std_logic;
signal \N__47634\ : std_logic;
signal \N__47629\ : std_logic;
signal \N__47626\ : std_logic;
signal \N__47621\ : std_logic;
signal \N__47618\ : std_logic;
signal \N__47617\ : std_logic;
signal \N__47612\ : std_logic;
signal \N__47609\ : std_logic;
signal \N__47608\ : std_logic;
signal \N__47603\ : std_logic;
signal \N__47602\ : std_logic;
signal \N__47599\ : std_logic;
signal \N__47596\ : std_logic;
signal \N__47593\ : std_logic;
signal \N__47588\ : std_logic;
signal \N__47587\ : std_logic;
signal \N__47584\ : std_logic;
signal \N__47581\ : std_logic;
signal \N__47576\ : std_logic;
signal \N__47575\ : std_logic;
signal \N__47572\ : std_logic;
signal \N__47569\ : std_logic;
signal \N__47566\ : std_logic;
signal \N__47561\ : std_logic;
signal \N__47560\ : std_logic;
signal \N__47555\ : std_logic;
signal \N__47552\ : std_logic;
signal \N__47549\ : std_logic;
signal \N__47546\ : std_logic;
signal \N__47543\ : std_logic;
signal \N__47540\ : std_logic;
signal \N__47537\ : std_logic;
signal \N__47534\ : std_logic;
signal \N__47533\ : std_logic;
signal \N__47530\ : std_logic;
signal \N__47527\ : std_logic;
signal \N__47522\ : std_logic;
signal \N__47521\ : std_logic;
signal \N__47520\ : std_logic;
signal \N__47515\ : std_logic;
signal \N__47512\ : std_logic;
signal \N__47509\ : std_logic;
signal \N__47508\ : std_logic;
signal \N__47505\ : std_logic;
signal \N__47502\ : std_logic;
signal \N__47499\ : std_logic;
signal \N__47492\ : std_logic;
signal \N__47489\ : std_logic;
signal \N__47486\ : std_logic;
signal \N__47483\ : std_logic;
signal \N__47480\ : std_logic;
signal \N__47477\ : std_logic;
signal \N__47476\ : std_logic;
signal \N__47475\ : std_logic;
signal \N__47472\ : std_logic;
signal \N__47469\ : std_logic;
signal \N__47466\ : std_logic;
signal \N__47461\ : std_logic;
signal \N__47456\ : std_logic;
signal \N__47455\ : std_logic;
signal \N__47452\ : std_logic;
signal \N__47449\ : std_logic;
signal \N__47448\ : std_logic;
signal \N__47447\ : std_logic;
signal \N__47444\ : std_logic;
signal \N__47441\ : std_logic;
signal \N__47438\ : std_logic;
signal \N__47435\ : std_logic;
signal \N__47430\ : std_logic;
signal \N__47427\ : std_logic;
signal \N__47424\ : std_logic;
signal \N__47419\ : std_logic;
signal \N__47416\ : std_logic;
signal \N__47413\ : std_logic;
signal \N__47408\ : std_logic;
signal \N__47405\ : std_logic;
signal \N__47402\ : std_logic;
signal \N__47399\ : std_logic;
signal \N__47396\ : std_logic;
signal \N__47395\ : std_logic;
signal \N__47394\ : std_logic;
signal \N__47389\ : std_logic;
signal \N__47386\ : std_logic;
signal \N__47383\ : std_logic;
signal \N__47378\ : std_logic;
signal \N__47375\ : std_logic;
signal \N__47374\ : std_logic;
signal \N__47373\ : std_logic;
signal \N__47368\ : std_logic;
signal \N__47365\ : std_logic;
signal \N__47362\ : std_logic;
signal \N__47357\ : std_logic;
signal \N__47354\ : std_logic;
signal \N__47353\ : std_logic;
signal \N__47348\ : std_logic;
signal \N__47345\ : std_logic;
signal \N__47342\ : std_logic;
signal \N__47339\ : std_logic;
signal \N__47336\ : std_logic;
signal \N__47333\ : std_logic;
signal \N__47330\ : std_logic;
signal \N__47327\ : std_logic;
signal \N__47324\ : std_logic;
signal \N__47323\ : std_logic;
signal \N__47320\ : std_logic;
signal \N__47317\ : std_logic;
signal \N__47312\ : std_logic;
signal \N__47311\ : std_logic;
signal \N__47306\ : std_logic;
signal \N__47305\ : std_logic;
signal \N__47302\ : std_logic;
signal \N__47301\ : std_logic;
signal \N__47298\ : std_logic;
signal \N__47295\ : std_logic;
signal \N__47292\ : std_logic;
signal \N__47289\ : std_logic;
signal \N__47284\ : std_logic;
signal \N__47281\ : std_logic;
signal \N__47278\ : std_logic;
signal \N__47273\ : std_logic;
signal \N__47270\ : std_logic;
signal \N__47269\ : std_logic;
signal \N__47264\ : std_logic;
signal \N__47261\ : std_logic;
signal \N__47260\ : std_logic;
signal \N__47255\ : std_logic;
signal \N__47252\ : std_logic;
signal \N__47249\ : std_logic;
signal \N__47248\ : std_logic;
signal \N__47245\ : std_logic;
signal \N__47242\ : std_logic;
signal \N__47237\ : std_logic;
signal \N__47234\ : std_logic;
signal \N__47231\ : std_logic;
signal \N__47228\ : std_logic;
signal \N__47227\ : std_logic;
signal \N__47224\ : std_logic;
signal \N__47221\ : std_logic;
signal \N__47216\ : std_logic;
signal \N__47215\ : std_logic;
signal \N__47210\ : std_logic;
signal \N__47209\ : std_logic;
signal \N__47206\ : std_logic;
signal \N__47203\ : std_logic;
signal \N__47200\ : std_logic;
signal \N__47199\ : std_logic;
signal \N__47196\ : std_logic;
signal \N__47193\ : std_logic;
signal \N__47190\ : std_logic;
signal \N__47183\ : std_logic;
signal \N__47180\ : std_logic;
signal \N__47179\ : std_logic;
signal \N__47178\ : std_logic;
signal \N__47175\ : std_logic;
signal \N__47170\ : std_logic;
signal \N__47165\ : std_logic;
signal \N__47162\ : std_logic;
signal \N__47161\ : std_logic;
signal \N__47158\ : std_logic;
signal \N__47155\ : std_logic;
signal \N__47150\ : std_logic;
signal \N__47149\ : std_logic;
signal \N__47146\ : std_logic;
signal \N__47143\ : std_logic;
signal \N__47140\ : std_logic;
signal \N__47135\ : std_logic;
signal \N__47132\ : std_logic;
signal \N__47131\ : std_logic;
signal \N__47126\ : std_logic;
signal \N__47123\ : std_logic;
signal \N__47120\ : std_logic;
signal \N__47117\ : std_logic;
signal \N__47114\ : std_logic;
signal \N__47111\ : std_logic;
signal \N__47108\ : std_logic;
signal \N__47107\ : std_logic;
signal \N__47104\ : std_logic;
signal \N__47101\ : std_logic;
signal \N__47098\ : std_logic;
signal \N__47093\ : std_logic;
signal \N__47092\ : std_logic;
signal \N__47091\ : std_logic;
signal \N__47086\ : std_logic;
signal \N__47083\ : std_logic;
signal \N__47080\ : std_logic;
signal \N__47079\ : std_logic;
signal \N__47076\ : std_logic;
signal \N__47073\ : std_logic;
signal \N__47070\ : std_logic;
signal \N__47063\ : std_logic;
signal \N__47060\ : std_logic;
signal \N__47057\ : std_logic;
signal \N__47054\ : std_logic;
signal \N__47051\ : std_logic;
signal \N__47048\ : std_logic;
signal \N__47047\ : std_logic;
signal \N__47042\ : std_logic;
signal \N__47039\ : std_logic;
signal \N__47036\ : std_logic;
signal \N__47033\ : std_logic;
signal \N__47032\ : std_logic;
signal \N__47027\ : std_logic;
signal \N__47024\ : std_logic;
signal \N__47021\ : std_logic;
signal \N__47018\ : std_logic;
signal \N__47015\ : std_logic;
signal \N__47012\ : std_logic;
signal \N__47009\ : std_logic;
signal \N__47006\ : std_logic;
signal \N__47003\ : std_logic;
signal \N__47002\ : std_logic;
signal \N__46999\ : std_logic;
signal \N__46996\ : std_logic;
signal \N__46993\ : std_logic;
signal \N__46988\ : std_logic;
signal \N__46987\ : std_logic;
signal \N__46986\ : std_logic;
signal \N__46985\ : std_logic;
signal \N__46982\ : std_logic;
signal \N__46981\ : std_logic;
signal \N__46974\ : std_logic;
signal \N__46971\ : std_logic;
signal \N__46968\ : std_logic;
signal \N__46965\ : std_logic;
signal \N__46958\ : std_logic;
signal \N__46957\ : std_logic;
signal \N__46954\ : std_logic;
signal \N__46951\ : std_logic;
signal \N__46950\ : std_logic;
signal \N__46947\ : std_logic;
signal \N__46942\ : std_logic;
signal \N__46939\ : std_logic;
signal \N__46936\ : std_logic;
signal \N__46931\ : std_logic;
signal \N__46930\ : std_logic;
signal \N__46927\ : std_logic;
signal \N__46926\ : std_logic;
signal \N__46923\ : std_logic;
signal \N__46920\ : std_logic;
signal \N__46917\ : std_logic;
signal \N__46916\ : std_logic;
signal \N__46913\ : std_logic;
signal \N__46910\ : std_logic;
signal \N__46907\ : std_logic;
signal \N__46904\ : std_logic;
signal \N__46901\ : std_logic;
signal \N__46896\ : std_logic;
signal \N__46895\ : std_logic;
signal \N__46894\ : std_logic;
signal \N__46891\ : std_logic;
signal \N__46888\ : std_logic;
signal \N__46885\ : std_logic;
signal \N__46880\ : std_logic;
signal \N__46871\ : std_logic;
signal \N__46868\ : std_logic;
signal \N__46865\ : std_logic;
signal \N__46862\ : std_logic;
signal \N__46859\ : std_logic;
signal \N__46856\ : std_logic;
signal \N__46853\ : std_logic;
signal \N__46852\ : std_logic;
signal \N__46851\ : std_logic;
signal \N__46850\ : std_logic;
signal \N__46845\ : std_logic;
signal \N__46840\ : std_logic;
signal \N__46835\ : std_logic;
signal \N__46834\ : std_logic;
signal \N__46833\ : std_logic;
signal \N__46828\ : std_logic;
signal \N__46825\ : std_logic;
signal \N__46822\ : std_logic;
signal \N__46821\ : std_logic;
signal \N__46820\ : std_logic;
signal \N__46817\ : std_logic;
signal \N__46814\ : std_logic;
signal \N__46809\ : std_logic;
signal \N__46802\ : std_logic;
signal \N__46799\ : std_logic;
signal \N__46796\ : std_logic;
signal \N__46793\ : std_logic;
signal \N__46790\ : std_logic;
signal \N__46787\ : std_logic;
signal \N__46784\ : std_logic;
signal \N__46781\ : std_logic;
signal \N__46778\ : std_logic;
signal \N__46777\ : std_logic;
signal \N__46776\ : std_logic;
signal \N__46773\ : std_logic;
signal \N__46770\ : std_logic;
signal \N__46767\ : std_logic;
signal \N__46762\ : std_logic;
signal \N__46757\ : std_logic;
signal \N__46754\ : std_logic;
signal \N__46751\ : std_logic;
signal \N__46748\ : std_logic;
signal \N__46747\ : std_logic;
signal \N__46744\ : std_logic;
signal \N__46741\ : std_logic;
signal \N__46740\ : std_logic;
signal \N__46735\ : std_logic;
signal \N__46732\ : std_logic;
signal \N__46729\ : std_logic;
signal \N__46724\ : std_logic;
signal \N__46721\ : std_logic;
signal \N__46718\ : std_logic;
signal \N__46717\ : std_logic;
signal \N__46714\ : std_logic;
signal \N__46711\ : std_logic;
signal \N__46708\ : std_logic;
signal \N__46703\ : std_logic;
signal \N__46700\ : std_logic;
signal \N__46699\ : std_logic;
signal \N__46698\ : std_logic;
signal \N__46697\ : std_logic;
signal \N__46696\ : std_logic;
signal \N__46695\ : std_logic;
signal \N__46694\ : std_logic;
signal \N__46693\ : std_logic;
signal \N__46684\ : std_logic;
signal \N__46675\ : std_logic;
signal \N__46674\ : std_logic;
signal \N__46673\ : std_logic;
signal \N__46672\ : std_logic;
signal \N__46671\ : std_logic;
signal \N__46670\ : std_logic;
signal \N__46669\ : std_logic;
signal \N__46668\ : std_logic;
signal \N__46667\ : std_logic;
signal \N__46666\ : std_logic;
signal \N__46665\ : std_logic;
signal \N__46664\ : std_logic;
signal \N__46663\ : std_logic;
signal \N__46662\ : std_logic;
signal \N__46661\ : std_logic;
signal \N__46660\ : std_logic;
signal \N__46659\ : std_logic;
signal \N__46658\ : std_logic;
signal \N__46657\ : std_logic;
signal \N__46656\ : std_logic;
signal \N__46655\ : std_logic;
signal \N__46654\ : std_logic;
signal \N__46653\ : std_logic;
signal \N__46648\ : std_logic;
signal \N__46639\ : std_logic;
signal \N__46634\ : std_logic;
signal \N__46625\ : std_logic;
signal \N__46616\ : std_logic;
signal \N__46607\ : std_logic;
signal \N__46598\ : std_logic;
signal \N__46591\ : std_logic;
signal \N__46582\ : std_logic;
signal \N__46577\ : std_logic;
signal \N__46574\ : std_logic;
signal \N__46571\ : std_logic;
signal \N__46568\ : std_logic;
signal \N__46567\ : std_logic;
signal \N__46564\ : std_logic;
signal \N__46561\ : std_logic;
signal \N__46558\ : std_logic;
signal \N__46553\ : std_logic;
signal \N__46552\ : std_logic;
signal \N__46551\ : std_logic;
signal \N__46548\ : std_logic;
signal \N__46545\ : std_logic;
signal \N__46544\ : std_logic;
signal \N__46541\ : std_logic;
signal \N__46538\ : std_logic;
signal \N__46535\ : std_logic;
signal \N__46532\ : std_logic;
signal \N__46529\ : std_logic;
signal \N__46526\ : std_logic;
signal \N__46523\ : std_logic;
signal \N__46520\ : std_logic;
signal \N__46517\ : std_logic;
signal \N__46514\ : std_logic;
signal \N__46509\ : std_logic;
signal \N__46502\ : std_logic;
signal \N__46499\ : std_logic;
signal \N__46498\ : std_logic;
signal \N__46495\ : std_logic;
signal \N__46492\ : std_logic;
signal \N__46487\ : std_logic;
signal \N__46484\ : std_logic;
signal \N__46483\ : std_logic;
signal \N__46480\ : std_logic;
signal \N__46477\ : std_logic;
signal \N__46476\ : std_logic;
signal \N__46471\ : std_logic;
signal \N__46468\ : std_logic;
signal \N__46465\ : std_logic;
signal \N__46460\ : std_logic;
signal \N__46459\ : std_logic;
signal \N__46458\ : std_logic;
signal \N__46455\ : std_logic;
signal \N__46452\ : std_logic;
signal \N__46449\ : std_logic;
signal \N__46448\ : std_logic;
signal \N__46445\ : std_logic;
signal \N__46442\ : std_logic;
signal \N__46439\ : std_logic;
signal \N__46436\ : std_logic;
signal \N__46431\ : std_logic;
signal \N__46428\ : std_logic;
signal \N__46421\ : std_logic;
signal \N__46418\ : std_logic;
signal \N__46415\ : std_logic;
signal \N__46414\ : std_logic;
signal \N__46413\ : std_logic;
signal \N__46410\ : std_logic;
signal \N__46409\ : std_logic;
signal \N__46406\ : std_logic;
signal \N__46403\ : std_logic;
signal \N__46400\ : std_logic;
signal \N__46397\ : std_logic;
signal \N__46394\ : std_logic;
signal \N__46385\ : std_logic;
signal \N__46384\ : std_logic;
signal \N__46383\ : std_logic;
signal \N__46380\ : std_logic;
signal \N__46379\ : std_logic;
signal \N__46376\ : std_logic;
signal \N__46373\ : std_logic;
signal \N__46370\ : std_logic;
signal \N__46367\ : std_logic;
signal \N__46364\ : std_logic;
signal \N__46361\ : std_logic;
signal \N__46358\ : std_logic;
signal \N__46355\ : std_logic;
signal \N__46350\ : std_logic;
signal \N__46347\ : std_logic;
signal \N__46340\ : std_logic;
signal \N__46339\ : std_logic;
signal \N__46336\ : std_logic;
signal \N__46335\ : std_logic;
signal \N__46332\ : std_logic;
signal \N__46331\ : std_logic;
signal \N__46328\ : std_logic;
signal \N__46325\ : std_logic;
signal \N__46322\ : std_logic;
signal \N__46319\ : std_logic;
signal \N__46316\ : std_logic;
signal \N__46309\ : std_logic;
signal \N__46304\ : std_logic;
signal \N__46301\ : std_logic;
signal \N__46298\ : std_logic;
signal \N__46297\ : std_logic;
signal \N__46296\ : std_logic;
signal \N__46293\ : std_logic;
signal \N__46290\ : std_logic;
signal \N__46287\ : std_logic;
signal \N__46282\ : std_logic;
signal \N__46277\ : std_logic;
signal \N__46274\ : std_logic;
signal \N__46271\ : std_logic;
signal \N__46270\ : std_logic;
signal \N__46265\ : std_logic;
signal \N__46264\ : std_logic;
signal \N__46261\ : std_logic;
signal \N__46258\ : std_logic;
signal \N__46255\ : std_logic;
signal \N__46250\ : std_logic;
signal \N__46247\ : std_logic;
signal \N__46244\ : std_logic;
signal \N__46243\ : std_logic;
signal \N__46240\ : std_logic;
signal \N__46237\ : std_logic;
signal \N__46236\ : std_logic;
signal \N__46231\ : std_logic;
signal \N__46228\ : std_logic;
signal \N__46225\ : std_logic;
signal \N__46220\ : std_logic;
signal \N__46217\ : std_logic;
signal \N__46216\ : std_logic;
signal \N__46213\ : std_logic;
signal \N__46210\ : std_logic;
signal \N__46205\ : std_logic;
signal \N__46204\ : std_logic;
signal \N__46201\ : std_logic;
signal \N__46198\ : std_logic;
signal \N__46195\ : std_logic;
signal \N__46190\ : std_logic;
signal \N__46187\ : std_logic;
signal \N__46186\ : std_logic;
signal \N__46181\ : std_logic;
signal \N__46180\ : std_logic;
signal \N__46177\ : std_logic;
signal \N__46174\ : std_logic;
signal \N__46171\ : std_logic;
signal \N__46166\ : std_logic;
signal \N__46163\ : std_logic;
signal \N__46162\ : std_logic;
signal \N__46157\ : std_logic;
signal \N__46156\ : std_logic;
signal \N__46153\ : std_logic;
signal \N__46150\ : std_logic;
signal \N__46147\ : std_logic;
signal \N__46142\ : std_logic;
signal \N__46139\ : std_logic;
signal \N__46138\ : std_logic;
signal \N__46135\ : std_logic;
signal \N__46132\ : std_logic;
signal \N__46129\ : std_logic;
signal \N__46126\ : std_logic;
signal \N__46125\ : std_logic;
signal \N__46122\ : std_logic;
signal \N__46119\ : std_logic;
signal \N__46116\ : std_logic;
signal \N__46113\ : std_logic;
signal \N__46110\ : std_logic;
signal \N__46103\ : std_logic;
signal \N__46100\ : std_logic;
signal \N__46099\ : std_logic;
signal \N__46096\ : std_logic;
signal \N__46093\ : std_logic;
signal \N__46090\ : std_logic;
signal \N__46087\ : std_logic;
signal \N__46086\ : std_logic;
signal \N__46083\ : std_logic;
signal \N__46080\ : std_logic;
signal \N__46077\ : std_logic;
signal \N__46074\ : std_logic;
signal \N__46071\ : std_logic;
signal \N__46064\ : std_logic;
signal \N__46061\ : std_logic;
signal \N__46058\ : std_logic;
signal \N__46057\ : std_logic;
signal \N__46054\ : std_logic;
signal \N__46051\ : std_logic;
signal \N__46050\ : std_logic;
signal \N__46047\ : std_logic;
signal \N__46044\ : std_logic;
signal \N__46041\ : std_logic;
signal \N__46038\ : std_logic;
signal \N__46035\ : std_logic;
signal \N__46028\ : std_logic;
signal \N__46025\ : std_logic;
signal \N__46024\ : std_logic;
signal \N__46023\ : std_logic;
signal \N__46018\ : std_logic;
signal \N__46015\ : std_logic;
signal \N__46012\ : std_logic;
signal \N__46007\ : std_logic;
signal \N__46004\ : std_logic;
signal \N__46001\ : std_logic;
signal \N__46000\ : std_logic;
signal \N__45995\ : std_logic;
signal \N__45994\ : std_logic;
signal \N__45991\ : std_logic;
signal \N__45988\ : std_logic;
signal \N__45985\ : std_logic;
signal \N__45980\ : std_logic;
signal \N__45977\ : std_logic;
signal \N__45976\ : std_logic;
signal \N__45973\ : std_logic;
signal \N__45970\ : std_logic;
signal \N__45965\ : std_logic;
signal \N__45964\ : std_logic;
signal \N__45961\ : std_logic;
signal \N__45958\ : std_logic;
signal \N__45955\ : std_logic;
signal \N__45950\ : std_logic;
signal \N__45947\ : std_logic;
signal \N__45946\ : std_logic;
signal \N__45943\ : std_logic;
signal \N__45940\ : std_logic;
signal \N__45935\ : std_logic;
signal \N__45934\ : std_logic;
signal \N__45931\ : std_logic;
signal \N__45928\ : std_logic;
signal \N__45925\ : std_logic;
signal \N__45920\ : std_logic;
signal \N__45917\ : std_logic;
signal \N__45916\ : std_logic;
signal \N__45911\ : std_logic;
signal \N__45910\ : std_logic;
signal \N__45907\ : std_logic;
signal \N__45904\ : std_logic;
signal \N__45901\ : std_logic;
signal \N__45896\ : std_logic;
signal \N__45893\ : std_logic;
signal \N__45890\ : std_logic;
signal \N__45889\ : std_logic;
signal \N__45886\ : std_logic;
signal \N__45883\ : std_logic;
signal \N__45882\ : std_logic;
signal \N__45877\ : std_logic;
signal \N__45874\ : std_logic;
signal \N__45871\ : std_logic;
signal \N__45866\ : std_logic;
signal \N__45863\ : std_logic;
signal \N__45862\ : std_logic;
signal \N__45859\ : std_logic;
signal \N__45856\ : std_logic;
signal \N__45853\ : std_logic;
signal \N__45850\ : std_logic;
signal \N__45849\ : std_logic;
signal \N__45846\ : std_logic;
signal \N__45843\ : std_logic;
signal \N__45840\ : std_logic;
signal \N__45837\ : std_logic;
signal \N__45834\ : std_logic;
signal \N__45827\ : std_logic;
signal \N__45824\ : std_logic;
signal \N__45821\ : std_logic;
signal \N__45820\ : std_logic;
signal \N__45817\ : std_logic;
signal \N__45814\ : std_logic;
signal \N__45813\ : std_logic;
signal \N__45810\ : std_logic;
signal \N__45807\ : std_logic;
signal \N__45804\ : std_logic;
signal \N__45801\ : std_logic;
signal \N__45798\ : std_logic;
signal \N__45791\ : std_logic;
signal \N__45790\ : std_logic;
signal \N__45787\ : std_logic;
signal \N__45784\ : std_logic;
signal \N__45783\ : std_logic;
signal \N__45780\ : std_logic;
signal \N__45777\ : std_logic;
signal \N__45774\ : std_logic;
signal \N__45771\ : std_logic;
signal \N__45764\ : std_logic;
signal \N__45761\ : std_logic;
signal \N__45760\ : std_logic;
signal \N__45757\ : std_logic;
signal \N__45754\ : std_logic;
signal \N__45753\ : std_logic;
signal \N__45748\ : std_logic;
signal \N__45745\ : std_logic;
signal \N__45742\ : std_logic;
signal \N__45737\ : std_logic;
signal \N__45734\ : std_logic;
signal \N__45731\ : std_logic;
signal \N__45730\ : std_logic;
signal \N__45727\ : std_logic;
signal \N__45724\ : std_logic;
signal \N__45719\ : std_logic;
signal \N__45718\ : std_logic;
signal \N__45715\ : std_logic;
signal \N__45712\ : std_logic;
signal \N__45709\ : std_logic;
signal \N__45704\ : std_logic;
signal \N__45701\ : std_logic;
signal \N__45698\ : std_logic;
signal \N__45697\ : std_logic;
signal \N__45694\ : std_logic;
signal \N__45691\ : std_logic;
signal \N__45690\ : std_logic;
signal \N__45685\ : std_logic;
signal \N__45682\ : std_logic;
signal \N__45679\ : std_logic;
signal \N__45674\ : std_logic;
signal \N__45671\ : std_logic;
signal \N__45668\ : std_logic;
signal \N__45667\ : std_logic;
signal \N__45664\ : std_logic;
signal \N__45661\ : std_logic;
signal \N__45660\ : std_logic;
signal \N__45655\ : std_logic;
signal \N__45652\ : std_logic;
signal \N__45649\ : std_logic;
signal \N__45644\ : std_logic;
signal \N__45641\ : std_logic;
signal \N__45638\ : std_logic;
signal \N__45637\ : std_logic;
signal \N__45634\ : std_logic;
signal \N__45631\ : std_logic;
signal \N__45630\ : std_logic;
signal \N__45625\ : std_logic;
signal \N__45622\ : std_logic;
signal \N__45619\ : std_logic;
signal \N__45614\ : std_logic;
signal \N__45611\ : std_logic;
signal \N__45608\ : std_logic;
signal \N__45607\ : std_logic;
signal \N__45604\ : std_logic;
signal \N__45601\ : std_logic;
signal \N__45600\ : std_logic;
signal \N__45595\ : std_logic;
signal \N__45592\ : std_logic;
signal \N__45589\ : std_logic;
signal \N__45584\ : std_logic;
signal \N__45581\ : std_logic;
signal \N__45578\ : std_logic;
signal \N__45577\ : std_logic;
signal \N__45574\ : std_logic;
signal \N__45571\ : std_logic;
signal \N__45570\ : std_logic;
signal \N__45567\ : std_logic;
signal \N__45564\ : std_logic;
signal \N__45561\ : std_logic;
signal \N__45558\ : std_logic;
signal \N__45555\ : std_logic;
signal \N__45548\ : std_logic;
signal \N__45545\ : std_logic;
signal \N__45544\ : std_logic;
signal \N__45539\ : std_logic;
signal \N__45536\ : std_logic;
signal \N__45533\ : std_logic;
signal \N__45532\ : std_logic;
signal \N__45527\ : std_logic;
signal \N__45526\ : std_logic;
signal \N__45523\ : std_logic;
signal \N__45520\ : std_logic;
signal \N__45517\ : std_logic;
signal \N__45512\ : std_logic;
signal \N__45511\ : std_logic;
signal \N__45506\ : std_logic;
signal \N__45505\ : std_logic;
signal \N__45502\ : std_logic;
signal \N__45499\ : std_logic;
signal \N__45496\ : std_logic;
signal \N__45491\ : std_logic;
signal \N__45488\ : std_logic;
signal \N__45485\ : std_logic;
signal \N__45482\ : std_logic;
signal \N__45481\ : std_logic;
signal \N__45480\ : std_logic;
signal \N__45477\ : std_logic;
signal \N__45474\ : std_logic;
signal \N__45471\ : std_logic;
signal \N__45468\ : std_logic;
signal \N__45461\ : std_logic;
signal \N__45458\ : std_logic;
signal \N__45455\ : std_logic;
signal \N__45454\ : std_logic;
signal \N__45453\ : std_logic;
signal \N__45452\ : std_logic;
signal \N__45451\ : std_logic;
signal \N__45450\ : std_logic;
signal \N__45449\ : std_logic;
signal \N__45448\ : std_logic;
signal \N__45447\ : std_logic;
signal \N__45446\ : std_logic;
signal \N__45445\ : std_logic;
signal \N__45444\ : std_logic;
signal \N__45443\ : std_logic;
signal \N__45442\ : std_logic;
signal \N__45441\ : std_logic;
signal \N__45440\ : std_logic;
signal \N__45439\ : std_logic;
signal \N__45438\ : std_logic;
signal \N__45437\ : std_logic;
signal \N__45436\ : std_logic;
signal \N__45435\ : std_logic;
signal \N__45434\ : std_logic;
signal \N__45433\ : std_logic;
signal \N__45432\ : std_logic;
signal \N__45431\ : std_logic;
signal \N__45426\ : std_logic;
signal \N__45425\ : std_logic;
signal \N__45424\ : std_logic;
signal \N__45419\ : std_logic;
signal \N__45418\ : std_logic;
signal \N__45417\ : std_logic;
signal \N__45416\ : std_logic;
signal \N__45415\ : std_logic;
signal \N__45414\ : std_logic;
signal \N__45411\ : std_logic;
signal \N__45410\ : std_logic;
signal \N__45409\ : std_logic;
signal \N__45408\ : std_logic;
signal \N__45407\ : std_logic;
signal \N__45406\ : std_logic;
signal \N__45405\ : std_logic;
signal \N__45404\ : std_logic;
signal \N__45401\ : std_logic;
signal \N__45400\ : std_logic;
signal \N__45399\ : std_logic;
signal \N__45398\ : std_logic;
signal \N__45397\ : std_logic;
signal \N__45396\ : std_logic;
signal \N__45393\ : std_logic;
signal \N__45392\ : std_logic;
signal \N__45391\ : std_logic;
signal \N__45390\ : std_logic;
signal \N__45387\ : std_logic;
signal \N__45386\ : std_logic;
signal \N__45385\ : std_logic;
signal \N__45384\ : std_logic;
signal \N__45383\ : std_logic;
signal \N__45382\ : std_logic;
signal \N__45379\ : std_logic;
signal \N__45378\ : std_logic;
signal \N__45377\ : std_logic;
signal \N__45376\ : std_logic;
signal \N__45369\ : std_logic;
signal \N__45362\ : std_logic;
signal \N__45359\ : std_logic;
signal \N__45352\ : std_logic;
signal \N__45339\ : std_logic;
signal \N__45336\ : std_logic;
signal \N__45335\ : std_logic;
signal \N__45330\ : std_logic;
signal \N__45327\ : std_logic;
signal \N__45324\ : std_logic;
signal \N__45319\ : std_logic;
signal \N__45304\ : std_logic;
signal \N__45297\ : std_logic;
signal \N__45294\ : std_logic;
signal \N__45285\ : std_logic;
signal \N__45284\ : std_logic;
signal \N__45283\ : std_logic;
signal \N__45282\ : std_logic;
signal \N__45281\ : std_logic;
signal \N__45280\ : std_logic;
signal \N__45279\ : std_logic;
signal \N__45278\ : std_logic;
signal \N__45277\ : std_logic;
signal \N__45262\ : std_logic;
signal \N__45247\ : std_logic;
signal \N__45244\ : std_logic;
signal \N__45241\ : std_logic;
signal \N__45236\ : std_logic;
signal \N__45233\ : std_logic;
signal \N__45228\ : std_logic;
signal \N__45225\ : std_logic;
signal \N__45224\ : std_logic;
signal \N__45223\ : std_logic;
signal \N__45222\ : std_logic;
signal \N__45221\ : std_logic;
signal \N__45220\ : std_logic;
signal \N__45219\ : std_logic;
signal \N__45218\ : std_logic;
signal \N__45209\ : std_logic;
signal \N__45206\ : std_logic;
signal \N__45203\ : std_logic;
signal \N__45198\ : std_logic;
signal \N__45195\ : std_logic;
signal \N__45190\ : std_logic;
signal \N__45185\ : std_logic;
signal \N__45178\ : std_logic;
signal \N__45173\ : std_logic;
signal \N__45170\ : std_logic;
signal \N__45165\ : std_logic;
signal \N__45158\ : std_logic;
signal \N__45151\ : std_logic;
signal \N__45142\ : std_logic;
signal \N__45139\ : std_logic;
signal \N__45132\ : std_logic;
signal \N__45107\ : std_logic;
signal \N__45104\ : std_logic;
signal \N__45103\ : std_logic;
signal \N__45102\ : std_logic;
signal \N__45101\ : std_logic;
signal \N__45098\ : std_logic;
signal \N__45095\ : std_logic;
signal \N__45090\ : std_logic;
signal \N__45083\ : std_logic;
signal \N__45080\ : std_logic;
signal \N__45077\ : std_logic;
signal \N__45076\ : std_logic;
signal \N__45073\ : std_logic;
signal \N__45070\ : std_logic;
signal \N__45067\ : std_logic;
signal \N__45062\ : std_logic;
signal \N__45059\ : std_logic;
signal \N__45058\ : std_logic;
signal \N__45055\ : std_logic;
signal \N__45052\ : std_logic;
signal \N__45049\ : std_logic;
signal \N__45044\ : std_logic;
signal \N__45043\ : std_logic;
signal \N__45042\ : std_logic;
signal \N__45041\ : std_logic;
signal \N__45038\ : std_logic;
signal \N__45035\ : std_logic;
signal \N__45034\ : std_logic;
signal \N__45033\ : std_logic;
signal \N__45028\ : std_logic;
signal \N__45023\ : std_logic;
signal \N__45020\ : std_logic;
signal \N__45017\ : std_logic;
signal \N__45014\ : std_logic;
signal \N__45011\ : std_logic;
signal \N__45002\ : std_logic;
signal \N__45001\ : std_logic;
signal \N__44998\ : std_logic;
signal \N__44997\ : std_logic;
signal \N__44994\ : std_logic;
signal \N__44991\ : std_logic;
signal \N__44988\ : std_logic;
signal \N__44985\ : std_logic;
signal \N__44982\ : std_logic;
signal \N__44979\ : std_logic;
signal \N__44976\ : std_logic;
signal \N__44971\ : std_logic;
signal \N__44966\ : std_logic;
signal \N__44963\ : std_logic;
signal \N__44960\ : std_logic;
signal \N__44959\ : std_logic;
signal \N__44958\ : std_logic;
signal \N__44957\ : std_logic;
signal \N__44956\ : std_logic;
signal \N__44955\ : std_logic;
signal \N__44954\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44936\ : std_logic;
signal \N__44933\ : std_logic;
signal \N__44930\ : std_logic;
signal \N__44929\ : std_logic;
signal \N__44928\ : std_logic;
signal \N__44923\ : std_logic;
signal \N__44920\ : std_logic;
signal \N__44917\ : std_logic;
signal \N__44916\ : std_logic;
signal \N__44915\ : std_logic;
signal \N__44914\ : std_logic;
signal \N__44913\ : std_logic;
signal \N__44912\ : std_logic;
signal \N__44911\ : std_logic;
signal \N__44910\ : std_logic;
signal \N__44909\ : std_logic;
signal \N__44908\ : std_logic;
signal \N__44907\ : std_logic;
signal \N__44906\ : std_logic;
signal \N__44905\ : std_logic;
signal \N__44904\ : std_logic;
signal \N__44903\ : std_logic;
signal \N__44902\ : std_logic;
signal \N__44901\ : std_logic;
signal \N__44900\ : std_logic;
signal \N__44899\ : std_logic;
signal \N__44898\ : std_logic;
signal \N__44893\ : std_logic;
signal \N__44884\ : std_logic;
signal \N__44873\ : std_logic;
signal \N__44866\ : std_logic;
signal \N__44865\ : std_logic;
signal \N__44864\ : std_logic;
signal \N__44863\ : std_logic;
signal \N__44860\ : std_logic;
signal \N__44849\ : std_logic;
signal \N__44846\ : std_logic;
signal \N__44837\ : std_logic;
signal \N__44834\ : std_logic;
signal \N__44829\ : std_logic;
signal \N__44816\ : std_logic;
signal \N__44813\ : std_logic;
signal \N__44812\ : std_logic;
signal \N__44811\ : std_logic;
signal \N__44808\ : std_logic;
signal \N__44805\ : std_logic;
signal \N__44802\ : std_logic;
signal \N__44799\ : std_logic;
signal \N__44794\ : std_logic;
signal \N__44789\ : std_logic;
signal \N__44786\ : std_logic;
signal \N__44783\ : std_logic;
signal \N__44780\ : std_logic;
signal \N__44777\ : std_logic;
signal \N__44776\ : std_logic;
signal \N__44775\ : std_logic;
signal \N__44774\ : std_logic;
signal \N__44771\ : std_logic;
signal \N__44768\ : std_logic;
signal \N__44763\ : std_logic;
signal \N__44760\ : std_logic;
signal \N__44757\ : std_logic;
signal \N__44754\ : std_logic;
signal \N__44751\ : std_logic;
signal \N__44746\ : std_logic;
signal \N__44741\ : std_logic;
signal \N__44738\ : std_logic;
signal \N__44735\ : std_logic;
signal \N__44732\ : std_logic;
signal \N__44731\ : std_logic;
signal \N__44728\ : std_logic;
signal \N__44725\ : std_logic;
signal \N__44724\ : std_logic;
signal \N__44721\ : std_logic;
signal \N__44718\ : std_logic;
signal \N__44715\ : std_logic;
signal \N__44712\ : std_logic;
signal \N__44705\ : std_logic;
signal \N__44702\ : std_logic;
signal \N__44699\ : std_logic;
signal \N__44696\ : std_logic;
signal \N__44693\ : std_logic;
signal \N__44692\ : std_logic;
signal \N__44689\ : std_logic;
signal \N__44686\ : std_logic;
signal \N__44681\ : std_logic;
signal \N__44680\ : std_logic;
signal \N__44677\ : std_logic;
signal \N__44674\ : std_logic;
signal \N__44671\ : std_logic;
signal \N__44666\ : std_logic;
signal \N__44663\ : std_logic;
signal \N__44660\ : std_logic;
signal \N__44659\ : std_logic;
signal \N__44654\ : std_logic;
signal \N__44653\ : std_logic;
signal \N__44650\ : std_logic;
signal \N__44647\ : std_logic;
signal \N__44644\ : std_logic;
signal \N__44639\ : std_logic;
signal \N__44636\ : std_logic;
signal \N__44633\ : std_logic;
signal \N__44630\ : std_logic;
signal \N__44627\ : std_logic;
signal \N__44624\ : std_logic;
signal \N__44623\ : std_logic;
signal \N__44620\ : std_logic;
signal \N__44615\ : std_logic;
signal \N__44614\ : std_logic;
signal \N__44611\ : std_logic;
signal \N__44608\ : std_logic;
signal \N__44605\ : std_logic;
signal \N__44600\ : std_logic;
signal \N__44597\ : std_logic;
signal \N__44596\ : std_logic;
signal \N__44593\ : std_logic;
signal \N__44590\ : std_logic;
signal \N__44589\ : std_logic;
signal \N__44584\ : std_logic;
signal \N__44581\ : std_logic;
signal \N__44578\ : std_logic;
signal \N__44573\ : std_logic;
signal \N__44570\ : std_logic;
signal \N__44567\ : std_logic;
signal \N__44564\ : std_logic;
signal \N__44561\ : std_logic;
signal \N__44558\ : std_logic;
signal \N__44555\ : std_logic;
signal \N__44552\ : std_logic;
signal \N__44549\ : std_logic;
signal \N__44548\ : std_logic;
signal \N__44547\ : std_logic;
signal \N__44542\ : std_logic;
signal \N__44539\ : std_logic;
signal \N__44536\ : std_logic;
signal \N__44531\ : std_logic;
signal \N__44528\ : std_logic;
signal \N__44527\ : std_logic;
signal \N__44526\ : std_logic;
signal \N__44521\ : std_logic;
signal \N__44518\ : std_logic;
signal \N__44515\ : std_logic;
signal \N__44510\ : std_logic;
signal \N__44507\ : std_logic;
signal \N__44506\ : std_logic;
signal \N__44503\ : std_logic;
signal \N__44502\ : std_logic;
signal \N__44497\ : std_logic;
signal \N__44494\ : std_logic;
signal \N__44491\ : std_logic;
signal \N__44486\ : std_logic;
signal \N__44483\ : std_logic;
signal \N__44480\ : std_logic;
signal \N__44479\ : std_logic;
signal \N__44478\ : std_logic;
signal \N__44475\ : std_logic;
signal \N__44472\ : std_logic;
signal \N__44469\ : std_logic;
signal \N__44464\ : std_logic;
signal \N__44459\ : std_logic;
signal \N__44456\ : std_logic;
signal \N__44453\ : std_logic;
signal \N__44450\ : std_logic;
signal \N__44449\ : std_logic;
signal \N__44448\ : std_logic;
signal \N__44445\ : std_logic;
signal \N__44440\ : std_logic;
signal \N__44435\ : std_logic;
signal \N__44432\ : std_logic;
signal \N__44431\ : std_logic;
signal \N__44430\ : std_logic;
signal \N__44427\ : std_logic;
signal \N__44424\ : std_logic;
signal \N__44419\ : std_logic;
signal \N__44414\ : std_logic;
signal \N__44411\ : std_logic;
signal \N__44408\ : std_logic;
signal \N__44407\ : std_logic;
signal \N__44404\ : std_logic;
signal \N__44401\ : std_logic;
signal \N__44396\ : std_logic;
signal \N__44393\ : std_logic;
signal \N__44392\ : std_logic;
signal \N__44389\ : std_logic;
signal \N__44386\ : std_logic;
signal \N__44381\ : std_logic;
signal \N__44378\ : std_logic;
signal \N__44375\ : std_logic;
signal \N__44374\ : std_logic;
signal \N__44371\ : std_logic;
signal \N__44368\ : std_logic;
signal \N__44365\ : std_logic;
signal \N__44360\ : std_logic;
signal \N__44357\ : std_logic;
signal \N__44356\ : std_logic;
signal \N__44353\ : std_logic;
signal \N__44350\ : std_logic;
signal \N__44345\ : std_logic;
signal \N__44342\ : std_logic;
signal \N__44341\ : std_logic;
signal \N__44338\ : std_logic;
signal \N__44335\ : std_logic;
signal \N__44330\ : std_logic;
signal \N__44327\ : std_logic;
signal \N__44326\ : std_logic;
signal \N__44323\ : std_logic;
signal \N__44320\ : std_logic;
signal \N__44315\ : std_logic;
signal \N__44312\ : std_logic;
signal \N__44309\ : std_logic;
signal \N__44306\ : std_logic;
signal \N__44303\ : std_logic;
signal \N__44300\ : std_logic;
signal \N__44297\ : std_logic;
signal \N__44296\ : std_logic;
signal \N__44293\ : std_logic;
signal \N__44292\ : std_logic;
signal \N__44289\ : std_logic;
signal \N__44286\ : std_logic;
signal \N__44283\ : std_logic;
signal \N__44280\ : std_logic;
signal \N__44277\ : std_logic;
signal \N__44274\ : std_logic;
signal \N__44267\ : std_logic;
signal \N__44266\ : std_logic;
signal \N__44263\ : std_logic;
signal \N__44260\ : std_logic;
signal \N__44255\ : std_logic;
signal \N__44252\ : std_logic;
signal \N__44249\ : std_logic;
signal \N__44246\ : std_logic;
signal \N__44243\ : std_logic;
signal \N__44242\ : std_logic;
signal \N__44239\ : std_logic;
signal \N__44236\ : std_logic;
signal \N__44231\ : std_logic;
signal \N__44228\ : std_logic;
signal \N__44227\ : std_logic;
signal \N__44224\ : std_logic;
signal \N__44221\ : std_logic;
signal \N__44216\ : std_logic;
signal \N__44213\ : std_logic;
signal \N__44212\ : std_logic;
signal \N__44209\ : std_logic;
signal \N__44206\ : std_logic;
signal \N__44201\ : std_logic;
signal \N__44198\ : std_logic;
signal \N__44197\ : std_logic;
signal \N__44194\ : std_logic;
signal \N__44191\ : std_logic;
signal \N__44186\ : std_logic;
signal \N__44183\ : std_logic;
signal \N__44182\ : std_logic;
signal \N__44179\ : std_logic;
signal \N__44176\ : std_logic;
signal \N__44171\ : std_logic;
signal \N__44168\ : std_logic;
signal \N__44167\ : std_logic;
signal \N__44164\ : std_logic;
signal \N__44161\ : std_logic;
signal \N__44156\ : std_logic;
signal \N__44153\ : std_logic;
signal \N__44152\ : std_logic;
signal \N__44149\ : std_logic;
signal \N__44146\ : std_logic;
signal \N__44141\ : std_logic;
signal \N__44138\ : std_logic;
signal \N__44135\ : std_logic;
signal \N__44132\ : std_logic;
signal \N__44129\ : std_logic;
signal \N__44126\ : std_logic;
signal \N__44123\ : std_logic;
signal \N__44120\ : std_logic;
signal \N__44119\ : std_logic;
signal \N__44116\ : std_logic;
signal \N__44113\ : std_logic;
signal \N__44108\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44104\ : std_logic;
signal \N__44103\ : std_logic;
signal \N__44100\ : std_logic;
signal \N__44095\ : std_logic;
signal \N__44094\ : std_logic;
signal \N__44091\ : std_logic;
signal \N__44088\ : std_logic;
signal \N__44085\ : std_logic;
signal \N__44080\ : std_logic;
signal \N__44077\ : std_logic;
signal \N__44072\ : std_logic;
signal \N__44071\ : std_logic;
signal \N__44068\ : std_logic;
signal \N__44063\ : std_logic;
signal \N__44060\ : std_logic;
signal \N__44059\ : std_logic;
signal \N__44056\ : std_logic;
signal \N__44055\ : std_logic;
signal \N__44052\ : std_logic;
signal \N__44049\ : std_logic;
signal \N__44046\ : std_logic;
signal \N__44039\ : std_logic;
signal \N__44036\ : std_logic;
signal \N__44035\ : std_logic;
signal \N__44032\ : std_logic;
signal \N__44029\ : std_logic;
signal \N__44028\ : std_logic;
signal \N__44027\ : std_logic;
signal \N__44022\ : std_logic;
signal \N__44017\ : std_logic;
signal \N__44012\ : std_logic;
signal \N__44009\ : std_logic;
signal \N__44006\ : std_logic;
signal \N__44003\ : std_logic;
signal \N__44002\ : std_logic;
signal \N__43997\ : std_logic;
signal \N__43994\ : std_logic;
signal \N__43991\ : std_logic;
signal \N__43988\ : std_logic;
signal \N__43985\ : std_logic;
signal \N__43984\ : std_logic;
signal \N__43981\ : std_logic;
signal \N__43978\ : std_logic;
signal \N__43973\ : std_logic;
signal \N__43972\ : std_logic;
signal \N__43967\ : std_logic;
signal \N__43964\ : std_logic;
signal \N__43963\ : std_logic;
signal \N__43960\ : std_logic;
signal \N__43957\ : std_logic;
signal \N__43952\ : std_logic;
signal \N__43949\ : std_logic;
signal \N__43946\ : std_logic;
signal \N__43943\ : std_logic;
signal \N__43940\ : std_logic;
signal \N__43939\ : std_logic;
signal \N__43938\ : std_logic;
signal \N__43935\ : std_logic;
signal \N__43932\ : std_logic;
signal \N__43929\ : std_logic;
signal \N__43926\ : std_logic;
signal \N__43923\ : std_logic;
signal \N__43920\ : std_logic;
signal \N__43919\ : std_logic;
signal \N__43916\ : std_logic;
signal \N__43913\ : std_logic;
signal \N__43910\ : std_logic;
signal \N__43907\ : std_logic;
signal \N__43904\ : std_logic;
signal \N__43901\ : std_logic;
signal \N__43898\ : std_logic;
signal \N__43889\ : std_logic;
signal \N__43886\ : std_logic;
signal \N__43885\ : std_logic;
signal \N__43882\ : std_logic;
signal \N__43881\ : std_logic;
signal \N__43878\ : std_logic;
signal \N__43875\ : std_logic;
signal \N__43872\ : std_logic;
signal \N__43865\ : std_logic;
signal \N__43862\ : std_logic;
signal \N__43861\ : std_logic;
signal \N__43858\ : std_logic;
signal \N__43855\ : std_logic;
signal \N__43854\ : std_logic;
signal \N__43851\ : std_logic;
signal \N__43848\ : std_logic;
signal \N__43845\ : std_logic;
signal \N__43838\ : std_logic;
signal \N__43837\ : std_logic;
signal \N__43834\ : std_logic;
signal \N__43831\ : std_logic;
signal \N__43828\ : std_logic;
signal \N__43825\ : std_logic;
signal \N__43824\ : std_logic;
signal \N__43821\ : std_logic;
signal \N__43818\ : std_logic;
signal \N__43815\ : std_logic;
signal \N__43812\ : std_logic;
signal \N__43805\ : std_logic;
signal \N__43802\ : std_logic;
signal \N__43801\ : std_logic;
signal \N__43800\ : std_logic;
signal \N__43797\ : std_logic;
signal \N__43794\ : std_logic;
signal \N__43793\ : std_logic;
signal \N__43792\ : std_logic;
signal \N__43789\ : std_logic;
signal \N__43784\ : std_logic;
signal \N__43781\ : std_logic;
signal \N__43778\ : std_logic;
signal \N__43775\ : std_logic;
signal \N__43772\ : std_logic;
signal \N__43769\ : std_logic;
signal \N__43766\ : std_logic;
signal \N__43763\ : std_logic;
signal \N__43758\ : std_logic;
signal \N__43755\ : std_logic;
signal \N__43748\ : std_logic;
signal \N__43745\ : std_logic;
signal \N__43744\ : std_logic;
signal \N__43741\ : std_logic;
signal \N__43740\ : std_logic;
signal \N__43737\ : std_logic;
signal \N__43734\ : std_logic;
signal \N__43731\ : std_logic;
signal \N__43724\ : std_logic;
signal \N__43721\ : std_logic;
signal \N__43720\ : std_logic;
signal \N__43717\ : std_logic;
signal \N__43716\ : std_logic;
signal \N__43713\ : std_logic;
signal \N__43710\ : std_logic;
signal \N__43707\ : std_logic;
signal \N__43700\ : std_logic;
signal \N__43697\ : std_logic;
signal \N__43696\ : std_logic;
signal \N__43693\ : std_logic;
signal \N__43692\ : std_logic;
signal \N__43689\ : std_logic;
signal \N__43686\ : std_logic;
signal \N__43683\ : std_logic;
signal \N__43676\ : std_logic;
signal \N__43673\ : std_logic;
signal \N__43670\ : std_logic;
signal \N__43667\ : std_logic;
signal \N__43664\ : std_logic;
signal \N__43661\ : std_logic;
signal \N__43658\ : std_logic;
signal \N__43655\ : std_logic;
signal \N__43652\ : std_logic;
signal \N__43649\ : std_logic;
signal \N__43646\ : std_logic;
signal \N__43643\ : std_logic;
signal \N__43640\ : std_logic;
signal \N__43637\ : std_logic;
signal \N__43634\ : std_logic;
signal \N__43631\ : std_logic;
signal \N__43628\ : std_logic;
signal \N__43625\ : std_logic;
signal \N__43622\ : std_logic;
signal \N__43619\ : std_logic;
signal \N__43616\ : std_logic;
signal \N__43613\ : std_logic;
signal \N__43610\ : std_logic;
signal \N__43607\ : std_logic;
signal \N__43604\ : std_logic;
signal \N__43601\ : std_logic;
signal \N__43598\ : std_logic;
signal \N__43595\ : std_logic;
signal \N__43592\ : std_logic;
signal \N__43591\ : std_logic;
signal \N__43590\ : std_logic;
signal \N__43589\ : std_logic;
signal \N__43586\ : std_logic;
signal \N__43583\ : std_logic;
signal \N__43582\ : std_logic;
signal \N__43581\ : std_logic;
signal \N__43580\ : std_logic;
signal \N__43579\ : std_logic;
signal \N__43578\ : std_logic;
signal \N__43577\ : std_logic;
signal \N__43576\ : std_logic;
signal \N__43575\ : std_logic;
signal \N__43574\ : std_logic;
signal \N__43573\ : std_logic;
signal \N__43572\ : std_logic;
signal \N__43571\ : std_logic;
signal \N__43568\ : std_logic;
signal \N__43567\ : std_logic;
signal \N__43566\ : std_logic;
signal \N__43563\ : std_logic;
signal \N__43562\ : std_logic;
signal \N__43561\ : std_logic;
signal \N__43560\ : std_logic;
signal \N__43559\ : std_logic;
signal \N__43558\ : std_logic;
signal \N__43557\ : std_logic;
signal \N__43556\ : std_logic;
signal \N__43555\ : std_logic;
signal \N__43554\ : std_logic;
signal \N__43553\ : std_logic;
signal \N__43552\ : std_logic;
signal \N__43551\ : std_logic;
signal \N__43546\ : std_logic;
signal \N__43543\ : std_logic;
signal \N__43532\ : std_logic;
signal \N__43529\ : std_logic;
signal \N__43520\ : std_logic;
signal \N__43517\ : std_logic;
signal \N__43516\ : std_logic;
signal \N__43515\ : std_logic;
signal \N__43512\ : std_logic;
signal \N__43501\ : std_logic;
signal \N__43496\ : std_logic;
signal \N__43491\ : std_logic;
signal \N__43488\ : std_logic;
signal \N__43477\ : std_logic;
signal \N__43466\ : std_logic;
signal \N__43463\ : std_logic;
signal \N__43458\ : std_logic;
signal \N__43451\ : std_logic;
signal \N__43442\ : std_logic;
signal \N__43439\ : std_logic;
signal \N__43436\ : std_logic;
signal \N__43433\ : std_logic;
signal \N__43430\ : std_logic;
signal \N__43427\ : std_logic;
signal \N__43424\ : std_logic;
signal \N__43419\ : std_logic;
signal \N__43412\ : std_logic;
signal \N__43409\ : std_logic;
signal \N__43406\ : std_logic;
signal \N__43403\ : std_logic;
signal \N__43400\ : std_logic;
signal \N__43397\ : std_logic;
signal \N__43394\ : std_logic;
signal \N__43391\ : std_logic;
signal \N__43388\ : std_logic;
signal \N__43385\ : std_logic;
signal \N__43382\ : std_logic;
signal \N__43379\ : std_logic;
signal \N__43376\ : std_logic;
signal \N__43373\ : std_logic;
signal \N__43370\ : std_logic;
signal \N__43367\ : std_logic;
signal \N__43364\ : std_logic;
signal \N__43361\ : std_logic;
signal \N__43358\ : std_logic;
signal \N__43355\ : std_logic;
signal \N__43352\ : std_logic;
signal \N__43349\ : std_logic;
signal \N__43346\ : std_logic;
signal \N__43343\ : std_logic;
signal \N__43340\ : std_logic;
signal \N__43337\ : std_logic;
signal \N__43334\ : std_logic;
signal \N__43331\ : std_logic;
signal \N__43328\ : std_logic;
signal \N__43325\ : std_logic;
signal \N__43322\ : std_logic;
signal \N__43319\ : std_logic;
signal \N__43316\ : std_logic;
signal \N__43313\ : std_logic;
signal \N__43310\ : std_logic;
signal \N__43307\ : std_logic;
signal \N__43304\ : std_logic;
signal \N__43301\ : std_logic;
signal \N__43298\ : std_logic;
signal \N__43295\ : std_logic;
signal \N__43292\ : std_logic;
signal \N__43289\ : std_logic;
signal \N__43286\ : std_logic;
signal \N__43283\ : std_logic;
signal \N__43280\ : std_logic;
signal \N__43277\ : std_logic;
signal \N__43274\ : std_logic;
signal \N__43271\ : std_logic;
signal \N__43268\ : std_logic;
signal \N__43265\ : std_logic;
signal \N__43262\ : std_logic;
signal \N__43259\ : std_logic;
signal \N__43256\ : std_logic;
signal \N__43253\ : std_logic;
signal \N__43250\ : std_logic;
signal \N__43247\ : std_logic;
signal \N__43244\ : std_logic;
signal \N__43241\ : std_logic;
signal \N__43238\ : std_logic;
signal \N__43235\ : std_logic;
signal \N__43232\ : std_logic;
signal \N__43229\ : std_logic;
signal \N__43226\ : std_logic;
signal \N__43223\ : std_logic;
signal \N__43220\ : std_logic;
signal \N__43217\ : std_logic;
signal \N__43214\ : std_logic;
signal \N__43211\ : std_logic;
signal \N__43208\ : std_logic;
signal \N__43205\ : std_logic;
signal \N__43202\ : std_logic;
signal \N__43199\ : std_logic;
signal \N__43196\ : std_logic;
signal \N__43193\ : std_logic;
signal \N__43190\ : std_logic;
signal \N__43187\ : std_logic;
signal \N__43184\ : std_logic;
signal \N__43181\ : std_logic;
signal \N__43178\ : std_logic;
signal \N__43175\ : std_logic;
signal \N__43172\ : std_logic;
signal \N__43169\ : std_logic;
signal \N__43166\ : std_logic;
signal \N__43163\ : std_logic;
signal \N__43160\ : std_logic;
signal \N__43157\ : std_logic;
signal \N__43154\ : std_logic;
signal \N__43151\ : std_logic;
signal \N__43148\ : std_logic;
signal \N__43145\ : std_logic;
signal \N__43142\ : std_logic;
signal \N__43139\ : std_logic;
signal \N__43138\ : std_logic;
signal \N__43137\ : std_logic;
signal \N__43136\ : std_logic;
signal \N__43133\ : std_logic;
signal \N__43130\ : std_logic;
signal \N__43125\ : std_logic;
signal \N__43122\ : std_logic;
signal \N__43119\ : std_logic;
signal \N__43116\ : std_logic;
signal \N__43113\ : std_logic;
signal \N__43108\ : std_logic;
signal \N__43105\ : std_logic;
signal \N__43102\ : std_logic;
signal \N__43097\ : std_logic;
signal \N__43094\ : std_logic;
signal \N__43091\ : std_logic;
signal \N__43090\ : std_logic;
signal \N__43089\ : std_logic;
signal \N__43086\ : std_logic;
signal \N__43083\ : std_logic;
signal \N__43080\ : std_logic;
signal \N__43073\ : std_logic;
signal \N__43070\ : std_logic;
signal \N__43069\ : std_logic;
signal \N__43068\ : std_logic;
signal \N__43065\ : std_logic;
signal \N__43062\ : std_logic;
signal \N__43059\ : std_logic;
signal \N__43056\ : std_logic;
signal \N__43055\ : std_logic;
signal \N__43050\ : std_logic;
signal \N__43047\ : std_logic;
signal \N__43044\ : std_logic;
signal \N__43041\ : std_logic;
signal \N__43034\ : std_logic;
signal \N__43033\ : std_logic;
signal \N__43030\ : std_logic;
signal \N__43029\ : std_logic;
signal \N__43026\ : std_logic;
signal \N__43023\ : std_logic;
signal \N__43020\ : std_logic;
signal \N__43017\ : std_logic;
signal \N__43014\ : std_logic;
signal \N__43011\ : std_logic;
signal \N__43008\ : std_logic;
signal \N__43001\ : std_logic;
signal \N__43000\ : std_logic;
signal \N__42997\ : std_logic;
signal \N__42996\ : std_logic;
signal \N__42993\ : std_logic;
signal \N__42990\ : std_logic;
signal \N__42987\ : std_logic;
signal \N__42984\ : std_logic;
signal \N__42981\ : std_logic;
signal \N__42978\ : std_logic;
signal \N__42975\ : std_logic;
signal \N__42968\ : std_logic;
signal \N__42965\ : std_logic;
signal \N__42962\ : std_logic;
signal \N__42959\ : std_logic;
signal \N__42956\ : std_logic;
signal \N__42953\ : std_logic;
signal \N__42952\ : std_logic;
signal \N__42949\ : std_logic;
signal \N__42948\ : std_logic;
signal \N__42945\ : std_logic;
signal \N__42940\ : std_logic;
signal \N__42935\ : std_logic;
signal \N__42934\ : std_logic;
signal \N__42931\ : std_logic;
signal \N__42928\ : std_logic;
signal \N__42923\ : std_logic;
signal \N__42920\ : std_logic;
signal \N__42917\ : std_logic;
signal \N__42914\ : std_logic;
signal \N__42911\ : std_logic;
signal \N__42910\ : std_logic;
signal \N__42909\ : std_logic;
signal \N__42908\ : std_logic;
signal \N__42907\ : std_logic;
signal \N__42906\ : std_logic;
signal \N__42903\ : std_logic;
signal \N__42902\ : std_logic;
signal \N__42899\ : std_logic;
signal \N__42898\ : std_logic;
signal \N__42897\ : std_logic;
signal \N__42896\ : std_logic;
signal \N__42895\ : std_logic;
signal \N__42894\ : std_logic;
signal \N__42893\ : std_logic;
signal \N__42892\ : std_logic;
signal \N__42891\ : std_logic;
signal \N__42890\ : std_logic;
signal \N__42889\ : std_logic;
signal \N__42888\ : std_logic;
signal \N__42887\ : std_logic;
signal \N__42884\ : std_logic;
signal \N__42883\ : std_logic;
signal \N__42882\ : std_logic;
signal \N__42881\ : std_logic;
signal \N__42880\ : std_logic;
signal \N__42879\ : std_logic;
signal \N__42878\ : std_logic;
signal \N__42877\ : std_logic;
signal \N__42876\ : std_logic;
signal \N__42871\ : std_logic;
signal \N__42866\ : std_logic;
signal \N__42865\ : std_logic;
signal \N__42864\ : std_logic;
signal \N__42863\ : std_logic;
signal \N__42862\ : std_logic;
signal \N__42861\ : std_logic;
signal \N__42860\ : std_logic;
signal \N__42859\ : std_logic;
signal \N__42858\ : std_logic;
signal \N__42857\ : std_logic;
signal \N__42856\ : std_logic;
signal \N__42855\ : std_logic;
signal \N__42854\ : std_logic;
signal \N__42851\ : std_logic;
signal \N__42848\ : std_logic;
signal \N__42847\ : std_logic;
signal \N__42846\ : std_logic;
signal \N__42843\ : std_logic;
signal \N__42842\ : std_logic;
signal \N__42841\ : std_logic;
signal \N__42840\ : std_logic;
signal \N__42839\ : std_logic;
signal \N__42838\ : std_logic;
signal \N__42837\ : std_logic;
signal \N__42834\ : std_logic;
signal \N__42833\ : std_logic;
signal \N__42832\ : std_logic;
signal \N__42831\ : std_logic;
signal \N__42828\ : std_logic;
signal \N__42827\ : std_logic;
signal \N__42826\ : std_logic;
signal \N__42825\ : std_logic;
signal \N__42824\ : std_logic;
signal \N__42823\ : std_logic;
signal \N__42820\ : std_logic;
signal \N__42819\ : std_logic;
signal \N__42816\ : std_logic;
signal \N__42815\ : std_logic;
signal \N__42812\ : std_logic;
signal \N__42809\ : std_logic;
signal \N__42808\ : std_logic;
signal \N__42805\ : std_logic;
signal \N__42804\ : std_logic;
signal \N__42801\ : std_logic;
signal \N__42800\ : std_logic;
signal \N__42797\ : std_logic;
signal \N__42796\ : std_logic;
signal \N__42795\ : std_logic;
signal \N__42794\ : std_logic;
signal \N__42793\ : std_logic;
signal \N__42792\ : std_logic;
signal \N__42789\ : std_logic;
signal \N__42788\ : std_logic;
signal \N__42787\ : std_logic;
signal \N__42786\ : std_logic;
signal \N__42785\ : std_logic;
signal \N__42784\ : std_logic;
signal \N__42783\ : std_logic;
signal \N__42782\ : std_logic;
signal \N__42781\ : std_logic;
signal \N__42780\ : std_logic;
signal \N__42779\ : std_logic;
signal \N__42778\ : std_logic;
signal \N__42773\ : std_logic;
signal \N__42772\ : std_logic;
signal \N__42771\ : std_logic;
signal \N__42768\ : std_logic;
signal \N__42765\ : std_logic;
signal \N__42762\ : std_logic;
signal \N__42757\ : std_logic;
signal \N__42754\ : std_logic;
signal \N__42753\ : std_logic;
signal \N__42750\ : std_logic;
signal \N__42749\ : std_logic;
signal \N__42746\ : std_logic;
signal \N__42745\ : std_logic;
signal \N__42740\ : std_logic;
signal \N__42737\ : std_logic;
signal \N__42734\ : std_logic;
signal \N__42731\ : std_logic;
signal \N__42730\ : std_logic;
signal \N__42727\ : std_logic;
signal \N__42724\ : std_logic;
signal \N__42723\ : std_logic;
signal \N__42722\ : std_logic;
signal \N__42721\ : std_logic;
signal \N__42720\ : std_logic;
signal \N__42719\ : std_logic;
signal \N__42718\ : std_logic;
signal \N__42717\ : std_logic;
signal \N__42716\ : std_logic;
signal \N__42713\ : std_logic;
signal \N__42710\ : std_logic;
signal \N__42697\ : std_logic;
signal \N__42694\ : std_logic;
signal \N__42689\ : std_logic;
signal \N__42674\ : std_logic;
signal \N__42659\ : std_logic;
signal \N__42656\ : std_logic;
signal \N__42641\ : std_logic;
signal \N__42624\ : std_logic;
signal \N__42621\ : std_logic;
signal \N__42620\ : std_logic;
signal \N__42617\ : std_logic;
signal \N__42616\ : std_logic;
signal \N__42613\ : std_logic;
signal \N__42612\ : std_logic;
signal \N__42609\ : std_logic;
signal \N__42608\ : std_logic;
signal \N__42607\ : std_logic;
signal \N__42606\ : std_logic;
signal \N__42605\ : std_logic;
signal \N__42602\ : std_logic;
signal \N__42595\ : std_logic;
signal \N__42592\ : std_logic;
signal \N__42591\ : std_logic;
signal \N__42588\ : std_logic;
signal \N__42587\ : std_logic;
signal \N__42584\ : std_logic;
signal \N__42583\ : std_logic;
signal \N__42580\ : std_logic;
signal \N__42579\ : std_logic;
signal \N__42576\ : std_logic;
signal \N__42575\ : std_logic;
signal \N__42572\ : std_logic;
signal \N__42571\ : std_logic;
signal \N__42568\ : std_logic;
signal \N__42567\ : std_logic;
signal \N__42564\ : std_logic;
signal \N__42563\ : std_logic;
signal \N__42560\ : std_logic;
signal \N__42553\ : std_logic;
signal \N__42550\ : std_logic;
signal \N__42545\ : std_logic;
signal \N__42532\ : std_logic;
signal \N__42529\ : std_logic;
signal \N__42524\ : std_logic;
signal \N__42513\ : std_logic;
signal \N__42512\ : std_logic;
signal \N__42511\ : std_logic;
signal \N__42508\ : std_logic;
signal \N__42505\ : std_logic;
signal \N__42504\ : std_logic;
signal \N__42503\ : std_logic;
signal \N__42502\ : std_logic;
signal \N__42499\ : std_logic;
signal \N__42498\ : std_logic;
signal \N__42495\ : std_logic;
signal \N__42494\ : std_logic;
signal \N__42491\ : std_logic;
signal \N__42490\ : std_logic;
signal \N__42487\ : std_logic;
signal \N__42486\ : std_logic;
signal \N__42483\ : std_logic;
signal \N__42482\ : std_logic;
signal \N__42475\ : std_logic;
signal \N__42460\ : std_logic;
signal \N__42443\ : std_logic;
signal \N__42440\ : std_logic;
signal \N__42439\ : std_logic;
signal \N__42436\ : std_logic;
signal \N__42435\ : std_logic;
signal \N__42432\ : std_logic;
signal \N__42431\ : std_logic;
signal \N__42426\ : std_logic;
signal \N__42423\ : std_logic;
signal \N__42408\ : std_logic;
signal \N__42391\ : std_logic;
signal \N__42380\ : std_logic;
signal \N__42377\ : std_logic;
signal \N__42372\ : std_logic;
signal \N__42359\ : std_logic;
signal \N__42352\ : std_logic;
signal \N__42335\ : std_logic;
signal \N__42328\ : std_logic;
signal \N__42315\ : std_logic;
signal \N__42304\ : std_logic;
signal \N__42287\ : std_logic;
signal \N__42286\ : std_logic;
signal \N__42285\ : std_logic;
signal \N__42282\ : std_logic;
signal \N__42279\ : std_logic;
signal \N__42276\ : std_logic;
signal \N__42273\ : std_logic;
signal \N__42270\ : std_logic;
signal \N__42263\ : std_logic;
signal \N__42260\ : std_logic;
signal \N__42257\ : std_logic;
signal \N__42256\ : std_logic;
signal \N__42255\ : std_logic;
signal \N__42252\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42246\ : std_logic;
signal \N__42245\ : std_logic;
signal \N__42242\ : std_logic;
signal \N__42239\ : std_logic;
signal \N__42236\ : std_logic;
signal \N__42233\ : std_logic;
signal \N__42224\ : std_logic;
signal \N__42221\ : std_logic;
signal \N__42218\ : std_logic;
signal \N__42215\ : std_logic;
signal \N__42212\ : std_logic;
signal \N__42209\ : std_logic;
signal \N__42208\ : std_logic;
signal \N__42205\ : std_logic;
signal \N__42202\ : std_logic;
signal \N__42199\ : std_logic;
signal \N__42198\ : std_logic;
signal \N__42195\ : std_logic;
signal \N__42192\ : std_logic;
signal \N__42189\ : std_logic;
signal \N__42188\ : std_logic;
signal \N__42185\ : std_logic;
signal \N__42180\ : std_logic;
signal \N__42177\ : std_logic;
signal \N__42170\ : std_logic;
signal \N__42169\ : std_logic;
signal \N__42166\ : std_logic;
signal \N__42163\ : std_logic;
signal \N__42162\ : std_logic;
signal \N__42159\ : std_logic;
signal \N__42156\ : std_logic;
signal \N__42153\ : std_logic;
signal \N__42146\ : std_logic;
signal \N__42145\ : std_logic;
signal \N__42142\ : std_logic;
signal \N__42139\ : std_logic;
signal \N__42136\ : std_logic;
signal \N__42133\ : std_logic;
signal \N__42132\ : std_logic;
signal \N__42131\ : std_logic;
signal \N__42126\ : std_logic;
signal \N__42123\ : std_logic;
signal \N__42120\ : std_logic;
signal \N__42113\ : std_logic;
signal \N__42110\ : std_logic;
signal \N__42109\ : std_logic;
signal \N__42108\ : std_logic;
signal \N__42105\ : std_logic;
signal \N__42102\ : std_logic;
signal \N__42099\ : std_logic;
signal \N__42094\ : std_logic;
signal \N__42091\ : std_logic;
signal \N__42086\ : std_logic;
signal \N__42083\ : std_logic;
signal \N__42080\ : std_logic;
signal \N__42077\ : std_logic;
signal \N__42076\ : std_logic;
signal \N__42075\ : std_logic;
signal \N__42072\ : std_logic;
signal \N__42069\ : std_logic;
signal \N__42066\ : std_logic;
signal \N__42065\ : std_logic;
signal \N__42060\ : std_logic;
signal \N__42057\ : std_logic;
signal \N__42054\ : std_logic;
signal \N__42047\ : std_logic;
signal \N__42044\ : std_logic;
signal \N__42041\ : std_logic;
signal \N__42038\ : std_logic;
signal \N__42035\ : std_logic;
signal \N__42034\ : std_logic;
signal \N__42031\ : std_logic;
signal \N__42028\ : std_logic;
signal \N__42023\ : std_logic;
signal \N__42022\ : std_logic;
signal \N__42021\ : std_logic;
signal \N__42018\ : std_logic;
signal \N__42015\ : std_logic;
signal \N__42012\ : std_logic;
signal \N__42007\ : std_logic;
signal \N__42004\ : std_logic;
signal \N__41999\ : std_logic;
signal \N__41998\ : std_logic;
signal \N__41993\ : std_logic;
signal \N__41992\ : std_logic;
signal \N__41989\ : std_logic;
signal \N__41986\ : std_logic;
signal \N__41981\ : std_logic;
signal \N__41978\ : std_logic;
signal \N__41975\ : std_logic;
signal \N__41974\ : std_logic;
signal \N__41971\ : std_logic;
signal \N__41968\ : std_logic;
signal \N__41965\ : std_logic;
signal \N__41962\ : std_logic;
signal \N__41959\ : std_logic;
signal \N__41958\ : std_logic;
signal \N__41955\ : std_logic;
signal \N__41952\ : std_logic;
signal \N__41949\ : std_logic;
signal \N__41948\ : std_logic;
signal \N__41945\ : std_logic;
signal \N__41942\ : std_logic;
signal \N__41939\ : std_logic;
signal \N__41936\ : std_logic;
signal \N__41927\ : std_logic;
signal \N__41926\ : std_logic;
signal \N__41923\ : std_logic;
signal \N__41920\ : std_logic;
signal \N__41917\ : std_logic;
signal \N__41916\ : std_logic;
signal \N__41911\ : std_logic;
signal \N__41908\ : std_logic;
signal \N__41903\ : std_logic;
signal \N__41900\ : std_logic;
signal \N__41897\ : std_logic;
signal \N__41896\ : std_logic;
signal \N__41895\ : std_logic;
signal \N__41892\ : std_logic;
signal \N__41889\ : std_logic;
signal \N__41886\ : std_logic;
signal \N__41885\ : std_logic;
signal \N__41880\ : std_logic;
signal \N__41877\ : std_logic;
signal \N__41874\ : std_logic;
signal \N__41867\ : std_logic;
signal \N__41864\ : std_logic;
signal \N__41861\ : std_logic;
signal \N__41858\ : std_logic;
signal \N__41857\ : std_logic;
signal \N__41856\ : std_logic;
signal \N__41853\ : std_logic;
signal \N__41850\ : std_logic;
signal \N__41847\ : std_logic;
signal \N__41844\ : std_logic;
signal \N__41843\ : std_logic;
signal \N__41840\ : std_logic;
signal \N__41837\ : std_logic;
signal \N__41834\ : std_logic;
signal \N__41831\ : std_logic;
signal \N__41828\ : std_logic;
signal \N__41825\ : std_logic;
signal \N__41820\ : std_logic;
signal \N__41813\ : std_logic;
signal \N__41810\ : std_logic;
signal \N__41809\ : std_logic;
signal \N__41808\ : std_logic;
signal \N__41805\ : std_logic;
signal \N__41802\ : std_logic;
signal \N__41799\ : std_logic;
signal \N__41792\ : std_logic;
signal \N__41791\ : std_logic;
signal \N__41788\ : std_logic;
signal \N__41785\ : std_logic;
signal \N__41782\ : std_logic;
signal \N__41781\ : std_logic;
signal \N__41778\ : std_logic;
signal \N__41775\ : std_logic;
signal \N__41772\ : std_logic;
signal \N__41771\ : std_logic;
signal \N__41766\ : std_logic;
signal \N__41763\ : std_logic;
signal \N__41760\ : std_logic;
signal \N__41753\ : std_logic;
signal \N__41752\ : std_logic;
signal \N__41749\ : std_logic;
signal \N__41746\ : std_logic;
signal \N__41743\ : std_logic;
signal \N__41742\ : std_logic;
signal \N__41739\ : std_logic;
signal \N__41736\ : std_logic;
signal \N__41733\ : std_logic;
signal \N__41726\ : std_logic;
signal \N__41725\ : std_logic;
signal \N__41722\ : std_logic;
signal \N__41721\ : std_logic;
signal \N__41716\ : std_logic;
signal \N__41713\ : std_logic;
signal \N__41708\ : std_logic;
signal \N__41707\ : std_logic;
signal \N__41706\ : std_logic;
signal \N__41705\ : std_logic;
signal \N__41700\ : std_logic;
signal \N__41695\ : std_logic;
signal \N__41692\ : std_logic;
signal \N__41689\ : std_logic;
signal \N__41684\ : std_logic;
signal \N__41681\ : std_logic;
signal \N__41678\ : std_logic;
signal \N__41675\ : std_logic;
signal \N__41672\ : std_logic;
signal \N__41671\ : std_logic;
signal \N__41670\ : std_logic;
signal \N__41667\ : std_logic;
signal \N__41664\ : std_logic;
signal \N__41661\ : std_logic;
signal \N__41660\ : std_logic;
signal \N__41657\ : std_logic;
signal \N__41654\ : std_logic;
signal \N__41651\ : std_logic;
signal \N__41648\ : std_logic;
signal \N__41639\ : std_logic;
signal \N__41638\ : std_logic;
signal \N__41635\ : std_logic;
signal \N__41632\ : std_logic;
signal \N__41631\ : std_logic;
signal \N__41628\ : std_logic;
signal \N__41625\ : std_logic;
signal \N__41622\ : std_logic;
signal \N__41615\ : std_logic;
signal \N__41614\ : std_logic;
signal \N__41611\ : std_logic;
signal \N__41608\ : std_logic;
signal \N__41607\ : std_logic;
signal \N__41604\ : std_logic;
signal \N__41599\ : std_logic;
signal \N__41598\ : std_logic;
signal \N__41595\ : std_logic;
signal \N__41592\ : std_logic;
signal \N__41589\ : std_logic;
signal \N__41586\ : std_logic;
signal \N__41583\ : std_logic;
signal \N__41580\ : std_logic;
signal \N__41573\ : std_logic;
signal \N__41570\ : std_logic;
signal \N__41567\ : std_logic;
signal \N__41566\ : std_logic;
signal \N__41565\ : std_logic;
signal \N__41562\ : std_logic;
signal \N__41557\ : std_logic;
signal \N__41552\ : std_logic;
signal \N__41549\ : std_logic;
signal \N__41546\ : std_logic;
signal \N__41543\ : std_logic;
signal \N__41540\ : std_logic;
signal \N__41537\ : std_logic;
signal \N__41536\ : std_logic;
signal \N__41535\ : std_logic;
signal \N__41532\ : std_logic;
signal \N__41529\ : std_logic;
signal \N__41526\ : std_logic;
signal \N__41519\ : std_logic;
signal \N__41518\ : std_logic;
signal \N__41517\ : std_logic;
signal \N__41514\ : std_logic;
signal \N__41513\ : std_logic;
signal \N__41508\ : std_logic;
signal \N__41505\ : std_logic;
signal \N__41502\ : std_logic;
signal \N__41499\ : std_logic;
signal \N__41496\ : std_logic;
signal \N__41493\ : std_logic;
signal \N__41490\ : std_logic;
signal \N__41483\ : std_logic;
signal \N__41480\ : std_logic;
signal \N__41479\ : std_logic;
signal \N__41476\ : std_logic;
signal \N__41473\ : std_logic;
signal \N__41472\ : std_logic;
signal \N__41469\ : std_logic;
signal \N__41466\ : std_logic;
signal \N__41463\ : std_logic;
signal \N__41456\ : std_logic;
signal \N__41453\ : std_logic;
signal \N__41450\ : std_logic;
signal \N__41447\ : std_logic;
signal \N__41444\ : std_logic;
signal \N__41441\ : std_logic;
signal \N__41440\ : std_logic;
signal \N__41437\ : std_logic;
signal \N__41434\ : std_logic;
signal \N__41431\ : std_logic;
signal \N__41428\ : std_logic;
signal \N__41427\ : std_logic;
signal \N__41422\ : std_logic;
signal \N__41419\ : std_logic;
signal \N__41418\ : std_logic;
signal \N__41413\ : std_logic;
signal \N__41410\ : std_logic;
signal \N__41405\ : std_logic;
signal \N__41402\ : std_logic;
signal \N__41401\ : std_logic;
signal \N__41398\ : std_logic;
signal \N__41397\ : std_logic;
signal \N__41394\ : std_logic;
signal \N__41391\ : std_logic;
signal \N__41388\ : std_logic;
signal \N__41381\ : std_logic;
signal \N__41378\ : std_logic;
signal \N__41377\ : std_logic;
signal \N__41376\ : std_logic;
signal \N__41373\ : std_logic;
signal \N__41370\ : std_logic;
signal \N__41369\ : std_logic;
signal \N__41366\ : std_logic;
signal \N__41361\ : std_logic;
signal \N__41358\ : std_logic;
signal \N__41355\ : std_logic;
signal \N__41350\ : std_logic;
signal \N__41345\ : std_logic;
signal \N__41344\ : std_logic;
signal \N__41341\ : std_logic;
signal \N__41338\ : std_logic;
signal \N__41337\ : std_logic;
signal \N__41334\ : std_logic;
signal \N__41331\ : std_logic;
signal \N__41328\ : std_logic;
signal \N__41321\ : std_logic;
signal \N__41318\ : std_logic;
signal \N__41315\ : std_logic;
signal \N__41312\ : std_logic;
signal \N__41309\ : std_logic;
signal \N__41306\ : std_logic;
signal \N__41303\ : std_logic;
signal \N__41302\ : std_logic;
signal \N__41301\ : std_logic;
signal \N__41298\ : std_logic;
signal \N__41295\ : std_logic;
signal \N__41292\ : std_logic;
signal \N__41289\ : std_logic;
signal \N__41286\ : std_logic;
signal \N__41283\ : std_logic;
signal \N__41280\ : std_logic;
signal \N__41275\ : std_logic;
signal \N__41274\ : std_logic;
signal \N__41269\ : std_logic;
signal \N__41266\ : std_logic;
signal \N__41263\ : std_logic;
signal \N__41258\ : std_logic;
signal \N__41255\ : std_logic;
signal \N__41252\ : std_logic;
signal \N__41251\ : std_logic;
signal \N__41250\ : std_logic;
signal \N__41247\ : std_logic;
signal \N__41244\ : std_logic;
signal \N__41241\ : std_logic;
signal \N__41238\ : std_logic;
signal \N__41235\ : std_logic;
signal \N__41232\ : std_logic;
signal \N__41231\ : std_logic;
signal \N__41228\ : std_logic;
signal \N__41225\ : std_logic;
signal \N__41222\ : std_logic;
signal \N__41219\ : std_logic;
signal \N__41210\ : std_logic;
signal \N__41209\ : std_logic;
signal \N__41206\ : std_logic;
signal \N__41203\ : std_logic;
signal \N__41200\ : std_logic;
signal \N__41199\ : std_logic;
signal \N__41196\ : std_logic;
signal \N__41193\ : std_logic;
signal \N__41190\ : std_logic;
signal \N__41183\ : std_logic;
signal \N__41180\ : std_logic;
signal \N__41179\ : std_logic;
signal \N__41176\ : std_logic;
signal \N__41173\ : std_logic;
signal \N__41170\ : std_logic;
signal \N__41167\ : std_logic;
signal \N__41164\ : std_logic;
signal \N__41159\ : std_logic;
signal \N__41156\ : std_logic;
signal \N__41153\ : std_logic;
signal \N__41150\ : std_logic;
signal \N__41147\ : std_logic;
signal \N__41144\ : std_logic;
signal \N__41141\ : std_logic;
signal \N__41138\ : std_logic;
signal \N__41135\ : std_logic;
signal \N__41134\ : std_logic;
signal \N__41133\ : std_logic;
signal \N__41132\ : std_logic;
signal \N__41129\ : std_logic;
signal \N__41126\ : std_logic;
signal \N__41121\ : std_logic;
signal \N__41116\ : std_logic;
signal \N__41113\ : std_logic;
signal \N__41108\ : std_logic;
signal \N__41105\ : std_logic;
signal \N__41104\ : std_logic;
signal \N__41103\ : std_logic;
signal \N__41100\ : std_logic;
signal \N__41097\ : std_logic;
signal \N__41094\ : std_logic;
signal \N__41087\ : std_logic;
signal \N__41084\ : std_logic;
signal \N__41081\ : std_logic;
signal \N__41080\ : std_logic;
signal \N__41079\ : std_logic;
signal \N__41076\ : std_logic;
signal \N__41073\ : std_logic;
signal \N__41070\ : std_logic;
signal \N__41065\ : std_logic;
signal \N__41060\ : std_logic;
signal \N__41059\ : std_logic;
signal \N__41056\ : std_logic;
signal \N__41055\ : std_logic;
signal \N__41052\ : std_logic;
signal \N__41049\ : std_logic;
signal \N__41048\ : std_logic;
signal \N__41045\ : std_logic;
signal \N__41042\ : std_logic;
signal \N__41039\ : std_logic;
signal \N__41036\ : std_logic;
signal \N__41033\ : std_logic;
signal \N__41030\ : std_logic;
signal \N__41025\ : std_logic;
signal \N__41018\ : std_logic;
signal \N__41017\ : std_logic;
signal \N__41014\ : std_logic;
signal \N__41011\ : std_logic;
signal \N__41008\ : std_logic;
signal \N__41005\ : std_logic;
signal \N__41002\ : std_logic;
signal \N__40999\ : std_logic;
signal \N__40998\ : std_logic;
signal \N__40993\ : std_logic;
signal \N__40990\ : std_logic;
signal \N__40985\ : std_logic;
signal \N__40984\ : std_logic;
signal \N__40983\ : std_logic;
signal \N__40980\ : std_logic;
signal \N__40977\ : std_logic;
signal \N__40974\ : std_logic;
signal \N__40971\ : std_logic;
signal \N__40968\ : std_logic;
signal \N__40965\ : std_logic;
signal \N__40964\ : std_logic;
signal \N__40957\ : std_logic;
signal \N__40954\ : std_logic;
signal \N__40949\ : std_logic;
signal \N__40948\ : std_logic;
signal \N__40945\ : std_logic;
signal \N__40942\ : std_logic;
signal \N__40939\ : std_logic;
signal \N__40936\ : std_logic;
signal \N__40933\ : std_logic;
signal \N__40932\ : std_logic;
signal \N__40929\ : std_logic;
signal \N__40926\ : std_logic;
signal \N__40923\ : std_logic;
signal \N__40916\ : std_logic;
signal \N__40913\ : std_logic;
signal \N__40910\ : std_logic;
signal \N__40909\ : std_logic;
signal \N__40906\ : std_logic;
signal \N__40903\ : std_logic;
signal \N__40900\ : std_logic;
signal \N__40899\ : std_logic;
signal \N__40896\ : std_logic;
signal \N__40893\ : std_logic;
signal \N__40890\ : std_logic;
signal \N__40887\ : std_logic;
signal \N__40886\ : std_logic;
signal \N__40883\ : std_logic;
signal \N__40880\ : std_logic;
signal \N__40877\ : std_logic;
signal \N__40874\ : std_logic;
signal \N__40869\ : std_logic;
signal \N__40862\ : std_logic;
signal \N__40859\ : std_logic;
signal \N__40856\ : std_logic;
signal \N__40853\ : std_logic;
signal \N__40850\ : std_logic;
signal \N__40847\ : std_logic;
signal \N__40844\ : std_logic;
signal \N__40841\ : std_logic;
signal \N__40838\ : std_logic;
signal \N__40837\ : std_logic;
signal \N__40836\ : std_logic;
signal \N__40835\ : std_logic;
signal \N__40832\ : std_logic;
signal \N__40829\ : std_logic;
signal \N__40824\ : std_logic;
signal \N__40817\ : std_logic;
signal \N__40814\ : std_logic;
signal \N__40811\ : std_logic;
signal \N__40810\ : std_logic;
signal \N__40809\ : std_logic;
signal \N__40806\ : std_logic;
signal \N__40803\ : std_logic;
signal \N__40800\ : std_logic;
signal \N__40793\ : std_logic;
signal \N__40790\ : std_logic;
signal \N__40787\ : std_logic;
signal \N__40784\ : std_logic;
signal \N__40781\ : std_logic;
signal \N__40778\ : std_logic;
signal \N__40775\ : std_logic;
signal \N__40772\ : std_logic;
signal \N__40769\ : std_logic;
signal \N__40766\ : std_logic;
signal \N__40763\ : std_logic;
signal \N__40760\ : std_logic;
signal \N__40757\ : std_logic;
signal \N__40754\ : std_logic;
signal \N__40751\ : std_logic;
signal \N__40750\ : std_logic;
signal \N__40747\ : std_logic;
signal \N__40746\ : std_logic;
signal \N__40739\ : std_logic;
signal \N__40736\ : std_logic;
signal \N__40733\ : std_logic;
signal \N__40730\ : std_logic;
signal \N__40727\ : std_logic;
signal \N__40724\ : std_logic;
signal \N__40721\ : std_logic;
signal \N__40718\ : std_logic;
signal \N__40715\ : std_logic;
signal \N__40712\ : std_logic;
signal \N__40709\ : std_logic;
signal \N__40706\ : std_logic;
signal \N__40703\ : std_logic;
signal \N__40700\ : std_logic;
signal \N__40697\ : std_logic;
signal \N__40694\ : std_logic;
signal \N__40691\ : std_logic;
signal \N__40690\ : std_logic;
signal \N__40687\ : std_logic;
signal \N__40684\ : std_logic;
signal \N__40679\ : std_logic;
signal \N__40678\ : std_logic;
signal \N__40675\ : std_logic;
signal \N__40672\ : std_logic;
signal \N__40671\ : std_logic;
signal \N__40670\ : std_logic;
signal \N__40667\ : std_logic;
signal \N__40664\ : std_logic;
signal \N__40659\ : std_logic;
signal \N__40656\ : std_logic;
signal \N__40651\ : std_logic;
signal \N__40648\ : std_logic;
signal \N__40643\ : std_logic;
signal \N__40640\ : std_logic;
signal \N__40639\ : std_logic;
signal \N__40636\ : std_logic;
signal \N__40631\ : std_logic;
signal \N__40628\ : std_logic;
signal \N__40627\ : std_logic;
signal \N__40626\ : std_logic;
signal \N__40623\ : std_logic;
signal \N__40622\ : std_logic;
signal \N__40619\ : std_logic;
signal \N__40616\ : std_logic;
signal \N__40613\ : std_logic;
signal \N__40610\ : std_logic;
signal \N__40607\ : std_logic;
signal \N__40604\ : std_logic;
signal \N__40601\ : std_logic;
signal \N__40598\ : std_logic;
signal \N__40595\ : std_logic;
signal \N__40586\ : std_logic;
signal \N__40583\ : std_logic;
signal \N__40582\ : std_logic;
signal \N__40579\ : std_logic;
signal \N__40578\ : std_logic;
signal \N__40575\ : std_logic;
signal \N__40572\ : std_logic;
signal \N__40569\ : std_logic;
signal \N__40566\ : std_logic;
signal \N__40563\ : std_logic;
signal \N__40556\ : std_logic;
signal \N__40555\ : std_logic;
signal \N__40550\ : std_logic;
signal \N__40547\ : std_logic;
signal \N__40544\ : std_logic;
signal \N__40541\ : std_logic;
signal \N__40538\ : std_logic;
signal \N__40535\ : std_logic;
signal \N__40532\ : std_logic;
signal \N__40529\ : std_logic;
signal \N__40526\ : std_logic;
signal \N__40523\ : std_logic;
signal \N__40520\ : std_logic;
signal \N__40517\ : std_logic;
signal \N__40514\ : std_logic;
signal \N__40511\ : std_logic;
signal \N__40508\ : std_logic;
signal \N__40505\ : std_logic;
signal \N__40502\ : std_logic;
signal \N__40499\ : std_logic;
signal \N__40496\ : std_logic;
signal \N__40493\ : std_logic;
signal \N__40490\ : std_logic;
signal \N__40487\ : std_logic;
signal \N__40484\ : std_logic;
signal \N__40481\ : std_logic;
signal \N__40478\ : std_logic;
signal \N__40475\ : std_logic;
signal \N__40472\ : std_logic;
signal \N__40469\ : std_logic;
signal \N__40466\ : std_logic;
signal \N__40463\ : std_logic;
signal \N__40460\ : std_logic;
signal \N__40457\ : std_logic;
signal \N__40454\ : std_logic;
signal \N__40451\ : std_logic;
signal \N__40448\ : std_logic;
signal \N__40445\ : std_logic;
signal \N__40442\ : std_logic;
signal \N__40439\ : std_logic;
signal \N__40436\ : std_logic;
signal \N__40433\ : std_logic;
signal \N__40430\ : std_logic;
signal \N__40427\ : std_logic;
signal \N__40424\ : std_logic;
signal \N__40421\ : std_logic;
signal \N__40418\ : std_logic;
signal \N__40415\ : std_logic;
signal \N__40412\ : std_logic;
signal \N__40409\ : std_logic;
signal \N__40406\ : std_logic;
signal \N__40403\ : std_logic;
signal \N__40400\ : std_logic;
signal \N__40397\ : std_logic;
signal \N__40394\ : std_logic;
signal \N__40391\ : std_logic;
signal \N__40388\ : std_logic;
signal \N__40385\ : std_logic;
signal \N__40382\ : std_logic;
signal \N__40379\ : std_logic;
signal \N__40376\ : std_logic;
signal \N__40373\ : std_logic;
signal \N__40370\ : std_logic;
signal \N__40367\ : std_logic;
signal \N__40364\ : std_logic;
signal \N__40361\ : std_logic;
signal \N__40358\ : std_logic;
signal \N__40357\ : std_logic;
signal \N__40352\ : std_logic;
signal \N__40349\ : std_logic;
signal \N__40346\ : std_logic;
signal \N__40343\ : std_logic;
signal \N__40342\ : std_logic;
signal \N__40337\ : std_logic;
signal \N__40334\ : std_logic;
signal \N__40331\ : std_logic;
signal \N__40328\ : std_logic;
signal \N__40325\ : std_logic;
signal \N__40324\ : std_logic;
signal \N__40323\ : std_logic;
signal \N__40322\ : std_logic;
signal \N__40319\ : std_logic;
signal \N__40316\ : std_logic;
signal \N__40313\ : std_logic;
signal \N__40310\ : std_logic;
signal \N__40301\ : std_logic;
signal \N__40298\ : std_logic;
signal \N__40297\ : std_logic;
signal \N__40294\ : std_logic;
signal \N__40293\ : std_logic;
signal \N__40290\ : std_logic;
signal \N__40287\ : std_logic;
signal \N__40284\ : std_logic;
signal \N__40277\ : std_logic;
signal \N__40276\ : std_logic;
signal \N__40275\ : std_logic;
signal \N__40272\ : std_logic;
signal \N__40269\ : std_logic;
signal \N__40266\ : std_logic;
signal \N__40265\ : std_logic;
signal \N__40262\ : std_logic;
signal \N__40259\ : std_logic;
signal \N__40256\ : std_logic;
signal \N__40253\ : std_logic;
signal \N__40250\ : std_logic;
signal \N__40247\ : std_logic;
signal \N__40244\ : std_logic;
signal \N__40241\ : std_logic;
signal \N__40232\ : std_logic;
signal \N__40229\ : std_logic;
signal \N__40226\ : std_logic;
signal \N__40223\ : std_logic;
signal \N__40220\ : std_logic;
signal \N__40217\ : std_logic;
signal \N__40214\ : std_logic;
signal \N__40211\ : std_logic;
signal \N__40208\ : std_logic;
signal \N__40205\ : std_logic;
signal \N__40202\ : std_logic;
signal \N__40199\ : std_logic;
signal \N__40196\ : std_logic;
signal \N__40193\ : std_logic;
signal \N__40190\ : std_logic;
signal \N__40187\ : std_logic;
signal \N__40184\ : std_logic;
signal \N__40181\ : std_logic;
signal \N__40178\ : std_logic;
signal \N__40175\ : std_logic;
signal \N__40172\ : std_logic;
signal \N__40169\ : std_logic;
signal \N__40166\ : std_logic;
signal \N__40163\ : std_logic;
signal \N__40160\ : std_logic;
signal \N__40157\ : std_logic;
signal \N__40154\ : std_logic;
signal \N__40151\ : std_logic;
signal \N__40148\ : std_logic;
signal \N__40145\ : std_logic;
signal \N__40142\ : std_logic;
signal \N__40139\ : std_logic;
signal \N__40136\ : std_logic;
signal \N__40133\ : std_logic;
signal \N__40130\ : std_logic;
signal \N__40127\ : std_logic;
signal \N__40124\ : std_logic;
signal \N__40121\ : std_logic;
signal \N__40120\ : std_logic;
signal \N__40119\ : std_logic;
signal \N__40118\ : std_logic;
signal \N__40115\ : std_logic;
signal \N__40112\ : std_logic;
signal \N__40109\ : std_logic;
signal \N__40106\ : std_logic;
signal \N__40097\ : std_logic;
signal \N__40094\ : std_logic;
signal \N__40093\ : std_logic;
signal \N__40090\ : std_logic;
signal \N__40089\ : std_logic;
signal \N__40086\ : std_logic;
signal \N__40083\ : std_logic;
signal \N__40080\ : std_logic;
signal \N__40073\ : std_logic;
signal \N__40072\ : std_logic;
signal \N__40069\ : std_logic;
signal \N__40066\ : std_logic;
signal \N__40065\ : std_logic;
signal \N__40064\ : std_logic;
signal \N__40061\ : std_logic;
signal \N__40058\ : std_logic;
signal \N__40055\ : std_logic;
signal \N__40052\ : std_logic;
signal \N__40043\ : std_logic;
signal \N__40040\ : std_logic;
signal \N__40039\ : std_logic;
signal \N__40036\ : std_logic;
signal \N__40035\ : std_logic;
signal \N__40032\ : std_logic;
signal \N__40029\ : std_logic;
signal \N__40026\ : std_logic;
signal \N__40019\ : std_logic;
signal \N__40016\ : std_logic;
signal \N__40013\ : std_logic;
signal \N__40010\ : std_logic;
signal \N__40009\ : std_logic;
signal \N__40008\ : std_logic;
signal \N__40003\ : std_logic;
signal \N__40002\ : std_logic;
signal \N__39999\ : std_logic;
signal \N__39996\ : std_logic;
signal \N__39993\ : std_logic;
signal \N__39990\ : std_logic;
signal \N__39985\ : std_logic;
signal \N__39980\ : std_logic;
signal \N__39979\ : std_logic;
signal \N__39978\ : std_logic;
signal \N__39975\ : std_logic;
signal \N__39972\ : std_logic;
signal \N__39967\ : std_logic;
signal \N__39964\ : std_logic;
signal \N__39961\ : std_logic;
signal \N__39958\ : std_logic;
signal \N__39953\ : std_logic;
signal \N__39950\ : std_logic;
signal \N__39949\ : std_logic;
signal \N__39946\ : std_logic;
signal \N__39943\ : std_logic;
signal \N__39940\ : std_logic;
signal \N__39939\ : std_logic;
signal \N__39938\ : std_logic;
signal \N__39935\ : std_logic;
signal \N__39932\ : std_logic;
signal \N__39929\ : std_logic;
signal \N__39926\ : std_logic;
signal \N__39923\ : std_logic;
signal \N__39920\ : std_logic;
signal \N__39915\ : std_logic;
signal \N__39908\ : std_logic;
signal \N__39905\ : std_logic;
signal \N__39904\ : std_logic;
signal \N__39903\ : std_logic;
signal \N__39900\ : std_logic;
signal \N__39897\ : std_logic;
signal \N__39894\ : std_logic;
signal \N__39891\ : std_logic;
signal \N__39886\ : std_logic;
signal \N__39881\ : std_logic;
signal \N__39878\ : std_logic;
signal \N__39875\ : std_logic;
signal \N__39872\ : std_logic;
signal \N__39869\ : std_logic;
signal \N__39866\ : std_logic;
signal \N__39863\ : std_logic;
signal \N__39860\ : std_logic;
signal \N__39857\ : std_logic;
signal \N__39856\ : std_logic;
signal \N__39853\ : std_logic;
signal \N__39850\ : std_logic;
signal \N__39847\ : std_logic;
signal \N__39846\ : std_logic;
signal \N__39845\ : std_logic;
signal \N__39840\ : std_logic;
signal \N__39839\ : std_logic;
signal \N__39836\ : std_logic;
signal \N__39833\ : std_logic;
signal \N__39830\ : std_logic;
signal \N__39827\ : std_logic;
signal \N__39818\ : std_logic;
signal \N__39815\ : std_logic;
signal \N__39812\ : std_logic;
signal \N__39811\ : std_logic;
signal \N__39808\ : std_logic;
signal \N__39805\ : std_logic;
signal \N__39800\ : std_logic;
signal \N__39799\ : std_logic;
signal \N__39796\ : std_logic;
signal \N__39793\ : std_logic;
signal \N__39792\ : std_logic;
signal \N__39789\ : std_logic;
signal \N__39786\ : std_logic;
signal \N__39783\ : std_logic;
signal \N__39780\ : std_logic;
signal \N__39777\ : std_logic;
signal \N__39770\ : std_logic;
signal \N__39769\ : std_logic;
signal \N__39768\ : std_logic;
signal \N__39767\ : std_logic;
signal \N__39764\ : std_logic;
signal \N__39761\ : std_logic;
signal \N__39758\ : std_logic;
signal \N__39755\ : std_logic;
signal \N__39752\ : std_logic;
signal \N__39747\ : std_logic;
signal \N__39744\ : std_logic;
signal \N__39739\ : std_logic;
signal \N__39736\ : std_logic;
signal \N__39731\ : std_logic;
signal \N__39728\ : std_logic;
signal \N__39725\ : std_logic;
signal \N__39722\ : std_logic;
signal \N__39719\ : std_logic;
signal \N__39716\ : std_logic;
signal \N__39713\ : std_logic;
signal \N__39710\ : std_logic;
signal \N__39707\ : std_logic;
signal \N__39704\ : std_logic;
signal \N__39701\ : std_logic;
signal \N__39700\ : std_logic;
signal \N__39699\ : std_logic;
signal \N__39696\ : std_logic;
signal \N__39691\ : std_logic;
signal \N__39690\ : std_logic;
signal \N__39687\ : std_logic;
signal \N__39684\ : std_logic;
signal \N__39681\ : std_logic;
signal \N__39674\ : std_logic;
signal \N__39671\ : std_logic;
signal \N__39668\ : std_logic;
signal \N__39665\ : std_logic;
signal \N__39662\ : std_logic;
signal \N__39659\ : std_logic;
signal \N__39656\ : std_logic;
signal \N__39655\ : std_logic;
signal \N__39652\ : std_logic;
signal \N__39649\ : std_logic;
signal \N__39646\ : std_logic;
signal \N__39643\ : std_logic;
signal \N__39642\ : std_logic;
signal \N__39641\ : std_logic;
signal \N__39636\ : std_logic;
signal \N__39633\ : std_logic;
signal \N__39630\ : std_logic;
signal \N__39623\ : std_logic;
signal \N__39620\ : std_logic;
signal \N__39619\ : std_logic;
signal \N__39618\ : std_logic;
signal \N__39615\ : std_logic;
signal \N__39612\ : std_logic;
signal \N__39609\ : std_logic;
signal \N__39606\ : std_logic;
signal \N__39599\ : std_logic;
signal \N__39598\ : std_logic;
signal \N__39597\ : std_logic;
signal \N__39594\ : std_logic;
signal \N__39591\ : std_logic;
signal \N__39588\ : std_logic;
signal \N__39585\ : std_logic;
signal \N__39582\ : std_logic;
signal \N__39579\ : std_logic;
signal \N__39576\ : std_logic;
signal \N__39573\ : std_logic;
signal \N__39566\ : std_logic;
signal \N__39563\ : std_logic;
signal \N__39560\ : std_logic;
signal \N__39557\ : std_logic;
signal \N__39554\ : std_logic;
signal \N__39551\ : std_logic;
signal \N__39548\ : std_logic;
signal \N__39545\ : std_logic;
signal \N__39542\ : std_logic;
signal \N__39539\ : std_logic;
signal \N__39536\ : std_logic;
signal \N__39533\ : std_logic;
signal \N__39530\ : std_logic;
signal \N__39527\ : std_logic;
signal \N__39524\ : std_logic;
signal \N__39521\ : std_logic;
signal \N__39518\ : std_logic;
signal \N__39515\ : std_logic;
signal \N__39512\ : std_logic;
signal \N__39509\ : std_logic;
signal \N__39506\ : std_logic;
signal \N__39503\ : std_logic;
signal \N__39500\ : std_logic;
signal \N__39497\ : std_logic;
signal \N__39494\ : std_logic;
signal \N__39491\ : std_logic;
signal \N__39488\ : std_logic;
signal \N__39485\ : std_logic;
signal \N__39482\ : std_logic;
signal \N__39479\ : std_logic;
signal \N__39476\ : std_logic;
signal \N__39473\ : std_logic;
signal \N__39470\ : std_logic;
signal \N__39467\ : std_logic;
signal \N__39464\ : std_logic;
signal \N__39461\ : std_logic;
signal \N__39458\ : std_logic;
signal \N__39455\ : std_logic;
signal \N__39452\ : std_logic;
signal \N__39449\ : std_logic;
signal \N__39446\ : std_logic;
signal \N__39443\ : std_logic;
signal \N__39442\ : std_logic;
signal \N__39439\ : std_logic;
signal \N__39436\ : std_logic;
signal \N__39435\ : std_logic;
signal \N__39432\ : std_logic;
signal \N__39427\ : std_logic;
signal \N__39422\ : std_logic;
signal \N__39419\ : std_logic;
signal \N__39416\ : std_logic;
signal \N__39413\ : std_logic;
signal \N__39410\ : std_logic;
signal \N__39407\ : std_logic;
signal \N__39404\ : std_logic;
signal \N__39401\ : std_logic;
signal \N__39398\ : std_logic;
signal \N__39395\ : std_logic;
signal \N__39392\ : std_logic;
signal \N__39389\ : std_logic;
signal \N__39386\ : std_logic;
signal \N__39383\ : std_logic;
signal \N__39380\ : std_logic;
signal \N__39377\ : std_logic;
signal \N__39374\ : std_logic;
signal \N__39371\ : std_logic;
signal \N__39368\ : std_logic;
signal \N__39365\ : std_logic;
signal \N__39362\ : std_logic;
signal \N__39359\ : std_logic;
signal \N__39356\ : std_logic;
signal \N__39353\ : std_logic;
signal \N__39350\ : std_logic;
signal \N__39347\ : std_logic;
signal \N__39344\ : std_logic;
signal \N__39341\ : std_logic;
signal \N__39338\ : std_logic;
signal \N__39335\ : std_logic;
signal \N__39332\ : std_logic;
signal \N__39329\ : std_logic;
signal \N__39326\ : std_logic;
signal \N__39323\ : std_logic;
signal \N__39320\ : std_logic;
signal \N__39317\ : std_logic;
signal \N__39314\ : std_logic;
signal \N__39311\ : std_logic;
signal \N__39308\ : std_logic;
signal \N__39305\ : std_logic;
signal \N__39302\ : std_logic;
signal \N__39299\ : std_logic;
signal \N__39296\ : std_logic;
signal \N__39293\ : std_logic;
signal \N__39290\ : std_logic;
signal \N__39287\ : std_logic;
signal \N__39284\ : std_logic;
signal \N__39281\ : std_logic;
signal \N__39278\ : std_logic;
signal \N__39275\ : std_logic;
signal \N__39272\ : std_logic;
signal \N__39269\ : std_logic;
signal \N__39266\ : std_logic;
signal \N__39263\ : std_logic;
signal \N__39260\ : std_logic;
signal \N__39257\ : std_logic;
signal \N__39254\ : std_logic;
signal \N__39251\ : std_logic;
signal \N__39248\ : std_logic;
signal \N__39245\ : std_logic;
signal \N__39242\ : std_logic;
signal \N__39239\ : std_logic;
signal \N__39236\ : std_logic;
signal \N__39233\ : std_logic;
signal \N__39230\ : std_logic;
signal \N__39227\ : std_logic;
signal \N__39224\ : std_logic;
signal \N__39221\ : std_logic;
signal \N__39218\ : std_logic;
signal \N__39217\ : std_logic;
signal \N__39214\ : std_logic;
signal \N__39211\ : std_logic;
signal \N__39208\ : std_logic;
signal \N__39203\ : std_logic;
signal \N__39200\ : std_logic;
signal \N__39199\ : std_logic;
signal \N__39198\ : std_logic;
signal \N__39195\ : std_logic;
signal \N__39192\ : std_logic;
signal \N__39189\ : std_logic;
signal \N__39184\ : std_logic;
signal \N__39179\ : std_logic;
signal \N__39176\ : std_logic;
signal \N__39175\ : std_logic;
signal \N__39174\ : std_logic;
signal \N__39173\ : std_logic;
signal \N__39170\ : std_logic;
signal \N__39167\ : std_logic;
signal \N__39162\ : std_logic;
signal \N__39159\ : std_logic;
signal \N__39156\ : std_logic;
signal \N__39153\ : std_logic;
signal \N__39150\ : std_logic;
signal \N__39147\ : std_logic;
signal \N__39144\ : std_logic;
signal \N__39137\ : std_logic;
signal \N__39134\ : std_logic;
signal \N__39131\ : std_logic;
signal \N__39128\ : std_logic;
signal \N__39125\ : std_logic;
signal \N__39124\ : std_logic;
signal \N__39121\ : std_logic;
signal \N__39116\ : std_logic;
signal \N__39115\ : std_logic;
signal \N__39112\ : std_logic;
signal \N__39109\ : std_logic;
signal \N__39106\ : std_logic;
signal \N__39101\ : std_logic;
signal \N__39100\ : std_logic;
signal \N__39099\ : std_logic;
signal \N__39096\ : std_logic;
signal \N__39093\ : std_logic;
signal \N__39088\ : std_logic;
signal \N__39083\ : std_logic;
signal \N__39080\ : std_logic;
signal \N__39077\ : std_logic;
signal \N__39074\ : std_logic;
signal \N__39071\ : std_logic;
signal \N__39070\ : std_logic;
signal \N__39065\ : std_logic;
signal \N__39062\ : std_logic;
signal \N__39059\ : std_logic;
signal \N__39056\ : std_logic;
signal \N__39053\ : std_logic;
signal \N__39050\ : std_logic;
signal \N__39049\ : std_logic;
signal \N__39048\ : std_logic;
signal \N__39043\ : std_logic;
signal \N__39040\ : std_logic;
signal \N__39037\ : std_logic;
signal \N__39032\ : std_logic;
signal \N__39029\ : std_logic;
signal \N__39026\ : std_logic;
signal \N__39025\ : std_logic;
signal \N__39024\ : std_logic;
signal \N__39021\ : std_logic;
signal \N__39018\ : std_logic;
signal \N__39015\ : std_logic;
signal \N__39010\ : std_logic;
signal \N__39005\ : std_logic;
signal \N__39002\ : std_logic;
signal \N__39001\ : std_logic;
signal \N__38998\ : std_logic;
signal \N__38995\ : std_logic;
signal \N__38992\ : std_logic;
signal \N__38991\ : std_logic;
signal \N__38988\ : std_logic;
signal \N__38985\ : std_logic;
signal \N__38982\ : std_logic;
signal \N__38977\ : std_logic;
signal \N__38972\ : std_logic;
signal \N__38969\ : std_logic;
signal \N__38968\ : std_logic;
signal \N__38963\ : std_logic;
signal \N__38962\ : std_logic;
signal \N__38959\ : std_logic;
signal \N__38956\ : std_logic;
signal \N__38953\ : std_logic;
signal \N__38948\ : std_logic;
signal \N__38945\ : std_logic;
signal \N__38944\ : std_logic;
signal \N__38941\ : std_logic;
signal \N__38938\ : std_logic;
signal \N__38933\ : std_logic;
signal \N__38932\ : std_logic;
signal \N__38929\ : std_logic;
signal \N__38926\ : std_logic;
signal \N__38923\ : std_logic;
signal \N__38918\ : std_logic;
signal \N__38915\ : std_logic;
signal \N__38914\ : std_logic;
signal \N__38911\ : std_logic;
signal \N__38908\ : std_logic;
signal \N__38905\ : std_logic;
signal \N__38902\ : std_logic;
signal \N__38901\ : std_logic;
signal \N__38896\ : std_logic;
signal \N__38893\ : std_logic;
signal \N__38890\ : std_logic;
signal \N__38885\ : std_logic;
signal \N__38882\ : std_logic;
signal \N__38879\ : std_logic;
signal \N__38878\ : std_logic;
signal \N__38877\ : std_logic;
signal \N__38874\ : std_logic;
signal \N__38871\ : std_logic;
signal \N__38868\ : std_logic;
signal \N__38863\ : std_logic;
signal \N__38858\ : std_logic;
signal \N__38855\ : std_logic;
signal \N__38854\ : std_logic;
signal \N__38853\ : std_logic;
signal \N__38848\ : std_logic;
signal \N__38845\ : std_logic;
signal \N__38842\ : std_logic;
signal \N__38837\ : std_logic;
signal \N__38834\ : std_logic;
signal \N__38833\ : std_logic;
signal \N__38830\ : std_logic;
signal \N__38827\ : std_logic;
signal \N__38824\ : std_logic;
signal \N__38819\ : std_logic;
signal \N__38816\ : std_logic;
signal \N__38815\ : std_logic;
signal \N__38814\ : std_logic;
signal \N__38811\ : std_logic;
signal \N__38808\ : std_logic;
signal \N__38805\ : std_logic;
signal \N__38802\ : std_logic;
signal \N__38797\ : std_logic;
signal \N__38796\ : std_logic;
signal \N__38791\ : std_logic;
signal \N__38788\ : std_logic;
signal \N__38783\ : std_logic;
signal \N__38780\ : std_logic;
signal \N__38779\ : std_logic;
signal \N__38774\ : std_logic;
signal \N__38773\ : std_logic;
signal \N__38770\ : std_logic;
signal \N__38767\ : std_logic;
signal \N__38764\ : std_logic;
signal \N__38759\ : std_logic;
signal \N__38756\ : std_logic;
signal \N__38755\ : std_logic;
signal \N__38752\ : std_logic;
signal \N__38749\ : std_logic;
signal \N__38748\ : std_logic;
signal \N__38743\ : std_logic;
signal \N__38740\ : std_logic;
signal \N__38737\ : std_logic;
signal \N__38732\ : std_logic;
signal \N__38729\ : std_logic;
signal \N__38728\ : std_logic;
signal \N__38725\ : std_logic;
signal \N__38722\ : std_logic;
signal \N__38721\ : std_logic;
signal \N__38716\ : std_logic;
signal \N__38713\ : std_logic;
signal \N__38710\ : std_logic;
signal \N__38705\ : std_logic;
signal \N__38702\ : std_logic;
signal \N__38701\ : std_logic;
signal \N__38696\ : std_logic;
signal \N__38695\ : std_logic;
signal \N__38692\ : std_logic;
signal \N__38689\ : std_logic;
signal \N__38686\ : std_logic;
signal \N__38681\ : std_logic;
signal \N__38678\ : std_logic;
signal \N__38675\ : std_logic;
signal \N__38674\ : std_logic;
signal \N__38673\ : std_logic;
signal \N__38670\ : std_logic;
signal \N__38667\ : std_logic;
signal \N__38664\ : std_logic;
signal \N__38659\ : std_logic;
signal \N__38654\ : std_logic;
signal \N__38651\ : std_logic;
signal \N__38650\ : std_logic;
signal \N__38647\ : std_logic;
signal \N__38644\ : std_logic;
signal \N__38641\ : std_logic;
signal \N__38640\ : std_logic;
signal \N__38635\ : std_logic;
signal \N__38632\ : std_logic;
signal \N__38629\ : std_logic;
signal \N__38624\ : std_logic;
signal \N__38621\ : std_logic;
signal \N__38618\ : std_logic;
signal \N__38617\ : std_logic;
signal \N__38616\ : std_logic;
signal \N__38613\ : std_logic;
signal \N__38610\ : std_logic;
signal \N__38607\ : std_logic;
signal \N__38602\ : std_logic;
signal \N__38597\ : std_logic;
signal \N__38594\ : std_logic;
signal \N__38593\ : std_logic;
signal \N__38590\ : std_logic;
signal \N__38587\ : std_logic;
signal \N__38586\ : std_logic;
signal \N__38581\ : std_logic;
signal \N__38578\ : std_logic;
signal \N__38575\ : std_logic;
signal \N__38570\ : std_logic;
signal \N__38567\ : std_logic;
signal \N__38566\ : std_logic;
signal \N__38563\ : std_logic;
signal \N__38560\ : std_logic;
signal \N__38559\ : std_logic;
signal \N__38556\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38550\ : std_logic;
signal \N__38545\ : std_logic;
signal \N__38540\ : std_logic;
signal \N__38537\ : std_logic;
signal \N__38536\ : std_logic;
signal \N__38531\ : std_logic;
signal \N__38530\ : std_logic;
signal \N__38527\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38521\ : std_logic;
signal \N__38516\ : std_logic;
signal \N__38513\ : std_logic;
signal \N__38512\ : std_logic;
signal \N__38509\ : std_logic;
signal \N__38506\ : std_logic;
signal \N__38505\ : std_logic;
signal \N__38504\ : std_logic;
signal \N__38501\ : std_logic;
signal \N__38498\ : std_logic;
signal \N__38495\ : std_logic;
signal \N__38492\ : std_logic;
signal \N__38483\ : std_logic;
signal \N__38480\ : std_logic;
signal \N__38479\ : std_logic;
signal \N__38476\ : std_logic;
signal \N__38473\ : std_logic;
signal \N__38472\ : std_logic;
signal \N__38467\ : std_logic;
signal \N__38464\ : std_logic;
signal \N__38461\ : std_logic;
signal \N__38456\ : std_logic;
signal \N__38453\ : std_logic;
signal \N__38452\ : std_logic;
signal \N__38449\ : std_logic;
signal \N__38446\ : std_logic;
signal \N__38445\ : std_logic;
signal \N__38440\ : std_logic;
signal \N__38437\ : std_logic;
signal \N__38434\ : std_logic;
signal \N__38429\ : std_logic;
signal \N__38426\ : std_logic;
signal \N__38425\ : std_logic;
signal \N__38420\ : std_logic;
signal \N__38419\ : std_logic;
signal \N__38416\ : std_logic;
signal \N__38413\ : std_logic;
signal \N__38410\ : std_logic;
signal \N__38405\ : std_logic;
signal \N__38404\ : std_logic;
signal \N__38401\ : std_logic;
signal \N__38400\ : std_logic;
signal \N__38399\ : std_logic;
signal \N__38396\ : std_logic;
signal \N__38393\ : std_logic;
signal \N__38390\ : std_logic;
signal \N__38387\ : std_logic;
signal \N__38384\ : std_logic;
signal \N__38381\ : std_logic;
signal \N__38378\ : std_logic;
signal \N__38369\ : std_logic;
signal \N__38366\ : std_logic;
signal \N__38365\ : std_logic;
signal \N__38360\ : std_logic;
signal \N__38359\ : std_logic;
signal \N__38356\ : std_logic;
signal \N__38353\ : std_logic;
signal \N__38350\ : std_logic;
signal \N__38345\ : std_logic;
signal \N__38342\ : std_logic;
signal \N__38339\ : std_logic;
signal \N__38338\ : std_logic;
signal \N__38337\ : std_logic;
signal \N__38336\ : std_logic;
signal \N__38333\ : std_logic;
signal \N__38328\ : std_logic;
signal \N__38325\ : std_logic;
signal \N__38318\ : std_logic;
signal \N__38315\ : std_logic;
signal \N__38314\ : std_logic;
signal \N__38311\ : std_logic;
signal \N__38308\ : std_logic;
signal \N__38305\ : std_logic;
signal \N__38302\ : std_logic;
signal \N__38301\ : std_logic;
signal \N__38296\ : std_logic;
signal \N__38293\ : std_logic;
signal \N__38290\ : std_logic;
signal \N__38285\ : std_logic;
signal \N__38284\ : std_logic;
signal \N__38281\ : std_logic;
signal \N__38278\ : std_logic;
signal \N__38275\ : std_logic;
signal \N__38274\ : std_logic;
signal \N__38273\ : std_logic;
signal \N__38270\ : std_logic;
signal \N__38267\ : std_logic;
signal \N__38262\ : std_logic;
signal \N__38255\ : std_logic;
signal \N__38252\ : std_logic;
signal \N__38251\ : std_logic;
signal \N__38248\ : std_logic;
signal \N__38245\ : std_logic;
signal \N__38242\ : std_logic;
signal \N__38239\ : std_logic;
signal \N__38238\ : std_logic;
signal \N__38233\ : std_logic;
signal \N__38230\ : std_logic;
signal \N__38227\ : std_logic;
signal \N__38222\ : std_logic;
signal \N__38219\ : std_logic;
signal \N__38218\ : std_logic;
signal \N__38213\ : std_logic;
signal \N__38212\ : std_logic;
signal \N__38209\ : std_logic;
signal \N__38206\ : std_logic;
signal \N__38203\ : std_logic;
signal \N__38198\ : std_logic;
signal \N__38195\ : std_logic;
signal \N__38192\ : std_logic;
signal \N__38189\ : std_logic;
signal \N__38186\ : std_logic;
signal \N__38183\ : std_logic;
signal \N__38182\ : std_logic;
signal \N__38181\ : std_logic;
signal \N__38180\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38178\ : std_logic;
signal \N__38177\ : std_logic;
signal \N__38176\ : std_logic;
signal \N__38175\ : std_logic;
signal \N__38174\ : std_logic;
signal \N__38173\ : std_logic;
signal \N__38172\ : std_logic;
signal \N__38171\ : std_logic;
signal \N__38170\ : std_logic;
signal \N__38169\ : std_logic;
signal \N__38168\ : std_logic;
signal \N__38167\ : std_logic;
signal \N__38166\ : std_logic;
signal \N__38165\ : std_logic;
signal \N__38164\ : std_logic;
signal \N__38163\ : std_logic;
signal \N__38162\ : std_logic;
signal \N__38161\ : std_logic;
signal \N__38160\ : std_logic;
signal \N__38159\ : std_logic;
signal \N__38158\ : std_logic;
signal \N__38157\ : std_logic;
signal \N__38156\ : std_logic;
signal \N__38155\ : std_logic;
signal \N__38154\ : std_logic;
signal \N__38149\ : std_logic;
signal \N__38140\ : std_logic;
signal \N__38131\ : std_logic;
signal \N__38122\ : std_logic;
signal \N__38113\ : std_logic;
signal \N__38104\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38086\ : std_logic;
signal \N__38081\ : std_logic;
signal \N__38068\ : std_logic;
signal \N__38063\ : std_logic;
signal \N__38060\ : std_logic;
signal \N__38057\ : std_logic;
signal \N__38056\ : std_logic;
signal \N__38055\ : std_logic;
signal \N__38054\ : std_logic;
signal \N__38051\ : std_logic;
signal \N__38048\ : std_logic;
signal \N__38045\ : std_logic;
signal \N__38042\ : std_logic;
signal \N__38039\ : std_logic;
signal \N__38036\ : std_logic;
signal \N__38033\ : std_logic;
signal \N__38030\ : std_logic;
signal \N__38027\ : std_logic;
signal \N__38024\ : std_logic;
signal \N__38021\ : std_logic;
signal \N__38018\ : std_logic;
signal \N__38009\ : std_logic;
signal \N__38006\ : std_logic;
signal \N__38003\ : std_logic;
signal \N__38000\ : std_logic;
signal \N__37997\ : std_logic;
signal \N__37994\ : std_logic;
signal \N__37991\ : std_logic;
signal \N__37988\ : std_logic;
signal \N__37985\ : std_logic;
signal \N__37982\ : std_logic;
signal \N__37979\ : std_logic;
signal \N__37976\ : std_logic;
signal \N__37973\ : std_logic;
signal \N__37970\ : std_logic;
signal \N__37967\ : std_logic;
signal \N__37964\ : std_logic;
signal \N__37961\ : std_logic;
signal \N__37958\ : std_logic;
signal \N__37955\ : std_logic;
signal \N__37952\ : std_logic;
signal \N__37949\ : std_logic;
signal \N__37948\ : std_logic;
signal \N__37947\ : std_logic;
signal \N__37944\ : std_logic;
signal \N__37943\ : std_logic;
signal \N__37940\ : std_logic;
signal \N__37937\ : std_logic;
signal \N__37934\ : std_logic;
signal \N__37931\ : std_logic;
signal \N__37922\ : std_logic;
signal \N__37919\ : std_logic;
signal \N__37916\ : std_logic;
signal \N__37913\ : std_logic;
signal \N__37910\ : std_logic;
signal \N__37907\ : std_logic;
signal \N__37904\ : std_logic;
signal \N__37901\ : std_logic;
signal \N__37898\ : std_logic;
signal \N__37895\ : std_logic;
signal \N__37892\ : std_logic;
signal \N__37889\ : std_logic;
signal \N__37886\ : std_logic;
signal \N__37883\ : std_logic;
signal \N__37880\ : std_logic;
signal \N__37877\ : std_logic;
signal \N__37874\ : std_logic;
signal \N__37871\ : std_logic;
signal \N__37868\ : std_logic;
signal \N__37865\ : std_logic;
signal \N__37862\ : std_logic;
signal \N__37859\ : std_logic;
signal \N__37856\ : std_logic;
signal \N__37853\ : std_logic;
signal \N__37850\ : std_logic;
signal \N__37847\ : std_logic;
signal \N__37844\ : std_logic;
signal \N__37841\ : std_logic;
signal \N__37838\ : std_logic;
signal \N__37835\ : std_logic;
signal \N__37832\ : std_logic;
signal \N__37829\ : std_logic;
signal \N__37826\ : std_logic;
signal \N__37823\ : std_logic;
signal \N__37820\ : std_logic;
signal \N__37817\ : std_logic;
signal \N__37814\ : std_logic;
signal \N__37811\ : std_logic;
signal \N__37808\ : std_logic;
signal \N__37805\ : std_logic;
signal \N__37802\ : std_logic;
signal \N__37799\ : std_logic;
signal \N__37796\ : std_logic;
signal \N__37793\ : std_logic;
signal \N__37790\ : std_logic;
signal \N__37787\ : std_logic;
signal \N__37784\ : std_logic;
signal \N__37781\ : std_logic;
signal \N__37778\ : std_logic;
signal \N__37775\ : std_logic;
signal \N__37772\ : std_logic;
signal \N__37769\ : std_logic;
signal \N__37766\ : std_logic;
signal \N__37763\ : std_logic;
signal \N__37760\ : std_logic;
signal \N__37757\ : std_logic;
signal \N__37754\ : std_logic;
signal \N__37751\ : std_logic;
signal \N__37748\ : std_logic;
signal \N__37745\ : std_logic;
signal \N__37742\ : std_logic;
signal \N__37739\ : std_logic;
signal \N__37736\ : std_logic;
signal \N__37733\ : std_logic;
signal \N__37730\ : std_logic;
signal \N__37727\ : std_logic;
signal \N__37724\ : std_logic;
signal \N__37721\ : std_logic;
signal \N__37718\ : std_logic;
signal \N__37715\ : std_logic;
signal \N__37712\ : std_logic;
signal \N__37709\ : std_logic;
signal \N__37706\ : std_logic;
signal \N__37703\ : std_logic;
signal \N__37700\ : std_logic;
signal \N__37697\ : std_logic;
signal \N__37694\ : std_logic;
signal \N__37691\ : std_logic;
signal \N__37688\ : std_logic;
signal \N__37685\ : std_logic;
signal \N__37682\ : std_logic;
signal \N__37679\ : std_logic;
signal \N__37676\ : std_logic;
signal \N__37673\ : std_logic;
signal \N__37670\ : std_logic;
signal \N__37667\ : std_logic;
signal \N__37664\ : std_logic;
signal \N__37661\ : std_logic;
signal \N__37658\ : std_logic;
signal \N__37657\ : std_logic;
signal \N__37656\ : std_logic;
signal \N__37653\ : std_logic;
signal \N__37648\ : std_logic;
signal \N__37645\ : std_logic;
signal \N__37642\ : std_logic;
signal \N__37637\ : std_logic;
signal \N__37634\ : std_logic;
signal \N__37631\ : std_logic;
signal \N__37628\ : std_logic;
signal \N__37625\ : std_logic;
signal \N__37622\ : std_logic;
signal \N__37619\ : std_logic;
signal \N__37616\ : std_logic;
signal \N__37613\ : std_logic;
signal \N__37610\ : std_logic;
signal \N__37607\ : std_logic;
signal \N__37604\ : std_logic;
signal \N__37601\ : std_logic;
signal \N__37598\ : std_logic;
signal \N__37595\ : std_logic;
signal \N__37594\ : std_logic;
signal \N__37591\ : std_logic;
signal \N__37588\ : std_logic;
signal \N__37585\ : std_logic;
signal \N__37580\ : std_logic;
signal \N__37577\ : std_logic;
signal \N__37574\ : std_logic;
signal \N__37571\ : std_logic;
signal \N__37570\ : std_logic;
signal \N__37567\ : std_logic;
signal \N__37564\ : std_logic;
signal \N__37561\ : std_logic;
signal \N__37556\ : std_logic;
signal \N__37553\ : std_logic;
signal \N__37550\ : std_logic;
signal \N__37547\ : std_logic;
signal \N__37544\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37538\ : std_logic;
signal \N__37535\ : std_logic;
signal \N__37534\ : std_logic;
signal \N__37531\ : std_logic;
signal \N__37528\ : std_logic;
signal \N__37525\ : std_logic;
signal \N__37520\ : std_logic;
signal \N__37517\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37511\ : std_logic;
signal \N__37508\ : std_logic;
signal \N__37505\ : std_logic;
signal \N__37502\ : std_logic;
signal \N__37499\ : std_logic;
signal \N__37496\ : std_logic;
signal \N__37495\ : std_logic;
signal \N__37492\ : std_logic;
signal \N__37489\ : std_logic;
signal \N__37486\ : std_logic;
signal \N__37481\ : std_logic;
signal \N__37478\ : std_logic;
signal \N__37475\ : std_logic;
signal \N__37472\ : std_logic;
signal \N__37469\ : std_logic;
signal \N__37466\ : std_logic;
signal \N__37463\ : std_logic;
signal \N__37460\ : std_logic;
signal \N__37457\ : std_logic;
signal \N__37454\ : std_logic;
signal \N__37451\ : std_logic;
signal \N__37448\ : std_logic;
signal \N__37445\ : std_logic;
signal \N__37442\ : std_logic;
signal \N__37439\ : std_logic;
signal \N__37436\ : std_logic;
signal \N__37433\ : std_logic;
signal \N__37430\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37421\ : std_logic;
signal \N__37418\ : std_logic;
signal \N__37415\ : std_logic;
signal \N__37412\ : std_logic;
signal \N__37409\ : std_logic;
signal \N__37406\ : std_logic;
signal \N__37403\ : std_logic;
signal \N__37400\ : std_logic;
signal \N__37399\ : std_logic;
signal \N__37396\ : std_logic;
signal \N__37393\ : std_logic;
signal \N__37390\ : std_logic;
signal \N__37385\ : std_logic;
signal \N__37382\ : std_logic;
signal \N__37379\ : std_logic;
signal \N__37376\ : std_logic;
signal \N__37373\ : std_logic;
signal \N__37370\ : std_logic;
signal \N__37369\ : std_logic;
signal \N__37366\ : std_logic;
signal \N__37363\ : std_logic;
signal \N__37360\ : std_logic;
signal \N__37355\ : std_logic;
signal \N__37352\ : std_logic;
signal \N__37349\ : std_logic;
signal \N__37346\ : std_logic;
signal \N__37343\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37334\ : std_logic;
signal \N__37331\ : std_logic;
signal \N__37328\ : std_logic;
signal \N__37327\ : std_logic;
signal \N__37324\ : std_logic;
signal \N__37321\ : std_logic;
signal \N__37318\ : std_logic;
signal \N__37313\ : std_logic;
signal \N__37310\ : std_logic;
signal \N__37307\ : std_logic;
signal \N__37306\ : std_logic;
signal \N__37303\ : std_logic;
signal \N__37300\ : std_logic;
signal \N__37297\ : std_logic;
signal \N__37292\ : std_logic;
signal \N__37289\ : std_logic;
signal \N__37286\ : std_logic;
signal \N__37283\ : std_logic;
signal \N__37280\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37274\ : std_logic;
signal \N__37271\ : std_logic;
signal \N__37268\ : std_logic;
signal \N__37265\ : std_logic;
signal \N__37262\ : std_logic;
signal \N__37259\ : std_logic;
signal \N__37258\ : std_logic;
signal \N__37255\ : std_logic;
signal \N__37252\ : std_logic;
signal \N__37249\ : std_logic;
signal \N__37244\ : std_logic;
signal \N__37241\ : std_logic;
signal \N__37238\ : std_logic;
signal \N__37235\ : std_logic;
signal \N__37232\ : std_logic;
signal \N__37229\ : std_logic;
signal \N__37226\ : std_logic;
signal \N__37223\ : std_logic;
signal \N__37220\ : std_logic;
signal \N__37219\ : std_logic;
signal \N__37216\ : std_logic;
signal \N__37213\ : std_logic;
signal \N__37210\ : std_logic;
signal \N__37205\ : std_logic;
signal \N__37202\ : std_logic;
signal \N__37199\ : std_logic;
signal \N__37196\ : std_logic;
signal \N__37193\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37184\ : std_logic;
signal \N__37181\ : std_logic;
signal \N__37180\ : std_logic;
signal \N__37177\ : std_logic;
signal \N__37174\ : std_logic;
signal \N__37171\ : std_logic;
signal \N__37166\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37157\ : std_logic;
signal \N__37156\ : std_logic;
signal \N__37153\ : std_logic;
signal \N__37152\ : std_logic;
signal \N__37149\ : std_logic;
signal \N__37146\ : std_logic;
signal \N__37143\ : std_logic;
signal \N__37136\ : std_logic;
signal \N__37133\ : std_logic;
signal \N__37130\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37121\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37117\ : std_logic;
signal \N__37116\ : std_logic;
signal \N__37113\ : std_logic;
signal \N__37110\ : std_logic;
signal \N__37107\ : std_logic;
signal \N__37104\ : std_logic;
signal \N__37101\ : std_logic;
signal \N__37094\ : std_logic;
signal \N__37091\ : std_logic;
signal \N__37088\ : std_logic;
signal \N__37087\ : std_logic;
signal \N__37084\ : std_logic;
signal \N__37081\ : std_logic;
signal \N__37078\ : std_logic;
signal \N__37073\ : std_logic;
signal \N__37070\ : std_logic;
signal \N__37067\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37061\ : std_logic;
signal \N__37058\ : std_logic;
signal \N__37055\ : std_logic;
signal \N__37054\ : std_logic;
signal \N__37051\ : std_logic;
signal \N__37048\ : std_logic;
signal \N__37045\ : std_logic;
signal \N__37040\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37034\ : std_logic;
signal \N__37031\ : std_logic;
signal \N__37028\ : std_logic;
signal \N__37027\ : std_logic;
signal \N__37024\ : std_logic;
signal \N__37021\ : std_logic;
signal \N__37018\ : std_logic;
signal \N__37013\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__37001\ : std_logic;
signal \N__36998\ : std_logic;
signal \N__36995\ : std_logic;
signal \N__36992\ : std_logic;
signal \N__36991\ : std_logic;
signal \N__36988\ : std_logic;
signal \N__36987\ : std_logic;
signal \N__36984\ : std_logic;
signal \N__36981\ : std_logic;
signal \N__36978\ : std_logic;
signal \N__36975\ : std_logic;
signal \N__36972\ : std_logic;
signal \N__36965\ : std_logic;
signal \N__36964\ : std_logic;
signal \N__36961\ : std_logic;
signal \N__36960\ : std_logic;
signal \N__36955\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36949\ : std_logic;
signal \N__36944\ : std_logic;
signal \N__36941\ : std_logic;
signal \N__36940\ : std_logic;
signal \N__36937\ : std_logic;
signal \N__36934\ : std_logic;
signal \N__36933\ : std_logic;
signal \N__36928\ : std_logic;
signal \N__36925\ : std_logic;
signal \N__36922\ : std_logic;
signal \N__36917\ : std_logic;
signal \N__36916\ : std_logic;
signal \N__36913\ : std_logic;
signal \N__36910\ : std_logic;
signal \N__36905\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36901\ : std_logic;
signal \N__36896\ : std_logic;
signal \N__36893\ : std_logic;
signal \N__36892\ : std_logic;
signal \N__36889\ : std_logic;
signal \N__36886\ : std_logic;
signal \N__36885\ : std_logic;
signal \N__36880\ : std_logic;
signal \N__36877\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36869\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36860\ : std_logic;
signal \N__36857\ : std_logic;
signal \N__36854\ : std_logic;
signal \N__36851\ : std_logic;
signal \N__36850\ : std_logic;
signal \N__36849\ : std_logic;
signal \N__36846\ : std_logic;
signal \N__36843\ : std_logic;
signal \N__36838\ : std_logic;
signal \N__36833\ : std_logic;
signal \N__36832\ : std_logic;
signal \N__36831\ : std_logic;
signal \N__36828\ : std_logic;
signal \N__36823\ : std_logic;
signal \N__36818\ : std_logic;
signal \N__36815\ : std_logic;
signal \N__36812\ : std_logic;
signal \N__36809\ : std_logic;
signal \N__36806\ : std_logic;
signal \N__36803\ : std_logic;
signal \N__36800\ : std_logic;
signal \N__36797\ : std_logic;
signal \N__36794\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36788\ : std_logic;
signal \N__36785\ : std_logic;
signal \N__36782\ : std_logic;
signal \N__36781\ : std_logic;
signal \N__36778\ : std_logic;
signal \N__36775\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36764\ : std_logic;
signal \N__36761\ : std_logic;
signal \N__36758\ : std_logic;
signal \N__36755\ : std_logic;
signal \N__36752\ : std_logic;
signal \N__36751\ : std_logic;
signal \N__36750\ : std_logic;
signal \N__36749\ : std_logic;
signal \N__36744\ : std_logic;
signal \N__36741\ : std_logic;
signal \N__36738\ : std_logic;
signal \N__36733\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36727\ : std_logic;
signal \N__36726\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36720\ : std_logic;
signal \N__36717\ : std_logic;
signal \N__36714\ : std_logic;
signal \N__36707\ : std_logic;
signal \N__36704\ : std_logic;
signal \N__36701\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36695\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36689\ : std_logic;
signal \N__36686\ : std_logic;
signal \N__36685\ : std_logic;
signal \N__36684\ : std_logic;
signal \N__36681\ : std_logic;
signal \N__36678\ : std_logic;
signal \N__36675\ : std_logic;
signal \N__36670\ : std_logic;
signal \N__36665\ : std_logic;
signal \N__36662\ : std_logic;
signal \N__36659\ : std_logic;
signal \N__36656\ : std_logic;
signal \N__36653\ : std_logic;
signal \N__36650\ : std_logic;
signal \N__36647\ : std_logic;
signal \N__36644\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36638\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36632\ : std_logic;
signal \N__36629\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36620\ : std_logic;
signal \N__36617\ : std_logic;
signal \N__36614\ : std_logic;
signal \N__36611\ : std_logic;
signal \N__36608\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36602\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36596\ : std_logic;
signal \N__36593\ : std_logic;
signal \N__36590\ : std_logic;
signal \N__36587\ : std_logic;
signal \N__36584\ : std_logic;
signal \N__36581\ : std_logic;
signal \N__36578\ : std_logic;
signal \N__36575\ : std_logic;
signal \N__36572\ : std_logic;
signal \N__36569\ : std_logic;
signal \N__36566\ : std_logic;
signal \N__36563\ : std_logic;
signal \N__36560\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36554\ : std_logic;
signal \N__36551\ : std_logic;
signal \N__36548\ : std_logic;
signal \N__36545\ : std_logic;
signal \N__36542\ : std_logic;
signal \N__36539\ : std_logic;
signal \N__36536\ : std_logic;
signal \N__36533\ : std_logic;
signal \N__36530\ : std_logic;
signal \N__36527\ : std_logic;
signal \N__36524\ : std_logic;
signal \N__36521\ : std_logic;
signal \N__36518\ : std_logic;
signal \N__36515\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36509\ : std_logic;
signal \N__36506\ : std_logic;
signal \N__36503\ : std_logic;
signal \N__36500\ : std_logic;
signal \N__36497\ : std_logic;
signal \N__36494\ : std_logic;
signal \N__36491\ : std_logic;
signal \N__36488\ : std_logic;
signal \N__36485\ : std_logic;
signal \N__36482\ : std_logic;
signal \N__36479\ : std_logic;
signal \N__36476\ : std_logic;
signal \N__36473\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36467\ : std_logic;
signal \N__36464\ : std_logic;
signal \N__36461\ : std_logic;
signal \N__36458\ : std_logic;
signal \N__36455\ : std_logic;
signal \N__36452\ : std_logic;
signal \N__36449\ : std_logic;
signal \N__36446\ : std_logic;
signal \N__36443\ : std_logic;
signal \N__36440\ : std_logic;
signal \N__36437\ : std_logic;
signal \N__36434\ : std_logic;
signal \N__36431\ : std_logic;
signal \N__36428\ : std_logic;
signal \N__36425\ : std_logic;
signal \N__36422\ : std_logic;
signal \N__36419\ : std_logic;
signal \N__36416\ : std_logic;
signal \N__36413\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36404\ : std_logic;
signal \N__36401\ : std_logic;
signal \N__36398\ : std_logic;
signal \N__36395\ : std_logic;
signal \N__36392\ : std_logic;
signal \N__36389\ : std_logic;
signal \N__36386\ : std_logic;
signal \N__36383\ : std_logic;
signal \N__36380\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36374\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36368\ : std_logic;
signal \N__36365\ : std_logic;
signal \N__36362\ : std_logic;
signal \N__36359\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36353\ : std_logic;
signal \N__36350\ : std_logic;
signal \N__36347\ : std_logic;
signal \N__36344\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36335\ : std_logic;
signal \N__36332\ : std_logic;
signal \N__36329\ : std_logic;
signal \N__36326\ : std_logic;
signal \N__36323\ : std_logic;
signal \N__36320\ : std_logic;
signal \N__36317\ : std_logic;
signal \N__36314\ : std_logic;
signal \N__36311\ : std_logic;
signal \N__36308\ : std_logic;
signal \N__36305\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36299\ : std_logic;
signal \N__36296\ : std_logic;
signal \N__36293\ : std_logic;
signal \N__36290\ : std_logic;
signal \N__36287\ : std_logic;
signal \N__36284\ : std_logic;
signal \N__36281\ : std_logic;
signal \N__36278\ : std_logic;
signal \N__36277\ : std_logic;
signal \N__36276\ : std_logic;
signal \N__36273\ : std_logic;
signal \N__36268\ : std_logic;
signal \N__36263\ : std_logic;
signal \N__36260\ : std_logic;
signal \N__36257\ : std_logic;
signal \N__36254\ : std_logic;
signal \N__36251\ : std_logic;
signal \N__36248\ : std_logic;
signal \N__36247\ : std_logic;
signal \N__36246\ : std_logic;
signal \N__36243\ : std_logic;
signal \N__36238\ : std_logic;
signal \N__36233\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36229\ : std_logic;
signal \N__36228\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36226\ : std_logic;
signal \N__36225\ : std_logic;
signal \N__36224\ : std_logic;
signal \N__36223\ : std_logic;
signal \N__36222\ : std_logic;
signal \N__36221\ : std_logic;
signal \N__36220\ : std_logic;
signal \N__36219\ : std_logic;
signal \N__36218\ : std_logic;
signal \N__36217\ : std_logic;
signal \N__36216\ : std_logic;
signal \N__36213\ : std_logic;
signal \N__36206\ : std_logic;
signal \N__36197\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36195\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36186\ : std_logic;
signal \N__36177\ : std_logic;
signal \N__36176\ : std_logic;
signal \N__36175\ : std_logic;
signal \N__36174\ : std_logic;
signal \N__36173\ : std_logic;
signal \N__36170\ : std_logic;
signal \N__36169\ : std_logic;
signal \N__36168\ : std_logic;
signal \N__36167\ : std_logic;
signal \N__36166\ : std_logic;
signal \N__36165\ : std_logic;
signal \N__36164\ : std_logic;
signal \N__36163\ : std_logic;
signal \N__36162\ : std_logic;
signal \N__36161\ : std_logic;
signal \N__36158\ : std_logic;
signal \N__36155\ : std_logic;
signal \N__36146\ : std_logic;
signal \N__36141\ : std_logic;
signal \N__36132\ : std_logic;
signal \N__36129\ : std_logic;
signal \N__36126\ : std_logic;
signal \N__36117\ : std_logic;
signal \N__36108\ : std_logic;
signal \N__36097\ : std_logic;
signal \N__36094\ : std_logic;
signal \N__36087\ : std_logic;
signal \N__36084\ : std_logic;
signal \N__36081\ : std_logic;
signal \N__36078\ : std_logic;
signal \N__36075\ : std_logic;
signal \N__36072\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36061\ : std_logic;
signal \N__36058\ : std_logic;
signal \N__36057\ : std_logic;
signal \N__36054\ : std_logic;
signal \N__36049\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36038\ : std_logic;
signal \N__36035\ : std_logic;
signal \N__36032\ : std_logic;
signal \N__36029\ : std_logic;
signal \N__36026\ : std_logic;
signal \N__36023\ : std_logic;
signal \N__36022\ : std_logic;
signal \N__36021\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36010\ : std_logic;
signal \N__36005\ : std_logic;
signal \N__36002\ : std_logic;
signal \N__36001\ : std_logic;
signal \N__36000\ : std_logic;
signal \N__35997\ : std_logic;
signal \N__35994\ : std_logic;
signal \N__35989\ : std_logic;
signal \N__35984\ : std_logic;
signal \N__35981\ : std_logic;
signal \N__35980\ : std_logic;
signal \N__35977\ : std_logic;
signal \N__35976\ : std_logic;
signal \N__35973\ : std_logic;
signal \N__35968\ : std_logic;
signal \N__35963\ : std_logic;
signal \N__35960\ : std_logic;
signal \N__35957\ : std_logic;
signal \N__35954\ : std_logic;
signal \N__35951\ : std_logic;
signal \N__35948\ : std_logic;
signal \N__35945\ : std_logic;
signal \N__35942\ : std_logic;
signal \N__35939\ : std_logic;
signal \N__35936\ : std_logic;
signal \N__35933\ : std_logic;
signal \N__35932\ : std_logic;
signal \N__35929\ : std_logic;
signal \N__35928\ : std_logic;
signal \N__35925\ : std_logic;
signal \N__35922\ : std_logic;
signal \N__35919\ : std_logic;
signal \N__35912\ : std_logic;
signal \N__35909\ : std_logic;
signal \N__35906\ : std_logic;
signal \N__35903\ : std_logic;
signal \N__35900\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35894\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35885\ : std_logic;
signal \N__35882\ : std_logic;
signal \N__35879\ : std_logic;
signal \N__35876\ : std_logic;
signal \N__35873\ : std_logic;
signal \N__35870\ : std_logic;
signal \N__35867\ : std_logic;
signal \N__35864\ : std_logic;
signal \N__35861\ : std_logic;
signal \N__35860\ : std_logic;
signal \N__35857\ : std_logic;
signal \N__35854\ : std_logic;
signal \N__35853\ : std_logic;
signal \N__35852\ : std_logic;
signal \N__35847\ : std_logic;
signal \N__35844\ : std_logic;
signal \N__35841\ : std_logic;
signal \N__35838\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35827\ : std_logic;
signal \N__35826\ : std_logic;
signal \N__35823\ : std_logic;
signal \N__35818\ : std_logic;
signal \N__35817\ : std_logic;
signal \N__35812\ : std_logic;
signal \N__35809\ : std_logic;
signal \N__35806\ : std_logic;
signal \N__35801\ : std_logic;
signal \N__35798\ : std_logic;
signal \N__35797\ : std_logic;
signal \N__35796\ : std_logic;
signal \N__35793\ : std_logic;
signal \N__35790\ : std_logic;
signal \N__35787\ : std_logic;
signal \N__35782\ : std_logic;
signal \N__35777\ : std_logic;
signal \N__35774\ : std_logic;
signal \N__35773\ : std_logic;
signal \N__35770\ : std_logic;
signal \N__35769\ : std_logic;
signal \N__35766\ : std_logic;
signal \N__35763\ : std_logic;
signal \N__35760\ : std_logic;
signal \N__35753\ : std_logic;
signal \N__35750\ : std_logic;
signal \N__35747\ : std_logic;
signal \N__35744\ : std_logic;
signal \N__35741\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35735\ : std_logic;
signal \N__35732\ : std_logic;
signal \N__35729\ : std_logic;
signal \N__35726\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35714\ : std_logic;
signal \N__35711\ : std_logic;
signal \N__35708\ : std_logic;
signal \N__35705\ : std_logic;
signal \N__35702\ : std_logic;
signal \N__35699\ : std_logic;
signal \N__35696\ : std_logic;
signal \N__35693\ : std_logic;
signal \N__35690\ : std_logic;
signal \N__35687\ : std_logic;
signal \N__35684\ : std_logic;
signal \N__35681\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35677\ : std_logic;
signal \N__35676\ : std_logic;
signal \N__35673\ : std_logic;
signal \N__35670\ : std_logic;
signal \N__35667\ : std_logic;
signal \N__35660\ : std_logic;
signal \N__35657\ : std_logic;
signal \N__35654\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35648\ : std_logic;
signal \N__35645\ : std_logic;
signal \N__35642\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35638\ : std_logic;
signal \N__35635\ : std_logic;
signal \N__35630\ : std_logic;
signal \N__35629\ : std_logic;
signal \N__35628\ : std_logic;
signal \N__35625\ : std_logic;
signal \N__35624\ : std_logic;
signal \N__35623\ : std_logic;
signal \N__35618\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35610\ : std_logic;
signal \N__35603\ : std_logic;
signal \N__35602\ : std_logic;
signal \N__35601\ : std_logic;
signal \N__35598\ : std_logic;
signal \N__35593\ : std_logic;
signal \N__35588\ : std_logic;
signal \N__35585\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35579\ : std_logic;
signal \N__35576\ : std_logic;
signal \N__35575\ : std_logic;
signal \N__35574\ : std_logic;
signal \N__35571\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35565\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35555\ : std_logic;
signal \N__35552\ : std_logic;
signal \N__35549\ : std_logic;
signal \N__35546\ : std_logic;
signal \N__35543\ : std_logic;
signal \N__35540\ : std_logic;
signal \N__35537\ : std_logic;
signal \N__35534\ : std_logic;
signal \N__35531\ : std_logic;
signal \N__35528\ : std_logic;
signal \N__35525\ : std_logic;
signal \N__35522\ : std_logic;
signal \N__35519\ : std_logic;
signal \N__35516\ : std_logic;
signal \N__35513\ : std_logic;
signal \N__35510\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35504\ : std_logic;
signal \N__35501\ : std_logic;
signal \N__35498\ : std_logic;
signal \N__35495\ : std_logic;
signal \N__35492\ : std_logic;
signal \N__35489\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35477\ : std_logic;
signal \N__35474\ : std_logic;
signal \N__35471\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35465\ : std_logic;
signal \N__35462\ : std_logic;
signal \N__35459\ : std_logic;
signal \N__35456\ : std_logic;
signal \N__35453\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35447\ : std_logic;
signal \N__35444\ : std_logic;
signal \N__35441\ : std_logic;
signal \N__35438\ : std_logic;
signal \N__35435\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35420\ : std_logic;
signal \N__35417\ : std_logic;
signal \N__35414\ : std_logic;
signal \N__35411\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35402\ : std_logic;
signal \N__35399\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35393\ : std_logic;
signal \N__35390\ : std_logic;
signal \N__35387\ : std_logic;
signal \N__35384\ : std_logic;
signal \N__35381\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35363\ : std_logic;
signal \N__35360\ : std_logic;
signal \N__35357\ : std_logic;
signal \N__35354\ : std_logic;
signal \N__35351\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35342\ : std_logic;
signal \N__35339\ : std_logic;
signal \N__35336\ : std_logic;
signal \N__35333\ : std_logic;
signal \N__35330\ : std_logic;
signal \N__35327\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35294\ : std_logic;
signal \N__35291\ : std_logic;
signal \N__35288\ : std_logic;
signal \N__35285\ : std_logic;
signal \N__35282\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35267\ : std_logic;
signal \N__35264\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35258\ : std_logic;
signal \N__35255\ : std_logic;
signal \N__35252\ : std_logic;
signal \N__35251\ : std_logic;
signal \N__35246\ : std_logic;
signal \N__35243\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35239\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35231\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35227\ : std_logic;
signal \N__35222\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35213\ : std_logic;
signal \N__35210\ : std_logic;
signal \N__35207\ : std_logic;
signal \N__35204\ : std_logic;
signal \N__35201\ : std_logic;
signal \N__35198\ : std_logic;
signal \N__35195\ : std_logic;
signal \N__35192\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35186\ : std_logic;
signal \N__35183\ : std_logic;
signal \N__35180\ : std_logic;
signal \N__35179\ : std_logic;
signal \N__35174\ : std_logic;
signal \N__35171\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35169\ : std_logic;
signal \N__35168\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35164\ : std_logic;
signal \N__35161\ : std_logic;
signal \N__35158\ : std_logic;
signal \N__35155\ : std_logic;
signal \N__35152\ : std_logic;
signal \N__35149\ : std_logic;
signal \N__35146\ : std_logic;
signal \N__35135\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35131\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35127\ : std_logic;
signal \N__35124\ : std_logic;
signal \N__35121\ : std_logic;
signal \N__35118\ : std_logic;
signal \N__35111\ : std_logic;
signal \N__35108\ : std_logic;
signal \N__35107\ : std_logic;
signal \N__35104\ : std_logic;
signal \N__35101\ : std_logic;
signal \N__35096\ : std_logic;
signal \N__35093\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35091\ : std_logic;
signal \N__35088\ : std_logic;
signal \N__35083\ : std_logic;
signal \N__35078\ : std_logic;
signal \N__35075\ : std_logic;
signal \N__35074\ : std_logic;
signal \N__35071\ : std_logic;
signal \N__35068\ : std_logic;
signal \N__35067\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35061\ : std_logic;
signal \N__35056\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35048\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35037\ : std_logic;
signal \N__35036\ : std_logic;
signal \N__35031\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35021\ : std_logic;
signal \N__35020\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35013\ : std_logic;
signal \N__35012\ : std_logic;
signal \N__35011\ : std_logic;
signal \N__35008\ : std_logic;
signal \N__35005\ : std_logic;
signal \N__35000\ : std_logic;
signal \N__34997\ : std_logic;
signal \N__34988\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34986\ : std_logic;
signal \N__34983\ : std_logic;
signal \N__34980\ : std_logic;
signal \N__34977\ : std_logic;
signal \N__34974\ : std_logic;
signal \N__34969\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34961\ : std_logic;
signal \N__34958\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34954\ : std_logic;
signal \N__34949\ : std_logic;
signal \N__34948\ : std_logic;
signal \N__34945\ : std_logic;
signal \N__34942\ : std_logic;
signal \N__34939\ : std_logic;
signal \N__34938\ : std_logic;
signal \N__34935\ : std_logic;
signal \N__34932\ : std_logic;
signal \N__34929\ : std_logic;
signal \N__34922\ : std_logic;
signal \N__34921\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34910\ : std_logic;
signal \N__34909\ : std_logic;
signal \N__34906\ : std_logic;
signal \N__34905\ : std_logic;
signal \N__34902\ : std_logic;
signal \N__34899\ : std_logic;
signal \N__34896\ : std_logic;
signal \N__34889\ : std_logic;
signal \N__34886\ : std_logic;
signal \N__34885\ : std_logic;
signal \N__34882\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34875\ : std_logic;
signal \N__34872\ : std_logic;
signal \N__34871\ : std_logic;
signal \N__34868\ : std_logic;
signal \N__34863\ : std_logic;
signal \N__34860\ : std_logic;
signal \N__34853\ : std_logic;
signal \N__34850\ : std_logic;
signal \N__34847\ : std_logic;
signal \N__34844\ : std_logic;
signal \N__34843\ : std_logic;
signal \N__34842\ : std_logic;
signal \N__34841\ : std_logic;
signal \N__34840\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34838\ : std_logic;
signal \N__34837\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34835\ : std_logic;
signal \N__34834\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34832\ : std_logic;
signal \N__34831\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34829\ : std_logic;
signal \N__34828\ : std_logic;
signal \N__34825\ : std_logic;
signal \N__34818\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34816\ : std_logic;
signal \N__34815\ : std_logic;
signal \N__34810\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34786\ : std_logic;
signal \N__34781\ : std_logic;
signal \N__34780\ : std_logic;
signal \N__34779\ : std_logic;
signal \N__34778\ : std_logic;
signal \N__34777\ : std_logic;
signal \N__34776\ : std_logic;
signal \N__34775\ : std_logic;
signal \N__34774\ : std_logic;
signal \N__34773\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34770\ : std_logic;
signal \N__34769\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34767\ : std_logic;
signal \N__34766\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34762\ : std_logic;
signal \N__34759\ : std_logic;
signal \N__34758\ : std_logic;
signal \N__34757\ : std_logic;
signal \N__34756\ : std_logic;
signal \N__34755\ : std_logic;
signal \N__34754\ : std_logic;
signal \N__34753\ : std_logic;
signal \N__34752\ : std_logic;
signal \N__34751\ : std_logic;
signal \N__34750\ : std_logic;
signal \N__34749\ : std_logic;
signal \N__34748\ : std_logic;
signal \N__34747\ : std_logic;
signal \N__34746\ : std_logic;
signal \N__34743\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34741\ : std_logic;
signal \N__34740\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34738\ : std_logic;
signal \N__34737\ : std_logic;
signal \N__34736\ : std_logic;
signal \N__34735\ : std_logic;
signal \N__34734\ : std_logic;
signal \N__34733\ : std_logic;
signal \N__34732\ : std_logic;
signal \N__34723\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34711\ : std_logic;
signal \N__34710\ : std_logic;
signal \N__34709\ : std_logic;
signal \N__34704\ : std_logic;
signal \N__34691\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34685\ : std_logic;
signal \N__34684\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34674\ : std_logic;
signal \N__34673\ : std_logic;
signal \N__34672\ : std_logic;
signal \N__34671\ : std_logic;
signal \N__34670\ : std_logic;
signal \N__34669\ : std_logic;
signal \N__34668\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34666\ : std_logic;
signal \N__34663\ : std_logic;
signal \N__34660\ : std_logic;
signal \N__34647\ : std_logic;
signal \N__34636\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34623\ : std_logic;
signal \N__34620\ : std_logic;
signal \N__34615\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34613\ : std_logic;
signal \N__34612\ : std_logic;
signal \N__34611\ : std_logic;
signal \N__34610\ : std_logic;
signal \N__34609\ : std_logic;
signal \N__34608\ : std_logic;
signal \N__34607\ : std_logic;
signal \N__34606\ : std_logic;
signal \N__34605\ : std_logic;
signal \N__34604\ : std_logic;
signal \N__34603\ : std_logic;
signal \N__34602\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34600\ : std_logic;
signal \N__34599\ : std_logic;
signal \N__34590\ : std_logic;
signal \N__34585\ : std_logic;
signal \N__34582\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34578\ : std_logic;
signal \N__34575\ : std_logic;
signal \N__34568\ : std_logic;
signal \N__34557\ : std_logic;
signal \N__34554\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34530\ : std_logic;
signal \N__34525\ : std_logic;
signal \N__34520\ : std_logic;
signal \N__34517\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34507\ : std_logic;
signal \N__34504\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34486\ : std_logic;
signal \N__34475\ : std_logic;
signal \N__34472\ : std_logic;
signal \N__34469\ : std_logic;
signal \N__34464\ : std_logic;
signal \N__34459\ : std_logic;
signal \N__34452\ : std_logic;
signal \N__34435\ : std_logic;
signal \N__34412\ : std_logic;
signal \N__34409\ : std_logic;
signal \N__34408\ : std_logic;
signal \N__34405\ : std_logic;
signal \N__34404\ : std_logic;
signal \N__34401\ : std_logic;
signal \N__34398\ : std_logic;
signal \N__34395\ : std_logic;
signal \N__34390\ : std_logic;
signal \N__34385\ : std_logic;
signal \N__34384\ : std_logic;
signal \N__34381\ : std_logic;
signal \N__34378\ : std_logic;
signal \N__34375\ : std_logic;
signal \N__34374\ : std_logic;
signal \N__34371\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34365\ : std_logic;
signal \N__34364\ : std_logic;
signal \N__34361\ : std_logic;
signal \N__34356\ : std_logic;
signal \N__34353\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34340\ : std_logic;
signal \N__34337\ : std_logic;
signal \N__34334\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34332\ : std_logic;
signal \N__34331\ : std_logic;
signal \N__34330\ : std_logic;
signal \N__34329\ : std_logic;
signal \N__34328\ : std_logic;
signal \N__34327\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34325\ : std_logic;
signal \N__34324\ : std_logic;
signal \N__34323\ : std_logic;
signal \N__34322\ : std_logic;
signal \N__34321\ : std_logic;
signal \N__34320\ : std_logic;
signal \N__34319\ : std_logic;
signal \N__34318\ : std_logic;
signal \N__34317\ : std_logic;
signal \N__34316\ : std_logic;
signal \N__34313\ : std_logic;
signal \N__34312\ : std_logic;
signal \N__34311\ : std_logic;
signal \N__34310\ : std_logic;
signal \N__34309\ : std_logic;
signal \N__34302\ : std_logic;
signal \N__34293\ : std_logic;
signal \N__34284\ : std_logic;
signal \N__34281\ : std_logic;
signal \N__34280\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34276\ : std_logic;
signal \N__34267\ : std_logic;
signal \N__34264\ : std_logic;
signal \N__34263\ : std_logic;
signal \N__34262\ : std_logic;
signal \N__34261\ : std_logic;
signal \N__34258\ : std_logic;
signal \N__34255\ : std_logic;
signal \N__34254\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34238\ : std_logic;
signal \N__34237\ : std_logic;
signal \N__34236\ : std_logic;
signal \N__34235\ : std_logic;
signal \N__34234\ : std_logic;
signal \N__34233\ : std_logic;
signal \N__34232\ : std_logic;
signal \N__34231\ : std_logic;
signal \N__34230\ : std_logic;
signal \N__34229\ : std_logic;
signal \N__34228\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34226\ : std_logic;
signal \N__34223\ : std_logic;
signal \N__34220\ : std_logic;
signal \N__34217\ : std_logic;
signal \N__34212\ : std_logic;
signal \N__34209\ : std_logic;
signal \N__34206\ : std_logic;
signal \N__34203\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34180\ : std_logic;
signal \N__34171\ : std_logic;
signal \N__34162\ : std_logic;
signal \N__34159\ : std_logic;
signal \N__34154\ : std_logic;
signal \N__34151\ : std_logic;
signal \N__34148\ : std_logic;
signal \N__34145\ : std_logic;
signal \N__34142\ : std_logic;
signal \N__34141\ : std_logic;
signal \N__34138\ : std_logic;
signal \N__34135\ : std_logic;
signal \N__34132\ : std_logic;
signal \N__34121\ : std_logic;
signal \N__34118\ : std_logic;
signal \N__34115\ : std_logic;
signal \N__34110\ : std_logic;
signal \N__34107\ : std_logic;
signal \N__34104\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34094\ : std_logic;
signal \N__34089\ : std_logic;
signal \N__34076\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34070\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34058\ : std_logic;
signal \N__34055\ : std_logic;
signal \N__34054\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34043\ : std_logic;
signal \N__34040\ : std_logic;
signal \N__34039\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34035\ : std_logic;
signal \N__34032\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34026\ : std_logic;
signal \N__34023\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34019\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34008\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__33998\ : std_logic;
signal \N__33997\ : std_logic;
signal \N__33996\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33990\ : std_logic;
signal \N__33987\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33981\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33971\ : std_logic;
signal \N__33968\ : std_logic;
signal \N__33965\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33959\ : std_logic;
signal \N__33956\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33954\ : std_logic;
signal \N__33951\ : std_logic;
signal \N__33946\ : std_logic;
signal \N__33941\ : std_logic;
signal \N__33938\ : std_logic;
signal \N__33937\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33931\ : std_logic;
signal \N__33928\ : std_logic;
signal \N__33925\ : std_logic;
signal \N__33920\ : std_logic;
signal \N__33917\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33908\ : std_logic;
signal \N__33905\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33901\ : std_logic;
signal \N__33900\ : std_logic;
signal \N__33897\ : std_logic;
signal \N__33894\ : std_logic;
signal \N__33891\ : std_logic;
signal \N__33888\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33878\ : std_logic;
signal \N__33875\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33870\ : std_logic;
signal \N__33867\ : std_logic;
signal \N__33864\ : std_logic;
signal \N__33861\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33857\ : std_logic;
signal \N__33852\ : std_logic;
signal \N__33849\ : std_logic;
signal \N__33842\ : std_logic;
signal \N__33839\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33833\ : std_logic;
signal \N__33830\ : std_logic;
signal \N__33827\ : std_logic;
signal \N__33824\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33820\ : std_logic;
signal \N__33817\ : std_logic;
signal \N__33812\ : std_logic;
signal \N__33809\ : std_logic;
signal \N__33806\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33800\ : std_logic;
signal \N__33797\ : std_logic;
signal \N__33794\ : std_logic;
signal \N__33791\ : std_logic;
signal \N__33788\ : std_logic;
signal \N__33785\ : std_logic;
signal \N__33782\ : std_logic;
signal \N__33779\ : std_logic;
signal \N__33776\ : std_logic;
signal \N__33773\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33767\ : std_logic;
signal \N__33764\ : std_logic;
signal \N__33761\ : std_logic;
signal \N__33758\ : std_logic;
signal \N__33755\ : std_logic;
signal \N__33752\ : std_logic;
signal \N__33749\ : std_logic;
signal \N__33746\ : std_logic;
signal \N__33743\ : std_logic;
signal \N__33740\ : std_logic;
signal \N__33737\ : std_logic;
signal \N__33734\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33728\ : std_logic;
signal \N__33725\ : std_logic;
signal \N__33722\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33710\ : std_logic;
signal \N__33707\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33701\ : std_logic;
signal \N__33698\ : std_logic;
signal \N__33695\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33677\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33665\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33653\ : std_logic;
signal \N__33650\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33638\ : std_logic;
signal \N__33635\ : std_logic;
signal \N__33632\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33623\ : std_logic;
signal \N__33620\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33614\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33599\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33593\ : std_logic;
signal \N__33590\ : std_logic;
signal \N__33587\ : std_logic;
signal \N__33584\ : std_logic;
signal \N__33581\ : std_logic;
signal \N__33578\ : std_logic;
signal \N__33575\ : std_logic;
signal \N__33572\ : std_logic;
signal \N__33571\ : std_logic;
signal \N__33568\ : std_logic;
signal \N__33565\ : std_logic;
signal \N__33560\ : std_logic;
signal \N__33557\ : std_logic;
signal \N__33554\ : std_logic;
signal \N__33553\ : std_logic;
signal \N__33550\ : std_logic;
signal \N__33547\ : std_logic;
signal \N__33546\ : std_logic;
signal \N__33545\ : std_logic;
signal \N__33540\ : std_logic;
signal \N__33535\ : std_logic;
signal \N__33532\ : std_logic;
signal \N__33529\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33520\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33511\ : std_logic;
signal \N__33506\ : std_logic;
signal \N__33503\ : std_logic;
signal \N__33500\ : std_logic;
signal \N__33497\ : std_logic;
signal \N__33494\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33488\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33482\ : std_logic;
signal \N__33479\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33473\ : std_logic;
signal \N__33470\ : std_logic;
signal \N__33469\ : std_logic;
signal \N__33468\ : std_logic;
signal \N__33461\ : std_logic;
signal \N__33458\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33454\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33450\ : std_logic;
signal \N__33447\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33437\ : std_logic;
signal \N__33434\ : std_logic;
signal \N__33431\ : std_logic;
signal \N__33428\ : std_logic;
signal \N__33427\ : std_logic;
signal \N__33424\ : std_logic;
signal \N__33421\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33412\ : std_logic;
signal \N__33411\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33405\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33399\ : std_logic;
signal \N__33396\ : std_logic;
signal \N__33393\ : std_logic;
signal \N__33390\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33381\ : std_logic;
signal \N__33374\ : std_logic;
signal \N__33371\ : std_logic;
signal \N__33368\ : std_logic;
signal \N__33365\ : std_logic;
signal \N__33362\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33355\ : std_logic;
signal \N__33354\ : std_logic;
signal \N__33349\ : std_logic;
signal \N__33346\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33338\ : std_logic;
signal \N__33335\ : std_logic;
signal \N__33334\ : std_logic;
signal \N__33329\ : std_logic;
signal \N__33326\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33324\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33316\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33308\ : std_logic;
signal \N__33305\ : std_logic;
signal \N__33302\ : std_logic;
signal \N__33299\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33292\ : std_logic;
signal \N__33289\ : std_logic;
signal \N__33286\ : std_logic;
signal \N__33281\ : std_logic;
signal \N__33278\ : std_logic;
signal \N__33277\ : std_logic;
signal \N__33276\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33267\ : std_logic;
signal \N__33264\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33255\ : std_logic;
signal \N__33252\ : std_logic;
signal \N__33249\ : std_logic;
signal \N__33242\ : std_logic;
signal \N__33239\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33233\ : std_logic;
signal \N__33230\ : std_logic;
signal \N__33227\ : std_logic;
signal \N__33226\ : std_logic;
signal \N__33223\ : std_logic;
signal \N__33220\ : std_logic;
signal \N__33217\ : std_logic;
signal \N__33212\ : std_logic;
signal \N__33209\ : std_logic;
signal \N__33206\ : std_logic;
signal \N__33203\ : std_logic;
signal \N__33200\ : std_logic;
signal \N__33197\ : std_logic;
signal \N__33196\ : std_logic;
signal \N__33195\ : std_logic;
signal \N__33192\ : std_logic;
signal \N__33189\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33179\ : std_logic;
signal \N__33176\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33174\ : std_logic;
signal \N__33171\ : std_logic;
signal \N__33168\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33158\ : std_logic;
signal \N__33155\ : std_logic;
signal \N__33154\ : std_logic;
signal \N__33153\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33145\ : std_logic;
signal \N__33142\ : std_logic;
signal \N__33137\ : std_logic;
signal \N__33134\ : std_logic;
signal \N__33133\ : std_logic;
signal \N__33132\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33113\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33111\ : std_logic;
signal \N__33108\ : std_logic;
signal \N__33105\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33099\ : std_logic;
signal \N__33096\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33086\ : std_logic;
signal \N__33083\ : std_logic;
signal \N__33080\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33075\ : std_logic;
signal \N__33072\ : std_logic;
signal \N__33069\ : std_logic;
signal \N__33066\ : std_logic;
signal \N__33059\ : std_logic;
signal \N__33056\ : std_logic;
signal \N__33055\ : std_logic;
signal \N__33052\ : std_logic;
signal \N__33049\ : std_logic;
signal \N__33046\ : std_logic;
signal \N__33041\ : std_logic;
signal \N__33038\ : std_logic;
signal \N__33037\ : std_logic;
signal \N__33036\ : std_logic;
signal \N__33033\ : std_logic;
signal \N__33028\ : std_logic;
signal \N__33023\ : std_logic;
signal \N__33022\ : std_logic;
signal \N__33019\ : std_logic;
signal \N__33016\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__33002\ : std_logic;
signal \N__32999\ : std_logic;
signal \N__32996\ : std_logic;
signal \N__32993\ : std_logic;
signal \N__32992\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32980\ : std_logic;
signal \N__32977\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32969\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32965\ : std_logic;
signal \N__32964\ : std_logic;
signal \N__32959\ : std_logic;
signal \N__32956\ : std_logic;
signal \N__32953\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32944\ : std_logic;
signal \N__32941\ : std_logic;
signal \N__32940\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32929\ : std_logic;
signal \N__32924\ : std_logic;
signal \N__32921\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32919\ : std_logic;
signal \N__32914\ : std_logic;
signal \N__32911\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32903\ : std_logic;
signal \N__32900\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32890\ : std_logic;
signal \N__32887\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32879\ : std_logic;
signal \N__32878\ : std_logic;
signal \N__32877\ : std_logic;
signal \N__32872\ : std_logic;
signal \N__32869\ : std_logic;
signal \N__32866\ : std_logic;
signal \N__32861\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32855\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32851\ : std_logic;
signal \N__32848\ : std_logic;
signal \N__32845\ : std_logic;
signal \N__32840\ : std_logic;
signal \N__32837\ : std_logic;
signal \N__32836\ : std_logic;
signal \N__32833\ : std_logic;
signal \N__32830\ : std_logic;
signal \N__32825\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32821\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32815\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32806\ : std_logic;
signal \N__32803\ : std_logic;
signal \N__32800\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32792\ : std_logic;
signal \N__32791\ : std_logic;
signal \N__32788\ : std_logic;
signal \N__32785\ : std_logic;
signal \N__32780\ : std_logic;
signal \N__32777\ : std_logic;
signal \N__32776\ : std_logic;
signal \N__32773\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32761\ : std_logic;
signal \N__32758\ : std_logic;
signal \N__32755\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32737\ : std_logic;
signal \N__32734\ : std_logic;
signal \N__32733\ : std_logic;
signal \N__32730\ : std_logic;
signal \N__32727\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32714\ : std_logic;
signal \N__32713\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32706\ : std_logic;
signal \N__32703\ : std_logic;
signal \N__32700\ : std_logic;
signal \N__32697\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32680\ : std_logic;
signal \N__32677\ : std_logic;
signal \N__32674\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32663\ : std_logic;
signal \N__32662\ : std_logic;
signal \N__32659\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32651\ : std_logic;
signal \N__32648\ : std_logic;
signal \N__32647\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32641\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32633\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32629\ : std_logic;
signal \N__32626\ : std_logic;
signal \N__32621\ : std_logic;
signal \N__32618\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32614\ : std_logic;
signal \N__32611\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32584\ : std_logic;
signal \N__32581\ : std_logic;
signal \N__32576\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32564\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32558\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32552\ : std_logic;
signal \N__32551\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32539\ : std_logic;
signal \N__32536\ : std_logic;
signal \N__32533\ : std_logic;
signal \N__32530\ : std_logic;
signal \N__32527\ : std_logic;
signal \N__32522\ : std_logic;
signal \N__32521\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32510\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32506\ : std_logic;
signal \N__32505\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32502\ : std_logic;
signal \N__32501\ : std_logic;
signal \N__32498\ : std_logic;
signal \N__32491\ : std_logic;
signal \N__32484\ : std_logic;
signal \N__32477\ : std_logic;
signal \N__32474\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32470\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32468\ : std_logic;
signal \N__32467\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32464\ : std_logic;
signal \N__32463\ : std_logic;
signal \N__32462\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32459\ : std_logic;
signal \N__32458\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32440\ : std_logic;
signal \N__32425\ : std_logic;
signal \N__32424\ : std_logic;
signal \N__32423\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32411\ : std_logic;
signal \N__32410\ : std_logic;
signal \N__32409\ : std_logic;
signal \N__32408\ : std_logic;
signal \N__32407\ : std_logic;
signal \N__32406\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32400\ : std_logic;
signal \N__32397\ : std_logic;
signal \N__32396\ : std_logic;
signal \N__32395\ : std_logic;
signal \N__32394\ : std_logic;
signal \N__32393\ : std_logic;
signal \N__32392\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32390\ : std_logic;
signal \N__32389\ : std_logic;
signal \N__32386\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32374\ : std_logic;
signal \N__32371\ : std_logic;
signal \N__32368\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32347\ : std_logic;
signal \N__32344\ : std_logic;
signal \N__32339\ : std_logic;
signal \N__32336\ : std_logic;
signal \N__32333\ : std_logic;
signal \N__32330\ : std_logic;
signal \N__32321\ : std_logic;
signal \N__32318\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32300\ : std_logic;
signal \N__32297\ : std_logic;
signal \N__32294\ : std_logic;
signal \N__32291\ : std_logic;
signal \N__32288\ : std_logic;
signal \N__32285\ : std_logic;
signal \N__32282\ : std_logic;
signal \N__32279\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32273\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32264\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32258\ : std_logic;
signal \N__32257\ : std_logic;
signal \N__32254\ : std_logic;
signal \N__32253\ : std_logic;
signal \N__32250\ : std_logic;
signal \N__32247\ : std_logic;
signal \N__32244\ : std_logic;
signal \N__32243\ : std_logic;
signal \N__32240\ : std_logic;
signal \N__32235\ : std_logic;
signal \N__32232\ : std_logic;
signal \N__32229\ : std_logic;
signal \N__32226\ : std_logic;
signal \N__32219\ : std_logic;
signal \N__32216\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32209\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32199\ : std_logic;
signal \N__32196\ : std_logic;
signal \N__32193\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32179\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32175\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32150\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32144\ : std_logic;
signal \N__32141\ : std_logic;
signal \N__32138\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32126\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32114\ : std_logic;
signal \N__32111\ : std_logic;
signal \N__32108\ : std_logic;
signal \N__32105\ : std_logic;
signal \N__32102\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32093\ : std_logic;
signal \N__32090\ : std_logic;
signal \N__32087\ : std_logic;
signal \N__32084\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32078\ : std_logic;
signal \N__32075\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32065\ : std_logic;
signal \N__32062\ : std_logic;
signal \N__32059\ : std_logic;
signal \N__32054\ : std_logic;
signal \N__32051\ : std_logic;
signal \N__32048\ : std_logic;
signal \N__32045\ : std_logic;
signal \N__32042\ : std_logic;
signal \N__32039\ : std_logic;
signal \N__32036\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32021\ : std_logic;
signal \N__32018\ : std_logic;
signal \N__32015\ : std_logic;
signal \N__32012\ : std_logic;
signal \N__32009\ : std_logic;
signal \N__32006\ : std_logic;
signal \N__32003\ : std_logic;
signal \N__32000\ : std_logic;
signal \N__31997\ : std_logic;
signal \N__31994\ : std_logic;
signal \N__31991\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31955\ : std_logic;
signal \N__31952\ : std_logic;
signal \N__31949\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31940\ : std_logic;
signal \N__31937\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31931\ : std_logic;
signal \N__31928\ : std_logic;
signal \N__31925\ : std_logic;
signal \N__31922\ : std_logic;
signal \N__31919\ : std_logic;
signal \N__31916\ : std_logic;
signal \N__31913\ : std_logic;
signal \N__31910\ : std_logic;
signal \N__31907\ : std_logic;
signal \N__31904\ : std_logic;
signal \N__31901\ : std_logic;
signal \N__31898\ : std_logic;
signal \N__31895\ : std_logic;
signal \N__31892\ : std_logic;
signal \N__31889\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31883\ : std_logic;
signal \N__31880\ : std_logic;
signal \N__31877\ : std_logic;
signal \N__31874\ : std_logic;
signal \N__31871\ : std_logic;
signal \N__31868\ : std_logic;
signal \N__31865\ : std_logic;
signal \N__31862\ : std_logic;
signal \N__31859\ : std_logic;
signal \N__31856\ : std_logic;
signal \N__31853\ : std_logic;
signal \N__31850\ : std_logic;
signal \N__31847\ : std_logic;
signal \N__31844\ : std_logic;
signal \N__31841\ : std_logic;
signal \N__31838\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31832\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31823\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31817\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31811\ : std_logic;
signal \N__31808\ : std_logic;
signal \N__31805\ : std_logic;
signal \N__31802\ : std_logic;
signal \N__31799\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31793\ : std_logic;
signal \N__31790\ : std_logic;
signal \N__31787\ : std_logic;
signal \N__31786\ : std_logic;
signal \N__31783\ : std_logic;
signal \N__31780\ : std_logic;
signal \N__31775\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31767\ : std_logic;
signal \N__31764\ : std_logic;
signal \N__31761\ : std_logic;
signal \N__31758\ : std_logic;
signal \N__31755\ : std_logic;
signal \N__31748\ : std_logic;
signal \N__31745\ : std_logic;
signal \N__31742\ : std_logic;
signal \N__31739\ : std_logic;
signal \N__31736\ : std_logic;
signal \N__31733\ : std_logic;
signal \N__31730\ : std_logic;
signal \N__31727\ : std_logic;
signal \N__31724\ : std_logic;
signal \N__31721\ : std_logic;
signal \N__31718\ : std_logic;
signal \N__31715\ : std_logic;
signal \N__31712\ : std_logic;
signal \N__31709\ : std_logic;
signal \N__31706\ : std_logic;
signal \N__31703\ : std_logic;
signal \N__31700\ : std_logic;
signal \N__31697\ : std_logic;
signal \N__31694\ : std_logic;
signal \N__31691\ : std_logic;
signal \N__31688\ : std_logic;
signal \N__31685\ : std_logic;
signal \N__31682\ : std_logic;
signal \N__31679\ : std_logic;
signal \N__31676\ : std_logic;
signal \N__31673\ : std_logic;
signal \N__31670\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31661\ : std_logic;
signal \N__31658\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31652\ : std_logic;
signal \N__31649\ : std_logic;
signal \N__31646\ : std_logic;
signal \N__31645\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31639\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31633\ : std_logic;
signal \N__31630\ : std_logic;
signal \N__31627\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31616\ : std_logic;
signal \N__31615\ : std_logic;
signal \N__31614\ : std_logic;
signal \N__31611\ : std_logic;
signal \N__31608\ : std_logic;
signal \N__31605\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31599\ : std_logic;
signal \N__31596\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31587\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31581\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31573\ : std_logic;
signal \N__31570\ : std_logic;
signal \N__31569\ : std_logic;
signal \N__31566\ : std_logic;
signal \N__31565\ : std_logic;
signal \N__31562\ : std_logic;
signal \N__31559\ : std_logic;
signal \N__31554\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31541\ : std_logic;
signal \N__31540\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31537\ : std_logic;
signal \N__31536\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31534\ : std_logic;
signal \N__31533\ : std_logic;
signal \N__31532\ : std_logic;
signal \N__31531\ : std_logic;
signal \N__31530\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31528\ : std_logic;
signal \N__31527\ : std_logic;
signal \N__31526\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31524\ : std_logic;
signal \N__31523\ : std_logic;
signal \N__31522\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31520\ : std_logic;
signal \N__31519\ : std_logic;
signal \N__31516\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31514\ : std_logic;
signal \N__31513\ : std_logic;
signal \N__31512\ : std_logic;
signal \N__31511\ : std_logic;
signal \N__31510\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31508\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31492\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31476\ : std_logic;
signal \N__31467\ : std_logic;
signal \N__31458\ : std_logic;
signal \N__31455\ : std_logic;
signal \N__31446\ : std_logic;
signal \N__31437\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31427\ : std_logic;
signal \N__31424\ : std_logic;
signal \N__31421\ : std_logic;
signal \N__31418\ : std_logic;
signal \N__31411\ : std_logic;
signal \N__31406\ : std_logic;
signal \N__31403\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31390\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31386\ : std_logic;
signal \N__31381\ : std_logic;
signal \N__31380\ : std_logic;
signal \N__31379\ : std_logic;
signal \N__31376\ : std_logic;
signal \N__31373\ : std_logic;
signal \N__31368\ : std_logic;
signal \N__31365\ : std_logic;
signal \N__31362\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31351\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31344\ : std_logic;
signal \N__31341\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31331\ : std_logic;
signal \N__31328\ : std_logic;
signal \N__31327\ : std_logic;
signal \N__31326\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31317\ : std_logic;
signal \N__31312\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31304\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31298\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31294\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31290\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31284\ : std_logic;
signal \N__31281\ : std_logic;
signal \N__31280\ : std_logic;
signal \N__31277\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31269\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31259\ : std_logic;
signal \N__31256\ : std_logic;
signal \N__31255\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31244\ : std_logic;
signal \N__31243\ : std_logic;
signal \N__31242\ : std_logic;
signal \N__31241\ : std_logic;
signal \N__31238\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31226\ : std_logic;
signal \N__31223\ : std_logic;
signal \N__31220\ : std_logic;
signal \N__31217\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31211\ : std_logic;
signal \N__31208\ : std_logic;
signal \N__31205\ : std_logic;
signal \N__31202\ : std_logic;
signal \N__31199\ : std_logic;
signal \N__31196\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31192\ : std_logic;
signal \N__31189\ : std_logic;
signal \N__31186\ : std_logic;
signal \N__31181\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31175\ : std_logic;
signal \N__31174\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31170\ : std_logic;
signal \N__31165\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31159\ : std_logic;
signal \N__31156\ : std_logic;
signal \N__31153\ : std_logic;
signal \N__31150\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31144\ : std_logic;
signal \N__31139\ : std_logic;
signal \N__31136\ : std_logic;
signal \N__31135\ : std_logic;
signal \N__31132\ : std_logic;
signal \N__31129\ : std_logic;
signal \N__31124\ : std_logic;
signal \N__31121\ : std_logic;
signal \N__31120\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31104\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31088\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31070\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31064\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31058\ : std_logic;
signal \N__31055\ : std_logic;
signal \N__31052\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31040\ : std_logic;
signal \N__31037\ : std_logic;
signal \N__31034\ : std_logic;
signal \N__31031\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31025\ : std_logic;
signal \N__31022\ : std_logic;
signal \N__31019\ : std_logic;
signal \N__31016\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31010\ : std_logic;
signal \N__31007\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__30998\ : std_logic;
signal \N__30995\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30986\ : std_logic;
signal \N__30983\ : std_logic;
signal \N__30980\ : std_logic;
signal \N__30977\ : std_logic;
signal \N__30974\ : std_logic;
signal \N__30971\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30965\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30959\ : std_logic;
signal \N__30956\ : std_logic;
signal \N__30953\ : std_logic;
signal \N__30950\ : std_logic;
signal \N__30947\ : std_logic;
signal \N__30944\ : std_logic;
signal \N__30941\ : std_logic;
signal \N__30938\ : std_logic;
signal \N__30935\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30926\ : std_logic;
signal \N__30923\ : std_logic;
signal \N__30920\ : std_logic;
signal \N__30917\ : std_logic;
signal \N__30914\ : std_logic;
signal \N__30911\ : std_logic;
signal \N__30908\ : std_logic;
signal \N__30905\ : std_logic;
signal \N__30902\ : std_logic;
signal \N__30899\ : std_logic;
signal \N__30896\ : std_logic;
signal \N__30893\ : std_logic;
signal \N__30890\ : std_logic;
signal \N__30887\ : std_logic;
signal \N__30884\ : std_logic;
signal \N__30881\ : std_logic;
signal \N__30878\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30872\ : std_logic;
signal \N__30869\ : std_logic;
signal \N__30868\ : std_logic;
signal \N__30865\ : std_logic;
signal \N__30862\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30848\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30842\ : std_logic;
signal \N__30839\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30831\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30823\ : std_logic;
signal \N__30820\ : std_logic;
signal \N__30815\ : std_logic;
signal \N__30814\ : std_logic;
signal \N__30811\ : std_logic;
signal \N__30808\ : std_logic;
signal \N__30807\ : std_logic;
signal \N__30804\ : std_logic;
signal \N__30801\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30792\ : std_logic;
signal \N__30787\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30776\ : std_logic;
signal \N__30773\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30767\ : std_logic;
signal \N__30764\ : std_logic;
signal \N__30761\ : std_logic;
signal \N__30758\ : std_logic;
signal \N__30755\ : std_logic;
signal \N__30752\ : std_logic;
signal \N__30749\ : std_logic;
signal \N__30746\ : std_logic;
signal \N__30743\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30737\ : std_logic;
signal \N__30734\ : std_logic;
signal \N__30731\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30725\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30719\ : std_logic;
signal \N__30716\ : std_logic;
signal \N__30713\ : std_logic;
signal \N__30710\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30692\ : std_logic;
signal \N__30689\ : std_logic;
signal \N__30686\ : std_logic;
signal \N__30683\ : std_logic;
signal \N__30680\ : std_logic;
signal \N__30677\ : std_logic;
signal \N__30674\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30656\ : std_logic;
signal \N__30653\ : std_logic;
signal \N__30650\ : std_logic;
signal \N__30647\ : std_logic;
signal \N__30644\ : std_logic;
signal \N__30641\ : std_logic;
signal \N__30638\ : std_logic;
signal \N__30635\ : std_logic;
signal \N__30632\ : std_logic;
signal \N__30629\ : std_logic;
signal \N__30626\ : std_logic;
signal \N__30623\ : std_logic;
signal \N__30620\ : std_logic;
signal \N__30617\ : std_logic;
signal \N__30614\ : std_logic;
signal \N__30611\ : std_logic;
signal \N__30608\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30596\ : std_logic;
signal \N__30593\ : std_logic;
signal \N__30590\ : std_logic;
signal \N__30587\ : std_logic;
signal \N__30584\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30578\ : std_logic;
signal \N__30575\ : std_logic;
signal \N__30572\ : std_logic;
signal \N__30569\ : std_logic;
signal \N__30566\ : std_logic;
signal \N__30563\ : std_logic;
signal \N__30560\ : std_logic;
signal \N__30557\ : std_logic;
signal \N__30554\ : std_logic;
signal \N__30551\ : std_logic;
signal \N__30548\ : std_logic;
signal \N__30545\ : std_logic;
signal \N__30542\ : std_logic;
signal \N__30539\ : std_logic;
signal \N__30536\ : std_logic;
signal \N__30533\ : std_logic;
signal \N__30530\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30521\ : std_logic;
signal \N__30520\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30516\ : std_logic;
signal \N__30513\ : std_logic;
signal \N__30510\ : std_logic;
signal \N__30507\ : std_logic;
signal \N__30504\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30502\ : std_logic;
signal \N__30501\ : std_logic;
signal \N__30500\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30487\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30474\ : std_logic;
signal \N__30471\ : std_logic;
signal \N__30468\ : std_logic;
signal \N__30465\ : std_logic;
signal \N__30462\ : std_logic;
signal \N__30457\ : std_logic;
signal \N__30454\ : std_logic;
signal \N__30449\ : std_logic;
signal \N__30440\ : std_logic;
signal \N__30437\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30420\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30404\ : std_logic;
signal \N__30401\ : std_logic;
signal \N__30398\ : std_logic;
signal \N__30395\ : std_logic;
signal \N__30392\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30383\ : std_logic;
signal \N__30380\ : std_logic;
signal \N__30377\ : std_logic;
signal \N__30374\ : std_logic;
signal \N__30371\ : std_logic;
signal \N__30368\ : std_logic;
signal \N__30365\ : std_logic;
signal \N__30362\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30356\ : std_logic;
signal \N__30353\ : std_logic;
signal \N__30350\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30344\ : std_logic;
signal \N__30341\ : std_logic;
signal \N__30338\ : std_logic;
signal \N__30335\ : std_logic;
signal \N__30332\ : std_logic;
signal \N__30329\ : std_logic;
signal \N__30326\ : std_logic;
signal \N__30323\ : std_logic;
signal \N__30320\ : std_logic;
signal \N__30317\ : std_logic;
signal \N__30314\ : std_logic;
signal \N__30311\ : std_logic;
signal \N__30308\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30302\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30293\ : std_logic;
signal \N__30290\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30272\ : std_logic;
signal \N__30269\ : std_logic;
signal \N__30266\ : std_logic;
signal \N__30263\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30257\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30245\ : std_logic;
signal \N__30242\ : std_logic;
signal \N__30239\ : std_logic;
signal \N__30236\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30230\ : std_logic;
signal \N__30227\ : std_logic;
signal \N__30224\ : std_logic;
signal \N__30221\ : std_logic;
signal \N__30218\ : std_logic;
signal \N__30215\ : std_logic;
signal \N__30212\ : std_logic;
signal \N__30209\ : std_logic;
signal \N__30206\ : std_logic;
signal \N__30203\ : std_logic;
signal \N__30200\ : std_logic;
signal \N__30197\ : std_logic;
signal \N__30194\ : std_logic;
signal \N__30191\ : std_logic;
signal \N__30188\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30182\ : std_logic;
signal \N__30179\ : std_logic;
signal \N__30176\ : std_logic;
signal \N__30173\ : std_logic;
signal \N__30170\ : std_logic;
signal \N__30167\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30161\ : std_logic;
signal \N__30158\ : std_logic;
signal \N__30155\ : std_logic;
signal \N__30152\ : std_logic;
signal \N__30149\ : std_logic;
signal \N__30146\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30131\ : std_logic;
signal \N__30128\ : std_logic;
signal \N__30125\ : std_logic;
signal \N__30122\ : std_logic;
signal \N__30119\ : std_logic;
signal \N__30116\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30104\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30098\ : std_logic;
signal \N__30095\ : std_logic;
signal \N__30092\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30086\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30080\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30071\ : std_logic;
signal \N__30068\ : std_logic;
signal \N__30065\ : std_logic;
signal \N__30062\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30053\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30047\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30041\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30035\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30023\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30017\ : std_logic;
signal \N__30014\ : std_logic;
signal \N__30011\ : std_logic;
signal \N__30008\ : std_logic;
signal \N__30005\ : std_logic;
signal \N__30002\ : std_logic;
signal \N__29999\ : std_logic;
signal \N__29996\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29981\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29972\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29963\ : std_logic;
signal \N__29960\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29954\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29933\ : std_logic;
signal \N__29930\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29915\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29909\ : std_logic;
signal \N__29906\ : std_logic;
signal \N__29903\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29893\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29881\ : std_logic;
signal \N__29878\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29864\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29854\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29842\ : std_logic;
signal \N__29837\ : std_logic;
signal \N__29834\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29830\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29822\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29817\ : std_logic;
signal \N__29814\ : std_logic;
signal \N__29809\ : std_logic;
signal \N__29804\ : std_logic;
signal \N__29803\ : std_logic;
signal \N__29800\ : std_logic;
signal \N__29797\ : std_logic;
signal \N__29792\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29788\ : std_logic;
signal \N__29785\ : std_logic;
signal \N__29782\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29766\ : std_logic;
signal \N__29765\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29763\ : std_logic;
signal \N__29762\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29759\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29725\ : std_logic;
signal \N__29722\ : std_logic;
signal \N__29719\ : std_logic;
signal \N__29716\ : std_logic;
signal \N__29713\ : std_logic;
signal \N__29710\ : std_logic;
signal \N__29707\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29690\ : std_logic;
signal \N__29687\ : std_logic;
signal \N__29684\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29679\ : std_logic;
signal \N__29678\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29663\ : std_logic;
signal \N__29660\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29656\ : std_logic;
signal \N__29653\ : std_logic;
signal \N__29650\ : std_logic;
signal \N__29645\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29641\ : std_logic;
signal \N__29640\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29632\ : std_logic;
signal \N__29631\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29622\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29612\ : std_logic;
signal \N__29611\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29605\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29593\ : std_logic;
signal \N__29592\ : std_logic;
signal \N__29589\ : std_logic;
signal \N__29584\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29578\ : std_logic;
signal \N__29575\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29567\ : std_logic;
signal \N__29564\ : std_logic;
signal \N__29563\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29552\ : std_logic;
signal \N__29549\ : std_logic;
signal \N__29546\ : std_logic;
signal \N__29543\ : std_logic;
signal \N__29540\ : std_logic;
signal \N__29537\ : std_logic;
signal \N__29534\ : std_logic;
signal \N__29531\ : std_logic;
signal \N__29528\ : std_logic;
signal \N__29527\ : std_logic;
signal \N__29522\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29518\ : std_logic;
signal \N__29517\ : std_logic;
signal \N__29512\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29501\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29497\ : std_logic;
signal \N__29496\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29488\ : std_logic;
signal \N__29485\ : std_logic;
signal \N__29480\ : std_logic;
signal \N__29479\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29471\ : std_logic;
signal \N__29468\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29458\ : std_logic;
signal \N__29455\ : std_logic;
signal \N__29454\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29441\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29423\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29419\ : std_logic;
signal \N__29416\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29378\ : std_logic;
signal \N__29377\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29368\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29359\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29347\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29339\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29332\ : std_logic;
signal \N__29329\ : std_logic;
signal \N__29324\ : std_logic;
signal \N__29321\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29312\ : std_logic;
signal \N__29309\ : std_logic;
signal \N__29308\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29293\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29287\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29283\ : std_logic;
signal \N__29280\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29274\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29270\ : std_logic;
signal \N__29267\ : std_logic;
signal \N__29264\ : std_logic;
signal \N__29261\ : std_logic;
signal \N__29258\ : std_logic;
signal \N__29249\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29237\ : std_logic;
signal \N__29234\ : std_logic;
signal \N__29231\ : std_logic;
signal \N__29228\ : std_logic;
signal \N__29225\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29218\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29212\ : std_logic;
signal \N__29209\ : std_logic;
signal \N__29206\ : std_logic;
signal \N__29201\ : std_logic;
signal \N__29198\ : std_logic;
signal \N__29197\ : std_logic;
signal \N__29194\ : std_logic;
signal \N__29191\ : std_logic;
signal \N__29190\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29184\ : std_logic;
signal \N__29179\ : std_logic;
signal \N__29174\ : std_logic;
signal \N__29171\ : std_logic;
signal \N__29168\ : std_logic;
signal \N__29165\ : std_logic;
signal \N__29162\ : std_logic;
signal \N__29161\ : std_logic;
signal \N__29156\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29138\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29132\ : std_logic;
signal \N__29131\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29119\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29107\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29099\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29090\ : std_logic;
signal \N__29085\ : std_logic;
signal \N__29082\ : std_logic;
signal \N__29075\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29070\ : std_logic;
signal \N__29067\ : std_logic;
signal \N__29064\ : std_logic;
signal \N__29061\ : std_logic;
signal \N__29054\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29045\ : std_logic;
signal \N__29044\ : std_logic;
signal \N__29041\ : std_logic;
signal \N__29038\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29027\ : std_logic;
signal \N__29026\ : std_logic;
signal \N__29025\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29016\ : std_logic;
signal \N__29011\ : std_logic;
signal \N__29006\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__29001\ : std_logic;
signal \N__28998\ : std_logic;
signal \N__28995\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28986\ : std_logic;
signal \N__28983\ : std_logic;
signal \N__28980\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28970\ : std_logic;
signal \N__28967\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28953\ : std_logic;
signal \N__28946\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28932\ : std_logic;
signal \N__28929\ : std_logic;
signal \N__28928\ : std_logic;
signal \N__28925\ : std_logic;
signal \N__28922\ : std_logic;
signal \N__28919\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28907\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28903\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28886\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28877\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28871\ : std_logic;
signal \N__28868\ : std_logic;
signal \N__28865\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28849\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28840\ : std_logic;
signal \N__28837\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28827\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28818\ : std_logic;
signal \N__28815\ : std_logic;
signal \N__28812\ : std_logic;
signal \N__28809\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28799\ : std_logic;
signal \N__28796\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28782\ : std_logic;
signal \N__28777\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28770\ : std_logic;
signal \N__28767\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28754\ : std_logic;
signal \N__28751\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28747\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28741\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28739\ : std_logic;
signal \N__28736\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28728\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28720\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28710\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28700\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28698\ : std_logic;
signal \N__28695\ : std_logic;
signal \N__28692\ : std_logic;
signal \N__28689\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28681\ : std_logic;
signal \N__28680\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28670\ : std_logic;
signal \N__28667\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28659\ : std_logic;
signal \N__28656\ : std_logic;
signal \N__28653\ : std_logic;
signal \N__28650\ : std_logic;
signal \N__28647\ : std_logic;
signal \N__28640\ : std_logic;
signal \N__28639\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28635\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28629\ : std_logic;
signal \N__28622\ : std_logic;
signal \N__28619\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28617\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28596\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28587\ : std_logic;
signal \N__28580\ : std_logic;
signal \N__28577\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28571\ : std_logic;
signal \N__28568\ : std_logic;
signal \N__28565\ : std_logic;
signal \N__28562\ : std_logic;
signal \N__28559\ : std_logic;
signal \N__28556\ : std_logic;
signal \N__28553\ : std_logic;
signal \N__28552\ : std_logic;
signal \N__28549\ : std_logic;
signal \N__28546\ : std_logic;
signal \N__28541\ : std_logic;
signal \N__28538\ : std_logic;
signal \N__28535\ : std_logic;
signal \N__28532\ : std_logic;
signal \N__28529\ : std_logic;
signal \N__28526\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28514\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28508\ : std_logic;
signal \N__28505\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28499\ : std_logic;
signal \N__28496\ : std_logic;
signal \N__28493\ : std_logic;
signal \N__28490\ : std_logic;
signal \N__28487\ : std_logic;
signal \N__28484\ : std_logic;
signal \N__28481\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28475\ : std_logic;
signal \N__28472\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28468\ : std_logic;
signal \N__28467\ : std_logic;
signal \N__28466\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28464\ : std_logic;
signal \N__28457\ : std_logic;
signal \N__28454\ : std_logic;
signal \N__28453\ : std_logic;
signal \N__28452\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28445\ : std_logic;
signal \N__28442\ : std_logic;
signal \N__28439\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28427\ : std_logic;
signal \N__28422\ : std_logic;
signal \N__28419\ : std_logic;
signal \N__28416\ : std_logic;
signal \N__28413\ : std_logic;
signal \N__28410\ : std_logic;
signal \N__28403\ : std_logic;
signal \N__28400\ : std_logic;
signal \N__28397\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28390\ : std_logic;
signal \N__28387\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28379\ : std_logic;
signal \N__28376\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28370\ : std_logic;
signal \N__28367\ : std_logic;
signal \N__28364\ : std_logic;
signal \N__28361\ : std_logic;
signal \N__28358\ : std_logic;
signal \N__28357\ : std_logic;
signal \N__28354\ : std_logic;
signal \N__28351\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28345\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28334\ : std_logic;
signal \N__28331\ : std_logic;
signal \N__28328\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28318\ : std_logic;
signal \N__28315\ : std_logic;
signal \N__28312\ : std_logic;
signal \N__28309\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28298\ : std_logic;
signal \N__28295\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28289\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28283\ : std_logic;
signal \N__28280\ : std_logic;
signal \N__28277\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28273\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28267\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28256\ : std_logic;
signal \N__28255\ : std_logic;
signal \N__28252\ : std_logic;
signal \N__28249\ : std_logic;
signal \N__28244\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28238\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28232\ : std_logic;
signal \N__28229\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28225\ : std_logic;
signal \N__28222\ : std_logic;
signal \N__28219\ : std_logic;
signal \N__28214\ : std_logic;
signal \N__28211\ : std_logic;
signal \N__28208\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28202\ : std_logic;
signal \N__28201\ : std_logic;
signal \N__28198\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28192\ : std_logic;
signal \N__28189\ : std_logic;
signal \N__28186\ : std_logic;
signal \N__28181\ : std_logic;
signal \N__28178\ : std_logic;
signal \N__28175\ : std_logic;
signal \N__28172\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28165\ : std_logic;
signal \N__28162\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28156\ : std_logic;
signal \N__28153\ : std_logic;
signal \N__28150\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28142\ : std_logic;
signal \N__28141\ : std_logic;
signal \N__28138\ : std_logic;
signal \N__28135\ : std_logic;
signal \N__28132\ : std_logic;
signal \N__28129\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28115\ : std_logic;
signal \N__28112\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28096\ : std_logic;
signal \N__28093\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28085\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28075\ : std_logic;
signal \N__28072\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28061\ : std_logic;
signal \N__28058\ : std_logic;
signal \N__28055\ : std_logic;
signal \N__28052\ : std_logic;
signal \N__28049\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28042\ : std_logic;
signal \N__28039\ : std_logic;
signal \N__28036\ : std_logic;
signal \N__28033\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28025\ : std_logic;
signal \N__28024\ : std_logic;
signal \N__28021\ : std_logic;
signal \N__28018\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28012\ : std_logic;
signal \N__28009\ : std_logic;
signal \N__28006\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__27998\ : std_logic;
signal \N__27995\ : std_logic;
signal \N__27992\ : std_logic;
signal \N__27991\ : std_logic;
signal \N__27988\ : std_logic;
signal \N__27985\ : std_logic;
signal \N__27982\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27973\ : std_logic;
signal \N__27970\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27955\ : std_logic;
signal \N__27952\ : std_logic;
signal \N__27949\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27935\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27922\ : std_logic;
signal \N__27919\ : std_logic;
signal \N__27916\ : std_logic;
signal \N__27913\ : std_logic;
signal \N__27910\ : std_logic;
signal \N__27907\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27893\ : std_logic;
signal \N__27892\ : std_logic;
signal \N__27889\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27880\ : std_logic;
signal \N__27877\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27866\ : std_logic;
signal \N__27863\ : std_logic;
signal \N__27860\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27847\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27836\ : std_logic;
signal \N__27833\ : std_logic;
signal \N__27830\ : std_logic;
signal \N__27827\ : std_logic;
signal \N__27826\ : std_logic;
signal \N__27823\ : std_logic;
signal \N__27820\ : std_logic;
signal \N__27817\ : std_logic;
signal \N__27814\ : std_logic;
signal \N__27811\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27800\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27790\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27772\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27760\ : std_logic;
signal \N__27757\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27740\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27733\ : std_logic;
signal \N__27730\ : std_logic;
signal \N__27727\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27718\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27697\ : std_logic;
signal \N__27694\ : std_logic;
signal \N__27691\ : std_logic;
signal \N__27686\ : std_logic;
signal \N__27683\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27673\ : std_logic;
signal \N__27670\ : std_logic;
signal \N__27667\ : std_logic;
signal \N__27664\ : std_logic;
signal \N__27661\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27653\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27649\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27640\ : std_logic;
signal \N__27637\ : std_logic;
signal \N__27634\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27623\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27619\ : std_logic;
signal \N__27616\ : std_logic;
signal \N__27613\ : std_logic;
signal \N__27610\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27593\ : std_logic;
signal \N__27592\ : std_logic;
signal \N__27589\ : std_logic;
signal \N__27586\ : std_logic;
signal \N__27583\ : std_logic;
signal \N__27580\ : std_logic;
signal \N__27577\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27560\ : std_logic;
signal \N__27557\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27550\ : std_logic;
signal \N__27547\ : std_logic;
signal \N__27544\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27535\ : std_logic;
signal \N__27530\ : std_logic;
signal \N__27527\ : std_logic;
signal \N__27524\ : std_logic;
signal \N__27521\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27511\ : std_logic;
signal \N__27508\ : std_logic;
signal \N__27505\ : std_logic;
signal \N__27500\ : std_logic;
signal \N__27497\ : std_logic;
signal \N__27494\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27487\ : std_logic;
signal \N__27484\ : std_logic;
signal \N__27481\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27470\ : std_logic;
signal \N__27467\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27463\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27446\ : std_logic;
signal \N__27443\ : std_logic;
signal \N__27440\ : std_logic;
signal \N__27437\ : std_logic;
signal \N__27434\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27428\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27413\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27409\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27397\ : std_logic;
signal \N__27392\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27385\ : std_logic;
signal \N__27382\ : std_logic;
signal \N__27379\ : std_logic;
signal \N__27376\ : std_logic;
signal \N__27373\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27367\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27352\ : std_logic;
signal \N__27349\ : std_logic;
signal \N__27346\ : std_logic;
signal \N__27343\ : std_logic;
signal \N__27340\ : std_logic;
signal \N__27337\ : std_logic;
signal \N__27332\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27328\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27322\ : std_logic;
signal \N__27319\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27308\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27295\ : std_logic;
signal \N__27292\ : std_logic;
signal \N__27289\ : std_logic;
signal \N__27286\ : std_logic;
signal \N__27281\ : std_logic;
signal \N__27278\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27268\ : std_logic;
signal \N__27265\ : std_logic;
signal \N__27262\ : std_logic;
signal \N__27259\ : std_logic;
signal \N__27254\ : std_logic;
signal \N__27251\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27247\ : std_logic;
signal \N__27244\ : std_logic;
signal \N__27241\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27233\ : std_logic;
signal \N__27230\ : std_logic;
signal \N__27227\ : std_logic;
signal \N__27224\ : std_logic;
signal \N__27221\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27203\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27191\ : std_logic;
signal \N__27188\ : std_logic;
signal \N__27185\ : std_logic;
signal \N__27182\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27173\ : std_logic;
signal \N__27170\ : std_logic;
signal \N__27167\ : std_logic;
signal \N__27164\ : std_logic;
signal \N__27161\ : std_logic;
signal \N__27158\ : std_logic;
signal \N__27155\ : std_logic;
signal \N__27152\ : std_logic;
signal \N__27149\ : std_logic;
signal \N__27146\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27140\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27127\ : std_logic;
signal \N__27124\ : std_logic;
signal \N__27121\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27106\ : std_logic;
signal \N__27103\ : std_logic;
signal \N__27100\ : std_logic;
signal \N__27095\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27089\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27071\ : std_logic;
signal \N__27068\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27062\ : std_logic;
signal \N__27059\ : std_logic;
signal \N__27058\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27049\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27025\ : std_logic;
signal \N__27022\ : std_logic;
signal \N__27019\ : std_logic;
signal \N__27014\ : std_logic;
signal \N__27011\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26996\ : std_logic;
signal \N__26993\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26986\ : std_logic;
signal \N__26981\ : std_logic;
signal \N__26978\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26968\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26957\ : std_logic;
signal \N__26954\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26948\ : std_logic;
signal \N__26945\ : std_logic;
signal \N__26942\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26938\ : std_logic;
signal \N__26935\ : std_logic;
signal \N__26930\ : std_logic;
signal \N__26927\ : std_logic;
signal \N__26924\ : std_logic;
signal \N__26923\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26906\ : std_logic;
signal \N__26905\ : std_logic;
signal \N__26902\ : std_logic;
signal \N__26897\ : std_logic;
signal \N__26894\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26884\ : std_logic;
signal \N__26881\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26875\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26869\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26858\ : std_logic;
signal \N__26855\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26840\ : std_logic;
signal \N__26837\ : std_logic;
signal \N__26834\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26830\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26816\ : std_logic;
signal \N__26813\ : std_logic;
signal \N__26810\ : std_logic;
signal \N__26809\ : std_logic;
signal \N__26806\ : std_logic;
signal \N__26803\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26795\ : std_logic;
signal \N__26792\ : std_logic;
signal \N__26789\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26776\ : std_logic;
signal \N__26773\ : std_logic;
signal \N__26770\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26756\ : std_logic;
signal \N__26755\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26744\ : std_logic;
signal \N__26741\ : std_logic;
signal \N__26738\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26734\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26723\ : std_logic;
signal \N__26722\ : std_logic;
signal \N__26719\ : std_logic;
signal \N__26718\ : std_logic;
signal \N__26717\ : std_logic;
signal \N__26714\ : std_logic;
signal \N__26711\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26692\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26687\ : std_logic;
signal \N__26682\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26672\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26660\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26649\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26633\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26629\ : std_logic;
signal \N__26628\ : std_logic;
signal \N__26623\ : std_logic;
signal \N__26620\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26612\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26597\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26588\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26579\ : std_logic;
signal \N__26576\ : std_logic;
signal \N__26573\ : std_logic;
signal \N__26570\ : std_logic;
signal \N__26567\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26546\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26534\ : std_logic;
signal \N__26531\ : std_logic;
signal \N__26528\ : std_logic;
signal \N__26527\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26507\ : std_logic;
signal \N__26506\ : std_logic;
signal \N__26503\ : std_logic;
signal \N__26500\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26479\ : std_logic;
signal \N__26476\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26470\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26462\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26453\ : std_logic;
signal \N__26450\ : std_logic;
signal \N__26447\ : std_logic;
signal \N__26446\ : std_logic;
signal \N__26443\ : std_logic;
signal \N__26440\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26422\ : std_logic;
signal \N__26419\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26413\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26407\ : std_logic;
signal \N__26406\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26379\ : std_logic;
signal \N__26376\ : std_logic;
signal \N__26373\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26371\ : std_logic;
signal \N__26368\ : std_logic;
signal \N__26365\ : std_logic;
signal \N__26362\ : std_logic;
signal \N__26359\ : std_logic;
signal \N__26356\ : std_logic;
signal \N__26353\ : std_logic;
signal \N__26346\ : std_logic;
signal \N__26343\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26337\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26328\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26324\ : std_logic;
signal \N__26319\ : std_logic;
signal \N__26316\ : std_logic;
signal \N__26313\ : std_logic;
signal \N__26306\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26302\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26295\ : std_logic;
signal \N__26292\ : std_logic;
signal \N__26289\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26269\ : std_logic;
signal \N__26268\ : std_logic;
signal \N__26265\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26255\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26247\ : std_logic;
signal \N__26244\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26228\ : std_logic;
signal \N__26225\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26217\ : std_logic;
signal \N__26214\ : std_logic;
signal \N__26211\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26195\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26168\ : std_logic;
signal \N__26165\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26158\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26154\ : std_logic;
signal \N__26151\ : std_logic;
signal \N__26146\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26137\ : std_logic;
signal \N__26136\ : std_logic;
signal \N__26133\ : std_logic;
signal \N__26128\ : std_logic;
signal \N__26123\ : std_logic;
signal \N__26120\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26110\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26101\ : std_logic;
signal \N__26100\ : std_logic;
signal \N__26097\ : std_logic;
signal \N__26094\ : std_logic;
signal \N__26089\ : std_logic;
signal \N__26084\ : std_logic;
signal \N__26081\ : std_logic;
signal \N__26078\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26064\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25999\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25974\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25960\ : std_logic;
signal \N__25957\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25949\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25941\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25928\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25919\ : std_logic;
signal \N__25916\ : std_logic;
signal \N__25913\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25892\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25890\ : std_logic;
signal \N__25887\ : std_logic;
signal \N__25884\ : std_logic;
signal \N__25881\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25867\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25863\ : std_logic;
signal \N__25860\ : std_logic;
signal \N__25857\ : std_logic;
signal \N__25850\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25844\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25842\ : std_logic;
signal \N__25839\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25833\ : std_logic;
signal \N__25826\ : std_logic;
signal \N__25823\ : std_logic;
signal \N__25820\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25815\ : std_logic;
signal \N__25812\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25795\ : std_logic;
signal \N__25794\ : std_logic;
signal \N__25791\ : std_logic;
signal \N__25788\ : std_logic;
signal \N__25785\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25770\ : std_logic;
signal \N__25767\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25743\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25730\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25722\ : std_logic;
signal \N__25719\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25700\ : std_logic;
signal \N__25699\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25695\ : std_logic;
signal \N__25692\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25678\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25674\ : std_logic;
signal \N__25671\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25661\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25653\ : std_logic;
signal \N__25650\ : std_logic;
signal \N__25647\ : std_logic;
signal \N__25644\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25631\ : std_logic;
signal \N__25630\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25626\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25620\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25610\ : std_logic;
signal \N__25607\ : std_logic;
signal \N__25606\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25575\ : std_logic;
signal \N__25572\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25558\ : std_logic;
signal \N__25557\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25534\ : std_logic;
signal \N__25533\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25527\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25510\ : std_logic;
signal \N__25509\ : std_logic;
signal \N__25506\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25485\ : std_logic;
signal \N__25482\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25465\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25458\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25448\ : std_logic;
signal \N__25445\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25421\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25413\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25397\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25383\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25369\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25346\ : std_logic;
signal \N__25345\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25338\ : std_logic;
signal \N__25335\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25311\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25297\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25287\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25276\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25249\ : std_logic;
signal \N__25246\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25237\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25228\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25186\ : std_logic;
signal \N__25185\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25177\ : std_logic;
signal \N__25174\ : std_logic;
signal \N__25171\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25156\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25150\ : std_logic;
signal \N__25149\ : std_logic;
signal \N__25148\ : std_logic;
signal \N__25143\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25124\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25115\ : std_logic;
signal \N__25112\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25103\ : std_logic;
signal \N__25102\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25097\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25083\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25080\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25078\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25075\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25072\ : std_logic;
signal \N__25071\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25069\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25067\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25064\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25049\ : std_logic;
signal \N__25040\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25022\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25004\ : std_logic;
signal \N__24997\ : std_logic;
signal \N__24988\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24976\ : std_logic;
signal \N__24975\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24971\ : std_logic;
signal \N__24968\ : std_logic;
signal \N__24963\ : std_logic;
signal \N__24960\ : std_logic;
signal \N__24957\ : std_logic;
signal \N__24950\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24945\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24929\ : std_logic;
signal \N__24926\ : std_logic;
signal \N__24923\ : std_logic;
signal \N__24920\ : std_logic;
signal \N__24917\ : std_logic;
signal \N__24914\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24905\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24881\ : std_logic;
signal \N__24878\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24869\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24860\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24828\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24819\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24799\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24771\ : std_logic;
signal \N__24766\ : std_logic;
signal \N__24761\ : std_logic;
signal \N__24758\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24722\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24716\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24709\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24702\ : std_logic;
signal \N__24699\ : std_logic;
signal \N__24696\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24686\ : std_logic;
signal \N__24685\ : std_logic;
signal \N__24684\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24672\ : std_logic;
signal \N__24665\ : std_logic;
signal \N__24662\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24648\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24638\ : std_logic;
signal \N__24637\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24630\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24613\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24606\ : std_logic;
signal \N__24603\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24593\ : std_logic;
signal \N__24590\ : std_logic;
signal \N__24589\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24579\ : std_logic;
signal \N__24576\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24566\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24564\ : std_logic;
signal \N__24561\ : std_logic;
signal \N__24558\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24497\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24482\ : std_logic;
signal \N__24479\ : std_logic;
signal \N__24476\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24455\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24431\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24425\ : std_logic;
signal \N__24422\ : std_logic;
signal \N__24419\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24389\ : std_logic;
signal \N__24386\ : std_logic;
signal \N__24383\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24374\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24368\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24356\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24341\ : std_logic;
signal \N__24338\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24299\ : std_logic;
signal \N__24296\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24281\ : std_logic;
signal \N__24278\ : std_logic;
signal \N__24275\ : std_logic;
signal \N__24272\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24245\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24238\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24200\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24182\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24166\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24151\ : std_logic;
signal \N__24146\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24142\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24116\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24110\ : std_logic;
signal \N__24109\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24090\ : std_logic;
signal \N__24083\ : std_logic;
signal \N__24080\ : std_logic;
signal \N__24077\ : std_logic;
signal \N__24076\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24070\ : std_logic;
signal \N__24069\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24034\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24026\ : std_logic;
signal \N__24023\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23983\ : std_logic;
signal \N__23980\ : std_logic;
signal \N__23977\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23970\ : std_logic;
signal \N__23967\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23961\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23926\ : std_logic;
signal \N__23923\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23851\ : std_logic;
signal \N__23850\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23847\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23844\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23838\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23820\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23805\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23802\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23766\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23761\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23755\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23725\ : std_logic;
signal \N__23718\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23700\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23689\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23686\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23683\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23662\ : std_logic;
signal \N__23661\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23659\ : std_logic;
signal \N__23658\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23646\ : std_logic;
signal \N__23643\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23611\ : std_logic;
signal \N__23608\ : std_logic;
signal \N__23593\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23577\ : std_logic;
signal \N__23574\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23556\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23525\ : std_logic;
signal \N__23522\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23515\ : std_logic;
signal \N__23514\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23512\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23505\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23476\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23470\ : std_logic;
signal \N__23467\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23461\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23454\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23452\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23440\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23415\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23401\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23364\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23350\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23237\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23169\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23165\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23112\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23014\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23006\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22984\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22962\ : std_logic;
signal \N__22959\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22955\ : std_logic;
signal \N__22952\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22936\ : std_logic;
signal \N__22931\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22867\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22837\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22819\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22811\ : std_logic;
signal \N__22808\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22796\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22754\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22712\ : std_logic;
signal \N__22709\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22705\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22675\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22517\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22495\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22381\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22371\ : std_logic;
signal \N__22368\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22336\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22161\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22153\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22104\ : std_logic;
signal \N__22101\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22032\ : std_logic;
signal \N__22029\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22002\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21952\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21940\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21841\ : std_logic;
signal \N__21838\ : std_logic;
signal \N__21835\ : std_logic;
signal \N__21832\ : std_logic;
signal \N__21829\ : std_logic;
signal \N__21826\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21789\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21783\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21739\ : std_logic;
signal \N__21736\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21726\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21702\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21684\ : std_logic;
signal \N__21681\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21594\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21536\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21503\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21483\ : std_logic;
signal \N__21480\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21443\ : std_logic;
signal \N__21442\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21435\ : std_logic;
signal \N__21432\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21419\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21393\ : std_logic;
signal \N__21390\ : std_logic;
signal \N__21387\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21316\ : std_logic;
signal \N__21311\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21306\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21276\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21256\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21241\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21188\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21068\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21027\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21014\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20884\ : std_logic;
signal \N__20881\ : std_logic;
signal \N__20880\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20871\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20794\ : std_logic;
signal \N__20791\ : std_logic;
signal \N__20788\ : std_logic;
signal \N__20785\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20747\ : std_logic;
signal \N__20744\ : std_logic;
signal \N__20741\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20729\ : std_logic;
signal \N__20726\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20721\ : std_logic;
signal \N__20718\ : std_logic;
signal \N__20715\ : std_logic;
signal \N__20712\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20698\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20639\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20601\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20570\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20501\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20474\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20303\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20288\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20261\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20231\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19485\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19482\ : std_logic;
signal \N__19479\ : std_logic;
signal \N__19476\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19464\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19449\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19443\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19422\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19181\ : std_logic;
signal delay_tr_input_ibuf_gb_io_gb_input : std_logic;
signal delay_hc_input_ibuf_gb_io_gb_input : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_15\ : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_8\ : std_logic;
signal \bfn_1_12_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\ : std_logic;
signal \bfn_1_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_9\ : std_logic;
signal \bfn_1_14_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_17\ : std_logic;
signal \bfn_1_15_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_25\ : std_logic;
signal \bfn_1_16_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_98_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_96_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_97\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_96\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_94\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_91\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_161\ : std_logic;
signal \pwm_generator_inst.O_0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_0\ : std_logic;
signal \bfn_1_24_0_\ : std_logic;
signal \pwm_generator_inst.O_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_0\ : std_logic;
signal \pwm_generator_inst.O_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_1\ : std_logic;
signal \pwm_generator_inst.O_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_2\ : std_logic;
signal \pwm_generator_inst.O_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_3\ : std_logic;
signal \pwm_generator_inst.O_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_4\ : std_logic;
signal \pwm_generator_inst.O_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_5\ : std_logic;
signal \pwm_generator_inst.O_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_7\ : std_logic;
signal \pwm_generator_inst.O_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_8\ : std_logic;
signal \bfn_1_25_0_\ : std_logic;
signal \pwm_generator_inst.O_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_15\ : std_logic;
signal \bfn_1_26_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_2_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_43_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31\ : std_logic;
signal pwm_duty_input_0 : std_logic;
signal pwm_duty_input_1 : std_logic;
signal pwm_duty_input_2 : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_15\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_15_cascade_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_18\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_14\ : std_logic;
signal \rgb_drv_RNOZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_44_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_19_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_77\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_159\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\ : std_logic;
signal \bfn_3_23_0_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_7\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_7\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_8\ : std_logic;
signal \bfn_3_24_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433_cascade_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_3\ : std_logic;
signal \pwm_generator_inst.un1_duty_inputlt3\ : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0\ : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\ : std_logic;
signal pwm_duty_input_9 : std_logic;
signal pwm_duty_input_8 : std_logic;
signal pwm_duty_input_6 : std_logic;
signal pwm_duty_input_7 : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_12\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_1\ : std_logic;
signal \bfn_4_17_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\ : std_logic;
signal \bfn_4_18_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\ : std_logic;
signal \bfn_4_19_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\ : std_logic;
signal \bfn_4_20_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23\ : std_logic;
signal pwm_duty_input_3 : std_logic;
signal pwm_duty_input_4 : std_logic;
signal pwm_duty_input_5 : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\ : std_logic;
signal \pwm_generator_inst.N_17\ : std_logic;
signal \pwm_generator_inst.N_16\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033\ : std_logic;
signal \pwm_generator_inst.N_17_cascade_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\ : std_logic;
signal \pwm_generator_inst.O_10\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_0\ : std_logic;
signal clk_12mhz : std_logic;
signal \GB_BUFFER_clk_12mhz_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_46\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_47\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\ : std_logic;
signal \pwm_generator_inst.threshold_0\ : std_logic;
signal \pwm_generator_inst.counter_i_0\ : std_logic;
signal \bfn_5_23_0_\ : std_logic;
signal \pwm_generator_inst.un14_counter_1\ : std_logic;
signal \pwm_generator_inst.counter_i_1\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_0\ : std_logic;
signal \pwm_generator_inst.threshold_2\ : std_logic;
signal \pwm_generator_inst.counter_i_2\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_1\ : std_logic;
signal \pwm_generator_inst.threshold_3\ : std_logic;
signal \pwm_generator_inst.counter_i_3\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_2\ : std_logic;
signal \pwm_generator_inst.threshold_4\ : std_logic;
signal \pwm_generator_inst.counter_i_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_3\ : std_logic;
signal \pwm_generator_inst.threshold_5\ : std_logic;
signal \pwm_generator_inst.counter_i_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_6\ : std_logic;
signal \pwm_generator_inst.counter_i_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_7\ : std_logic;
signal \pwm_generator_inst.counter_i_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_8\ : std_logic;
signal \pwm_generator_inst.counter_i_8\ : std_logic;
signal \bfn_5_24_0_\ : std_logic;
signal \pwm_generator_inst.threshold_9\ : std_logic;
signal \pwm_generator_inst.counter_i_9\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_8\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_9\ : std_logic;
signal pwm_output_c : std_logic;
signal \N_38_i_i\ : std_logic;
signal \pwm_generator_inst.un1_counterlto9_2_cascade_\ : std_logic;
signal \pwm_generator_inst.un1_counterlto2_0_cascade_\ : std_logic;
signal \pwm_generator_inst.un1_counterlt9\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_0\ : std_logic;
signal \bfn_5_26_0_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_1\ : std_logic;
signal \pwm_generator_inst.counter_cry_0\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_3\ : std_logic;
signal \pwm_generator_inst.counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_5\ : std_logic;
signal \pwm_generator_inst.counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counter_cry_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_7\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_8\ : std_logic;
signal \bfn_5_27_0_\ : std_logic;
signal \pwm_generator_inst.un1_counter_0\ : std_logic;
signal \pwm_generator_inst.counter_cry_8\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_9\ : std_logic;
signal \bfn_7_7_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_7\ : std_logic;
signal \bfn_7_8_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_15\ : std_logic;
signal \bfn_7_9_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_23\ : std_logic;
signal \bfn_7_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.running_i\ : std_logic;
signal \phase_controller_inst2.start_timer_tr_RNO_0_0\ : std_logic;
signal \phase_controller_inst2.hc_time_passed\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_28\ : std_logic;
signal il_max_comp2_c : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_201_i\ : std_logic;
signal \phase_controller_inst2.state_RNI9M3OZ0Z_0\ : std_logic;
signal il_min_comp2_c : std_logic;
signal \phase_controller_inst2.stateZ0Z_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\ : std_logic;
signal \bfn_8_7_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\ : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\ : std_logic;
signal \bfn_8_9_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\ : std_logic;
signal \bfn_8_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\ : std_logic;
signal \bfn_8_11_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1Z0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \bfn_8_12_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_8_13_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\ : std_logic;
signal \bfn_8_14_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst2.tr_time_passed\ : std_logic;
signal \phase_controller_inst2.stoper_tr.runningZ0\ : std_logic;
signal \phase_controller_inst2.start_timer_hc_0_sqmuxa\ : std_logic;
signal \phase_controller_inst2.state_RNIG7JFZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_200_i\ : std_logic;
signal \delay_measurement_inst.start_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_trZ0\ : std_logic;
signal delay_tr_input_c_g : std_logic;
signal \phase_controller_inst2.stateZ0Z_3\ : std_logic;
signal s3_phy_c : std_logic;
signal \phase_controller_inst2.stateZ0Z_1\ : std_logic;
signal s4_phy_c : std_logic;
signal \GB_BUFFER_clock_output_0_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20\ : std_logic;
signal \elapsed_time_ns_1_RNIV9PBB_0_21_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI5FOBB_0_18_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \elapsed_time_ns_1_RNI1BOBB_0_14_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI1BOBB_0_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\ : std_logic;
signal \elapsed_time_ns_1_RNI5FOBB_0_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_9_12_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_9_13_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_16\ : std_logic;
signal \bfn_9_14_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axb_0\ : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_8\ : std_logic;
signal \bfn_9_16_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_16\ : std_logic;
signal \bfn_9_17_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_24\ : std_logic;
signal \bfn_9_18_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.un8_enablelto31\ : std_logic;
signal \pwm_generator_inst.un3_threshold\ : std_logic;
signal \bfn_9_26_0_\ : std_logic;
signal \pwm_generator_inst.O_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_0\ : std_logic;
signal \pwm_generator_inst.O_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_1\ : std_logic;
signal \pwm_generator_inst.O_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_2\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_3\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_4\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_5\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_6\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_7\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11\ : std_logic;
signal \bfn_9_27_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_9\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_15\ : std_logic;
signal \bfn_9_28_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_16\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_17\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19\ : std_logic;
signal il_min_comp1_c : std_logic;
signal \il_min_comp1_D1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\ : std_logic;
signal \elapsed_time_ns_1_RNIHG91B_0_5\ : std_logic;
signal \elapsed_time_ns_1_RNIV8OBB_0_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\ : std_logic;
signal \elapsed_time_ns_1_RNI0BPBB_0_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\ : std_logic;
signal \elapsed_time_ns_1_RNI1CPBB_0_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\ : std_logic;
signal \elapsed_time_ns_1_RNI7IPBB_0_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\ : std_logic;
signal \elapsed_time_ns_1_RNIU7OBB_0_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\ : std_logic;
signal \elapsed_time_ns_1_RNIU7OBB_0_11_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIT6OBB_0_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\ : std_logic;
signal \elapsed_time_ns_1_RNIT6OBB_0_10_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNILK91B_0_9_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIU8PBB_0_20_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI2COBB_0_15_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\ : std_logic;
signal \elapsed_time_ns_1_RNI6HPBB_0_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_29\ : std_logic;
signal \elapsed_time_ns_1_RNIVAQBB_0_30\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\ : std_logic;
signal \elapsed_time_ns_1_RNI6GOBB_0_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \elapsed_time_ns_1_RNIFE91B_0_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\ : std_logic;
signal \elapsed_time_ns_1_RNIV9PBB_0_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\ : std_logic;
signal \elapsed_time_ns_1_RNIU8PBB_0_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\ : std_logic;
signal \elapsed_time_ns_1_RNILK91B_0_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\ : std_logic;
signal \elapsed_time_ns_1_RNIIH91B_0_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\ : std_logic;
signal \elapsed_time_ns_1_RNI2COBB_0_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_start_g\ : std_logic;
signal \current_shift_inst.control_input_axb_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_axbZ0Z_4\ : std_logic;
signal \bfn_10_26_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_18\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_20\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_21\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_22\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_23\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0\ : std_logic;
signal \bfn_10_27_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_24\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_9\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\ : std_logic;
signal \bfn_10_28_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_23\ : std_logic;
signal \elapsed_time_ns_1_RNIGF91B_0_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_11_8_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\ : std_logic;
signal \bfn_11_10_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26\ : std_logic;
signal \elapsed_time_ns_1_RNI5GPBB_0_27\ : std_logic;
signal \elapsed_time_ns_1_RNI5GPBB_0_27_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\ : std_logic;
signal \elapsed_time_ns_1_RNI4FPBB_0_26\ : std_logic;
signal \elapsed_time_ns_1_RNI4FPBB_0_26_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latchedZ0\ : std_logic;
signal \phase_controller_inst2.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un2_start_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un2_start_0_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.runningZ0\ : std_logic;
signal \phase_controller_inst2.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latchedZ0\ : std_logic;
signal \T45_c\ : std_logic;
signal \current_shift_inst.control_input_axb_0\ : std_logic;
signal \current_shift_inst.N_1269_i\ : std_logic;
signal \current_shift_inst.control_input_1\ : std_logic;
signal \bfn_11_15_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\ : std_logic;
signal \current_shift_inst.control_input_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\ : std_logic;
signal \current_shift_inst.control_input_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\ : std_logic;
signal \current_shift_inst.control_input_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\ : std_logic;
signal \current_shift_inst.control_input_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\ : std_logic;
signal \current_shift_inst.control_input_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\ : std_logic;
signal \current_shift_inst.control_input_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\ : std_logic;
signal \current_shift_inst.control_input_cry_6\ : std_logic;
signal \current_shift_inst.control_input_cry_7\ : std_logic;
signal \current_shift_inst.control_input_axb_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\ : std_logic;
signal \bfn_11_16_0_\ : std_logic;
signal \current_shift_inst.control_input_axb_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\ : std_logic;
signal \current_shift_inst.control_input_cry_8\ : std_logic;
signal \current_shift_inst.control_input_axb_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\ : std_logic;
signal \current_shift_inst.control_input_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\ : std_logic;
signal \current_shift_inst.control_input_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\ : std_logic;
signal \current_shift_inst.control_input_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\ : std_logic;
signal \current_shift_inst.control_input_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14\ : std_logic;
signal \current_shift_inst.control_input_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15\ : std_logic;
signal \current_shift_inst.control_input_cry_14\ : std_logic;
signal \current_shift_inst.control_input_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16\ : std_logic;
signal \bfn_11_17_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17\ : std_logic;
signal \current_shift_inst.control_input_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18\ : std_logic;
signal \current_shift_inst.control_input_cry_17\ : std_logic;
signal \current_shift_inst.control_input_axb_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19\ : std_logic;
signal \current_shift_inst.control_input_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20\ : std_logic;
signal \current_shift_inst.control_input_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21\ : std_logic;
signal \current_shift_inst.control_input_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22\ : std_logic;
signal \current_shift_inst.control_input_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23\ : std_logic;
signal \current_shift_inst.control_input_cry_22\ : std_logic;
signal \current_shift_inst.control_input_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24\ : std_logic;
signal \bfn_11_18_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25\ : std_logic;
signal \current_shift_inst.control_input_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26\ : std_logic;
signal \current_shift_inst.control_input_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27\ : std_logic;
signal \current_shift_inst.control_input_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28\ : std_logic;
signal \current_shift_inst.control_input_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29\ : std_logic;
signal \current_shift_inst.control_input_cry_28\ : std_logic;
signal \current_shift_inst.control_input_cry_29\ : std_logic;
signal \current_shift_inst.control_input_31\ : std_logic;
signal \current_shift_inst.control_input_axb_27\ : std_logic;
signal \current_shift_inst.control_input_axb_18\ : std_logic;
signal \current_shift_inst.control_input_axb_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_25\ : std_logic;
signal \N_19_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\ : std_logic;
signal il_max_comp1_c : std_logic;
signal \il_max_comp1_D1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\ : std_logic;
signal \elapsed_time_ns_1_RNI0CQBB_0_31\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\ : std_logic;
signal \elapsed_time_ns_1_RNIDC91B_0_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\ : std_logic;
signal \bfn_12_7_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_12_8_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_12_9_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\ : std_logic;
signal \bfn_12_10_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\ : std_logic;
signal \elapsed_time_ns_1_RNI0AOBB_0_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\ : std_logic;
signal \elapsed_time_ns_1_RNI0AOBB_0_13_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \elapsed_time_ns_1_RNI4EOBB_0_17\ : std_logic;
signal \elapsed_time_ns_1_RNI4EOBB_0_17_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt16\ : std_logic;
signal \elapsed_time_ns_1_RNI3DOBB_0_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\ : std_logic;
signal \elapsed_time_ns_1_RNI3DOBB_0_16_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1Z0Z_30\ : std_logic;
signal \phase_controller_inst1.tr_time_passed\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.state_RNI7NN7Z0Z_0_cascade_\ : std_logic;
signal state_ns_i_a3_1 : std_logic;
signal start_stop_c : std_logic;
signal \current_shift_inst.control_input_axb_1\ : std_logic;
signal \current_shift_inst.control_input_axb_2\ : std_logic;
signal \current_shift_inst.control_input_axb_3\ : std_logic;
signal \current_shift_inst.control_input_axb_4\ : std_logic;
signal \current_shift_inst.control_input_axb_5\ : std_logic;
signal \current_shift_inst.control_input_axb_6\ : std_logic;
signal \bfn_12_16_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_3\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_4\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_5\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_6\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_7\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_8\ : std_logic;
signal \bfn_12_17_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_9\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_11\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_12\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_13\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s0\ : std_logic;
signal \bfn_12_18_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s0\ : std_logic;
signal \bfn_12_19_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s0\ : std_logic;
signal \current_shift_inst.control_input_axb_28\ : std_logic;
signal \current_shift_inst.control_input_axb_29\ : std_logic;
signal \pll_inst.red_c_i\ : std_logic;
signal delay_hc_input_c_g : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\ : std_logic;
signal \elapsed_time_ns_1_RNIED91B_0_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24\ : std_logic;
signal \elapsed_time_ns_1_RNI3EPBB_0_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_25\ : std_logic;
signal \elapsed_time_ns_1_RNI2DPBB_0_24\ : std_logic;
signal \elapsed_time_ns_1_RNI2DPBB_0_24_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_24\ : std_logic;
signal \elapsed_time_ns_1_RNIJI91B_0_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3\ : std_logic;
signal \elapsed_time_ns_1_RNIKJ91B_0_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_start_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.runningZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un2_start_0\ : std_logic;
signal \phase_controller_inst1.state_RNI7NN7Z0Z_0\ : std_logic;
signal \phase_controller_inst1.start_timer_tr_RNOZ0Z_0\ : std_logic;
signal \phase_controller_inst1.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latchedZ0\ : std_logic;
signal \il_min_comp1_D2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_30\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_10\ : std_logic;
signal \current_shift_inst.control_input_axb_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_14\ : std_logic;
signal \current_shift_inst.control_input_axb_11\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_15\ : std_logic;
signal \current_shift_inst.control_input_axb_12\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_16\ : std_logic;
signal \current_shift_inst.control_input_axb_13\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_17\ : std_logic;
signal \current_shift_inst.control_input_axb_14\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_18\ : std_logic;
signal \current_shift_inst.control_input_axb_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_19\ : std_logic;
signal \current_shift_inst.control_input_axb_16\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_28\ : std_logic;
signal \current_shift_inst.control_input_axb_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_27\ : std_logic;
signal \current_shift_inst.control_input_axb_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_29\ : std_logic;
signal \current_shift_inst.control_input_axb_26\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_23\ : std_logic;
signal \current_shift_inst.control_input_axb_20\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_24\ : std_logic;
signal \current_shift_inst.control_input_axb_21\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_25\ : std_logic;
signal \current_shift_inst.control_input_axb_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_26\ : std_logic;
signal \current_shift_inst.control_input_axb_23\ : std_logic;
signal \il_max_comp1_D2\ : std_logic;
signal \T01_c\ : std_logic;
signal state_3 : std_logic;
signal s1_phy_c : std_logic;
signal \current_shift_inst.timer_s1.N_162_i\ : std_logic;
signal s2_phy_c : std_logic;
signal \delay_measurement_inst.start_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_hcZ0\ : std_logic;
signal \elapsed_time_ns_1_RNIV2EN9_0_30\ : std_logic;
signal \elapsed_time_ns_1_RNI02CN9_0_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\ : std_logic;
signal \bfn_14_11_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1Z0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \bfn_14_12_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_14_13_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\ : std_logic;
signal \bfn_14_14_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\ : std_logic;
signal \bfn_14_15_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_3\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_4\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_5\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_6\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_7\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_8\ : std_logic;
signal \bfn_14_16_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_9\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_10\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_11\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_12\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_13\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_14\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_15\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_16\ : std_logic;
signal \bfn_14_17_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_17\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_18\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_19\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_24\ : std_logic;
signal \bfn_14_18_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_25\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI00M61_4\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\ : std_logic;
signal \current_shift_inst.start_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.stop_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\ : std_logic;
signal \elapsed_time_ns_1_RNI04EN9_0_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3\ : std_logic;
signal \elapsed_time_ns_1_RNITUBN9_0_10\ : std_logic;
signal \elapsed_time_ns_1_RNITUBN9_0_10_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIUVBN9_0_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_20\ : std_logic;
signal \elapsed_time_ns_1_RNIL73T9_0_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \elapsed_time_ns_1_RNII43T9_0_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_15_13_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_15_14_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\ : std_logic;
signal \bfn_15_15_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI25021_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\ : std_logic;
signal \current_shift_inst.timer_s1.runningZ0\ : std_logic;
signal \bfn_16_5_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_7\ : std_logic;
signal \bfn_16_6_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_15\ : std_logic;
signal \bfn_16_7_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_23\ : std_logic;
signal \bfn_16_8_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_199_i\ : std_logic;
signal \bfn_16_9_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\ : std_logic;
signal \bfn_16_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\ : std_logic;
signal \bfn_16_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\ : std_logic;
signal \bfn_16_12_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI68O61_6\ : std_logic;
signal \bfn_16_15_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_8\ : std_logic;
signal \bfn_16_16_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_16\ : std_logic;
signal \bfn_16_17_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_17\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_25\ : std_logic;
signal \bfn_16_18_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_26\ : std_logic;
signal \current_shift_inst.un4_control_input1_29\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_31\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_24\ : std_logic;
signal \bfn_16_19_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \bfn_16_20_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \bfn_16_21_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \bfn_16_22_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_29\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_28\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_23\ : std_logic;
signal \current_shift_inst.un4_control_input1_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_25\ : std_logic;
signal \current_shift_inst.un4_control_input1_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISST11_17\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_1\ : std_logic;
signal \T23_c\ : std_logic;
signal \elapsed_time_ns_1_RNIV1DN9_0_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\ : std_logic;
signal \elapsed_time_ns_1_RNIK63T9_0_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\ : std_logic;
signal \elapsed_time_ns_1_RNIV0CN9_0_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\ : std_logic;
signal \elapsed_time_ns_1_RNIH33T9_0_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_17_10_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_17_11_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_16\ : std_logic;
signal \bfn_17_12_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24\ : std_logic;
signal \elapsed_time_ns_1_RNI36DN9_0_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\ : std_logic;
signal \elapsed_time_ns_1_RNI36DN9_0_25_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\ : std_logic;
signal \elapsed_time_ns_1_RNI25DN9_0_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_1\ : std_logic;
signal \current_shift_inst.un38_control_input_5_1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_2\ : std_logic;
signal \current_shift_inst.un4_control_input1_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\ : std_logic;
signal \current_shift_inst.un38_control_input_axb_31_s0\ : std_logic;
signal \current_shift_inst.un4_control_input1_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\ : std_logic;
signal \current_shift_inst.un38_control_input_5_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_6\ : std_logic;
signal \current_shift_inst.un4_control_input1_6\ : std_logic;
signal \current_shift_inst.un4_control_input1_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_7\ : std_logic;
signal \current_shift_inst.un4_control_input1_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_11\ : std_logic;
signal \current_shift_inst.un4_control_input1_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_9\ : std_logic;
signal \current_shift_inst.un4_control_input1_9\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0_sf\ : std_logic;
signal \current_shift_inst.un4_control_input1_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_5\ : std_logic;
signal \current_shift_inst.un4_control_input1_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI34N61_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_16\ : std_logic;
signal \current_shift_inst.un4_control_input1_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_13\ : std_logic;
signal \current_shift_inst.un4_control_input1_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_17\ : std_logic;
signal \current_shift_inst.un4_control_input1_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_15\ : std_logic;
signal \current_shift_inst.un4_control_input1_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_20\ : std_logic;
signal \current_shift_inst.un4_control_input1_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_19\ : std_logic;
signal \current_shift_inst.un4_control_input1_19\ : std_logic;
signal \current_shift_inst.un4_control_input1_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_22\ : std_logic;
signal \current_shift_inst.un4_control_input1_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_24\ : std_logic;
signal \current_shift_inst.un4_control_input1_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_8\ : std_logic;
signal \current_shift_inst.un4_control_input1_8\ : std_logic;
signal \current_shift_inst.un4_control_input1_31_THRU_CO\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_9\ : std_logic;
signal \current_shift_inst.un38_control_input_5_2\ : std_logic;
signal \current_shift_inst.un4_control_input1_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_30\ : std_logic;
signal \current_shift_inst.un4_control_input1_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_3\ : std_logic;
signal \current_shift_inst.un4_control_input1_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_4\ : std_logic;
signal \current_shift_inst.un4_control_input1_4\ : std_logic;
signal \bfn_17_20_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\ : std_logic;
signal \bfn_17_21_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\ : std_logic;
signal \bfn_17_22_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\ : std_logic;
signal \bfn_17_23_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\ : std_logic;
signal \elapsed_time_ns_1_RNIU0DN9_0_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_198_i\ : std_logic;
signal \elapsed_time_ns_1_RNIE03T9_0_2\ : std_logic;
signal \elapsed_time_ns_1_RNIF13T9_0_3\ : std_logic;
signal \elapsed_time_ns_1_RNIG23T9_0_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\ : std_logic;
signal \elapsed_time_ns_1_RNI68CN9_0_19\ : std_logic;
signal \elapsed_time_ns_1_RNI68CN9_0_19_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \elapsed_time_ns_1_RNI24CN9_0_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_18_11_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1Z0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_18_12_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_18_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\ : std_logic;
signal \bfn_18_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31\ : std_logic;
signal \current_shift_inst.un4_control_input1_1_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_fast_31\ : std_logic;
signal \current_shift_inst.timer_s1.N_162_i_g\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31_rep1\ : std_logic;
signal \current_shift_inst.un4_control_input1_12\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_11\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_0\ : std_logic;
signal \bfn_18_17_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_1\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_0\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_2\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_1\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_3\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_4\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_5\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_7\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_8\ : std_logic;
signal \bfn_18_18_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_10\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_11\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_12\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_13\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_15\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_16\ : std_logic;
signal \bfn_18_19_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_17\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_18\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_19\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_20\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_21\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_23\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_24\ : std_logic;
signal \bfn_18_20_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_25\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_26\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_27\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_28\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.running_i\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_29\ : std_logic;
signal \current_shift_inst.timer_s1.N_163_i\ : std_logic;
signal \T12_c\ : std_logic;
signal \elapsed_time_ns_1_RNIDV2T9_0_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.runningZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_start_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\ : std_logic;
signal phase_controller_inst1_state_4 : std_logic;
signal \phase_controller_inst1.start_timer_hc_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latchedZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt16\ : std_logic;
signal \elapsed_time_ns_1_RNI46CN9_0_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\ : std_logic;
signal \elapsed_time_ns_1_RNI46CN9_0_17_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\ : std_logic;
signal \elapsed_time_ns_1_RNI13CN9_0_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\ : std_logic;
signal \elapsed_time_ns_1_RNI13CN9_0_14_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_29\ : std_logic;
signal \elapsed_time_ns_1_RNIJ53T9_0_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\ : std_logic;
signal \elapsed_time_ns_1_RNIJ53T9_0_7_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \elapsed_time_ns_1_RNI7ADN9_0_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt28\ : std_logic;
signal \elapsed_time_ns_1_RNI69DN9_0_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\ : std_logic;
signal \elapsed_time_ns_1_RNI69DN9_0_28_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst1.hc_time_passed\ : std_logic;
signal \phase_controller_inst1.state_RNIE87FZ0Z_2\ : std_logic;
signal \elapsed_time_ns_1_RNI57CN9_0_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_start_g\ : std_logic;
signal \elapsed_time_ns_1_RNI35CN9_0_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \elapsed_time_ns_1_RNI03DN9_0_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt22\ : std_logic;
signal \elapsed_time_ns_1_RNI14DN9_0_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\ : std_logic;
signal \elapsed_time_ns_1_RNI14DN9_0_23_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22\ : std_logic;
signal \elapsed_time_ns_1_RNI47DN9_0_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\ : std_logic;
signal clock_output_0 : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\ : std_logic;
signal red_c_g : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3\ : std_logic;
signal \elapsed_time_ns_1_RNI58DN9_0_27\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal reset_wire : std_logic;
signal clock_output_wire : std_logic;
signal \T01_wire\ : std_logic;
signal start_stop_wire : std_logic;
signal il_max_comp2_wire : std_logic;
signal \T23_wire\ : std_logic;
signal pwm_output_wire : std_logic;
signal il_max_comp1_wire : std_logic;
signal s2_phy_wire : std_logic;
signal \T12_wire\ : std_logic;
signal il_min_comp2_wire : std_logic;
signal s1_phy_wire : std_logic;
signal s4_phy_wire : std_logic;
signal il_min_comp1_wire : std_logic;
signal s3_phy_wire : std_logic;
signal \T45_wire\ : std_logic;
signal delay_hc_input_wire : std_logic;
signal delay_tr_input_wire : std_logic;
signal rgb_b_wire : std_logic;
signal rgb_g_wire : std_logic;
signal rgb_r_wire : std_logic;
signal \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\ : std_logic_vector(31 downto 0);

begin
    reset_wire <= reset;
    clock_output <= clock_output_wire;
    T01 <= \T01_wire\;
    start_stop_wire <= start_stop;
    il_max_comp2_wire <= il_max_comp2;
    T23 <= \T23_wire\;
    pwm_output <= pwm_output_wire;
    il_max_comp1_wire <= il_max_comp1;
    s2_phy <= s2_phy_wire;
    T12 <= \T12_wire\;
    il_min_comp2_wire <= il_min_comp2;
    s1_phy <= s1_phy_wire;
    s4_phy <= s4_phy_wire;
    il_min_comp1_wire <= il_min_comp1;
    s3_phy <= s3_phy_wire;
    T45 <= \T45_wire\;
    delay_hc_input_wire <= delay_hc_input;
    delay_tr_input_wire <= delay_tr_input;
    rgb_b <= rgb_b_wire;
    rgb_g <= rgb_g_wire;
    rgb_r <= rgb_r_wire;
    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\ <= \N__27998\&\N__28024\&\N__28055\&\N__28082\&\N__28115\&\N__28141\&\N__28175\&\N__28208\&\N__27737\&\N__27763\&\N__27800\&\N__27833\&\N__27859\&\N__27899\&\N__27929\&\N__27962\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__48410\&'0'&\N__48409\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(15);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_14\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(14);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_13\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(13);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_12\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(12);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_11\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(11);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_10\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(10);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_9\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(9);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_8\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(8);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_7\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(7);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_6\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(6);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_5\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(5);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_4\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(4);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_3\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(3);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_2\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(2);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_1\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(1);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_0\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\ <= '0'&\N__32470\&\N__32463\&\N__32468\&\N__32462\&\N__32469\&\N__32461\&\N__32471\&\N__32458\&\N__32464\&\N__32457\&\N__32465\&\N__32459\&\N__32466\&\N__32460\&\N__32467\;
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__48305\&\N__48302\&'0'&'0'&'0'&\N__48300\&\N__48304\&\N__48301\&\N__48303\;
    \pwm_generator_inst.un2_threshold_2_1_16\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_2_1_15\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.un2_threshold_2_14\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.un2_threshold_2_13\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.un2_threshold_2_12\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un2_threshold_2_11\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.un2_threshold_2_10\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.un2_threshold_2_9\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.un2_threshold_2_8\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.un2_threshold_2_7\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.un2_threshold_2_6\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.un2_threshold_2_5\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.un2_threshold_2_4\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.un2_threshold_2_3\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.un2_threshold_2_2\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.un2_threshold_2_1\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.un2_threshold_2_0\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\ <= '0'&\N__32406\&\N__32409\&\N__32407\&\N__32410\&\N__32408\&\N__21328\&\N__21306\&\N__21250\&\N__21276\&\N__24108\&\N__24135\&\N__24165\&\N__20555\&\N__20573\&\N__20588\;
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__48418\&\N__48415\&'0'&'0'&'0'&\N__48413\&\N__48417\&\N__48414\&\N__48416\;
    \pwm_generator_inst.un2_threshold_1_25\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(25);
    \pwm_generator_inst.un2_threshold_1_24\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(24);
    \pwm_generator_inst.un2_threshold_1_23\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(23);
    \pwm_generator_inst.un2_threshold_1_22\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(22);
    \pwm_generator_inst.un2_threshold_1_21\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(21);
    \pwm_generator_inst.un2_threshold_1_20\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(20);
    \pwm_generator_inst.un2_threshold_1_19\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(19);
    \pwm_generator_inst.un2_threshold_1_18\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(18);
    \pwm_generator_inst.un2_threshold_1_17\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(17);
    \pwm_generator_inst.un2_threshold_1_16\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_1_15\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.O_14\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.O_13\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.O_12\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un3_threshold\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.O_10\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.O_9\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.O_8\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.O_7\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.O_6\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.O_5\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.O_4\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.O_3\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.O_2\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.O_1\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.O_0\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(0);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\ <= '0'&\N__27470\&\N__27493\&\N__27527\&\N__27557\&\N__27593\&\N__27626\&\N__27650\&\N__27680\&\N__27704\&\N__27271\&\N__27299\&\N__27329\&\N__27359\&\N__27385\&\N__29726\;
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__48407\&'0'&\N__48406\;
    \current_shift_inst.PI_CTRL.integrator_1_0_1_19\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(19);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_18\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(18);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_17\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(17);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_16\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(16);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(15);
    \current_shift_inst.PI_CTRL.integrator_1_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(14);
    \current_shift_inst.PI_CTRL.integrator_1_14\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(13);
    \current_shift_inst.PI_CTRL.integrator_1_13\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(12);
    \current_shift_inst.PI_CTRL.integrator_1_12\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(11);
    \current_shift_inst.PI_CTRL.integrator_1_11\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(10);
    \current_shift_inst.PI_CTRL.integrator_1_10\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(9);
    \current_shift_inst.PI_CTRL.integrator_1_9\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(8);
    \current_shift_inst.PI_CTRL.integrator_1_8\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(7);
    \current_shift_inst.PI_CTRL.integrator_1_7\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(6);
    \current_shift_inst.PI_CTRL.integrator_1_6\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(5);
    \current_shift_inst.PI_CTRL.integrator_1_5\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(4);
    \current_shift_inst.PI_CTRL.integrator_1_4\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(3);
    \current_shift_inst.PI_CTRL.integrator_1_3\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(2);
    \current_shift_inst.PI_CTRL.integrator_1_2\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(1);
    \current_shift_inst.PI_CTRL.un1_integrator\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(0);

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__23894\,
            RESETB => \N__34067\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => clock_output_0
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__48411\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__48408\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\,
            ADDSUBBOT => '0',
            A => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\,
            C => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\,
            B => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\,
            OHOLDTOP => '0',
            O => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__48348\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__48299\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__48436\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__48412\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__48371\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__48405\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\,
            ADDSUBBOT => '0',
            A => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\,
            C => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\,
            B => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\,
            OHOLDTOP => '0',
            O => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\
        );

    \reset_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__50562\,
            GLOBALBUFFEROUTPUT => red_c_g
        );

    \reset_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50564\,
            DIN => \N__50563\,
            DOUT => \N__50562\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50564\,
            PADOUT => \N__50563\,
            PADIN => \N__50562\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clock_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50553\,
            DIN => \N__50552\,
            DOUT => \N__50551\,
            PACKAGEPIN => clock_output_wire
        );

    \clock_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50553\,
            PADOUT => \N__50552\,
            PADIN => \N__50551\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__26171\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T01_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50544\,
            DIN => \N__50543\,
            DOUT => \N__50542\,
            PACKAGEPIN => \T01_wire\
        );

    \T01_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50544\,
            PADOUT => \N__50543\,
            PADIN => \N__50542\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__35654\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \start_stop_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50535\,
            DIN => \N__50534\,
            DOUT => \N__50533\,
            PACKAGEPIN => start_stop_wire
        );

    \start_stop_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50535\,
            PADOUT => \N__50534\,
            PADIN => \N__50533\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => start_stop_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50526\,
            DIN => \N__50525\,
            DOUT => \N__50524\,
            PACKAGEPIN => il_max_comp2_wire
        );

    \il_max_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50526\,
            PADOUT => \N__50525\,
            PADIN => \N__50524\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T23_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50517\,
            DIN => \N__50516\,
            DOUT => \N__50515\,
            PACKAGEPIN => \T23_wire\
        );

    \T23_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50517\,
            PADOUT => \N__50516\,
            PADIN => \N__50515\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__39818\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50508\,
            DIN => \N__50507\,
            DOUT => \N__50506\,
            PACKAGEPIN => pwm_output_wire
        );

    \pwm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50508\,
            PADOUT => \N__50507\,
            PADIN => \N__50506\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__24476\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50499\,
            DIN => \N__50498\,
            DOUT => \N__50497\,
            PACKAGEPIN => il_max_comp1_wire
        );

    \il_max_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50499\,
            PADOUT => \N__50498\,
            PADIN => \N__50497\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s2_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50490\,
            DIN => \N__50489\,
            DOUT => \N__50488\,
            PACKAGEPIN => s2_phy_wire
        );

    \s2_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50490\,
            PADOUT => \N__50489\,
            PADIN => \N__50488\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__35870\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T12_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50481\,
            DIN => \N__50480\,
            DOUT => \N__50479\,
            PACKAGEPIN => \T12_wire\
        );

    \T12_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50481\,
            PADOUT => \N__50480\,
            PADIN => \N__50479\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__46502\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50472\,
            DIN => \N__50471\,
            DOUT => \N__50470\,
            PACKAGEPIN => il_min_comp2_wire
        );

    \il_min_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50472\,
            PADOUT => \N__50471\,
            PADIN => \N__50470\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s1_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50463\,
            DIN => \N__50462\,
            DOUT => \N__50461\,
            PACKAGEPIN => s1_phy_wire
        );

    \s1_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50463\,
            PADOUT => \N__50462\,
            PADIN => \N__50461\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__35588\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s4_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50454\,
            DIN => \N__50453\,
            DOUT => \N__50452\,
            PACKAGEPIN => s4_phy_wire
        );

    \s4_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50454\,
            PADOUT => \N__50453\,
            PADIN => \N__50452\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__26180\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50445\,
            DIN => \N__50444\,
            DOUT => \N__50443\,
            PACKAGEPIN => il_min_comp1_wire
        );

    \il_min_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50445\,
            PADOUT => \N__50444\,
            PADIN => \N__50443\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s3_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50436\,
            DIN => \N__50435\,
            DOUT => \N__50434\,
            PACKAGEPIN => s3_phy_wire
        );

    \s3_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50436\,
            PADOUT => \N__50435\,
            PADIN => \N__50434\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__26234\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T45_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50427\,
            DIN => \N__50426\,
            DOUT => \N__50425\,
            PACKAGEPIN => \T45_wire\
        );

    \T45_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50427\,
            PADOUT => \N__50426\,
            PADIN => \N__50425\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__31802\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_hc_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50418\,
            DIN => \N__50417\,
            DOUT => \N__50416\,
            PACKAGEPIN => delay_hc_input_wire
        );

    \delay_hc_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50418\,
            PADOUT => \N__50417\,
            PADIN => \N__50416\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_hc_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_tr_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50409\,
            DIN => \N__50408\,
            DOUT => \N__50407\,
            PACKAGEPIN => delay_tr_input_wire
        );

    \delay_tr_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50409\,
            PADOUT => \N__50408\,
            PADIN => \N__50407\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_tr_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__11986\ : InMux
    port map (
            O => \N__50390\,
            I => \N__50387\
        );

    \I__11985\ : LocalMux
    port map (
            O => \N__50387\,
            I => \N__50382\
        );

    \I__11984\ : InMux
    port map (
            O => \N__50386\,
            I => \N__50379\
        );

    \I__11983\ : InMux
    port map (
            O => \N__50385\,
            I => \N__50376\
        );

    \I__11982\ : Span4Mux_v
    port map (
            O => \N__50382\,
            I => \N__50371\
        );

    \I__11981\ : LocalMux
    port map (
            O => \N__50379\,
            I => \N__50371\
        );

    \I__11980\ : LocalMux
    port map (
            O => \N__50376\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26\
        );

    \I__11979\ : Odrv4
    port map (
            O => \N__50371\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26\
        );

    \I__11978\ : InMux
    port map (
            O => \N__50366\,
            I => \N__50363\
        );

    \I__11977\ : LocalMux
    port map (
            O => \N__50363\,
            I => \N__50359\
        );

    \I__11976\ : InMux
    port map (
            O => \N__50362\,
            I => \N__50356\
        );

    \I__11975\ : Span4Mux_v
    port map (
            O => \N__50359\,
            I => \N__50349\
        );

    \I__11974\ : LocalMux
    port map (
            O => \N__50356\,
            I => \N__50349\
        );

    \I__11973\ : InMux
    port map (
            O => \N__50355\,
            I => \N__50346\
        );

    \I__11972\ : InMux
    port map (
            O => \N__50354\,
            I => \N__50343\
        );

    \I__11971\ : Span4Mux_v
    port map (
            O => \N__50349\,
            I => \N__50338\
        );

    \I__11970\ : LocalMux
    port map (
            O => \N__50346\,
            I => \N__50338\
        );

    \I__11969\ : LocalMux
    port map (
            O => \N__50343\,
            I => \N__50335\
        );

    \I__11968\ : Span4Mux_h
    port map (
            O => \N__50338\,
            I => \N__50332\
        );

    \I__11967\ : Span4Mux_h
    port map (
            O => \N__50335\,
            I => \N__50329\
        );

    \I__11966\ : Odrv4
    port map (
            O => \N__50332\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__11965\ : Odrv4
    port map (
            O => \N__50329\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__11964\ : InMux
    port map (
            O => \N__50324\,
            I => \N__50321\
        );

    \I__11963\ : LocalMux
    port map (
            O => \N__50321\,
            I => \N__50166\
        );

    \I__11962\ : ClkMux
    port map (
            O => \N__50320\,
            I => \N__49856\
        );

    \I__11961\ : ClkMux
    port map (
            O => \N__50319\,
            I => \N__49856\
        );

    \I__11960\ : ClkMux
    port map (
            O => \N__50318\,
            I => \N__49856\
        );

    \I__11959\ : ClkMux
    port map (
            O => \N__50317\,
            I => \N__49856\
        );

    \I__11958\ : ClkMux
    port map (
            O => \N__50316\,
            I => \N__49856\
        );

    \I__11957\ : ClkMux
    port map (
            O => \N__50315\,
            I => \N__49856\
        );

    \I__11956\ : ClkMux
    port map (
            O => \N__50314\,
            I => \N__49856\
        );

    \I__11955\ : ClkMux
    port map (
            O => \N__50313\,
            I => \N__49856\
        );

    \I__11954\ : ClkMux
    port map (
            O => \N__50312\,
            I => \N__49856\
        );

    \I__11953\ : ClkMux
    port map (
            O => \N__50311\,
            I => \N__49856\
        );

    \I__11952\ : ClkMux
    port map (
            O => \N__50310\,
            I => \N__49856\
        );

    \I__11951\ : ClkMux
    port map (
            O => \N__50309\,
            I => \N__49856\
        );

    \I__11950\ : ClkMux
    port map (
            O => \N__50308\,
            I => \N__49856\
        );

    \I__11949\ : ClkMux
    port map (
            O => \N__50307\,
            I => \N__49856\
        );

    \I__11948\ : ClkMux
    port map (
            O => \N__50306\,
            I => \N__49856\
        );

    \I__11947\ : ClkMux
    port map (
            O => \N__50305\,
            I => \N__49856\
        );

    \I__11946\ : ClkMux
    port map (
            O => \N__50304\,
            I => \N__49856\
        );

    \I__11945\ : ClkMux
    port map (
            O => \N__50303\,
            I => \N__49856\
        );

    \I__11944\ : ClkMux
    port map (
            O => \N__50302\,
            I => \N__49856\
        );

    \I__11943\ : ClkMux
    port map (
            O => \N__50301\,
            I => \N__49856\
        );

    \I__11942\ : ClkMux
    port map (
            O => \N__50300\,
            I => \N__49856\
        );

    \I__11941\ : ClkMux
    port map (
            O => \N__50299\,
            I => \N__49856\
        );

    \I__11940\ : ClkMux
    port map (
            O => \N__50298\,
            I => \N__49856\
        );

    \I__11939\ : ClkMux
    port map (
            O => \N__50297\,
            I => \N__49856\
        );

    \I__11938\ : ClkMux
    port map (
            O => \N__50296\,
            I => \N__49856\
        );

    \I__11937\ : ClkMux
    port map (
            O => \N__50295\,
            I => \N__49856\
        );

    \I__11936\ : ClkMux
    port map (
            O => \N__50294\,
            I => \N__49856\
        );

    \I__11935\ : ClkMux
    port map (
            O => \N__50293\,
            I => \N__49856\
        );

    \I__11934\ : ClkMux
    port map (
            O => \N__50292\,
            I => \N__49856\
        );

    \I__11933\ : ClkMux
    port map (
            O => \N__50291\,
            I => \N__49856\
        );

    \I__11932\ : ClkMux
    port map (
            O => \N__50290\,
            I => \N__49856\
        );

    \I__11931\ : ClkMux
    port map (
            O => \N__50289\,
            I => \N__49856\
        );

    \I__11930\ : ClkMux
    port map (
            O => \N__50288\,
            I => \N__49856\
        );

    \I__11929\ : ClkMux
    port map (
            O => \N__50287\,
            I => \N__49856\
        );

    \I__11928\ : ClkMux
    port map (
            O => \N__50286\,
            I => \N__49856\
        );

    \I__11927\ : ClkMux
    port map (
            O => \N__50285\,
            I => \N__49856\
        );

    \I__11926\ : ClkMux
    port map (
            O => \N__50284\,
            I => \N__49856\
        );

    \I__11925\ : ClkMux
    port map (
            O => \N__50283\,
            I => \N__49856\
        );

    \I__11924\ : ClkMux
    port map (
            O => \N__50282\,
            I => \N__49856\
        );

    \I__11923\ : ClkMux
    port map (
            O => \N__50281\,
            I => \N__49856\
        );

    \I__11922\ : ClkMux
    port map (
            O => \N__50280\,
            I => \N__49856\
        );

    \I__11921\ : ClkMux
    port map (
            O => \N__50279\,
            I => \N__49856\
        );

    \I__11920\ : ClkMux
    port map (
            O => \N__50278\,
            I => \N__49856\
        );

    \I__11919\ : ClkMux
    port map (
            O => \N__50277\,
            I => \N__49856\
        );

    \I__11918\ : ClkMux
    port map (
            O => \N__50276\,
            I => \N__49856\
        );

    \I__11917\ : ClkMux
    port map (
            O => \N__50275\,
            I => \N__49856\
        );

    \I__11916\ : ClkMux
    port map (
            O => \N__50274\,
            I => \N__49856\
        );

    \I__11915\ : ClkMux
    port map (
            O => \N__50273\,
            I => \N__49856\
        );

    \I__11914\ : ClkMux
    port map (
            O => \N__50272\,
            I => \N__49856\
        );

    \I__11913\ : ClkMux
    port map (
            O => \N__50271\,
            I => \N__49856\
        );

    \I__11912\ : ClkMux
    port map (
            O => \N__50270\,
            I => \N__49856\
        );

    \I__11911\ : ClkMux
    port map (
            O => \N__50269\,
            I => \N__49856\
        );

    \I__11910\ : ClkMux
    port map (
            O => \N__50268\,
            I => \N__49856\
        );

    \I__11909\ : ClkMux
    port map (
            O => \N__50267\,
            I => \N__49856\
        );

    \I__11908\ : ClkMux
    port map (
            O => \N__50266\,
            I => \N__49856\
        );

    \I__11907\ : ClkMux
    port map (
            O => \N__50265\,
            I => \N__49856\
        );

    \I__11906\ : ClkMux
    port map (
            O => \N__50264\,
            I => \N__49856\
        );

    \I__11905\ : ClkMux
    port map (
            O => \N__50263\,
            I => \N__49856\
        );

    \I__11904\ : ClkMux
    port map (
            O => \N__50262\,
            I => \N__49856\
        );

    \I__11903\ : ClkMux
    port map (
            O => \N__50261\,
            I => \N__49856\
        );

    \I__11902\ : ClkMux
    port map (
            O => \N__50260\,
            I => \N__49856\
        );

    \I__11901\ : ClkMux
    port map (
            O => \N__50259\,
            I => \N__49856\
        );

    \I__11900\ : ClkMux
    port map (
            O => \N__50258\,
            I => \N__49856\
        );

    \I__11899\ : ClkMux
    port map (
            O => \N__50257\,
            I => \N__49856\
        );

    \I__11898\ : ClkMux
    port map (
            O => \N__50256\,
            I => \N__49856\
        );

    \I__11897\ : ClkMux
    port map (
            O => \N__50255\,
            I => \N__49856\
        );

    \I__11896\ : ClkMux
    port map (
            O => \N__50254\,
            I => \N__49856\
        );

    \I__11895\ : ClkMux
    port map (
            O => \N__50253\,
            I => \N__49856\
        );

    \I__11894\ : ClkMux
    port map (
            O => \N__50252\,
            I => \N__49856\
        );

    \I__11893\ : ClkMux
    port map (
            O => \N__50251\,
            I => \N__49856\
        );

    \I__11892\ : ClkMux
    port map (
            O => \N__50250\,
            I => \N__49856\
        );

    \I__11891\ : ClkMux
    port map (
            O => \N__50249\,
            I => \N__49856\
        );

    \I__11890\ : ClkMux
    port map (
            O => \N__50248\,
            I => \N__49856\
        );

    \I__11889\ : ClkMux
    port map (
            O => \N__50247\,
            I => \N__49856\
        );

    \I__11888\ : ClkMux
    port map (
            O => \N__50246\,
            I => \N__49856\
        );

    \I__11887\ : ClkMux
    port map (
            O => \N__50245\,
            I => \N__49856\
        );

    \I__11886\ : ClkMux
    port map (
            O => \N__50244\,
            I => \N__49856\
        );

    \I__11885\ : ClkMux
    port map (
            O => \N__50243\,
            I => \N__49856\
        );

    \I__11884\ : ClkMux
    port map (
            O => \N__50242\,
            I => \N__49856\
        );

    \I__11883\ : ClkMux
    port map (
            O => \N__50241\,
            I => \N__49856\
        );

    \I__11882\ : ClkMux
    port map (
            O => \N__50240\,
            I => \N__49856\
        );

    \I__11881\ : ClkMux
    port map (
            O => \N__50239\,
            I => \N__49856\
        );

    \I__11880\ : ClkMux
    port map (
            O => \N__50238\,
            I => \N__49856\
        );

    \I__11879\ : ClkMux
    port map (
            O => \N__50237\,
            I => \N__49856\
        );

    \I__11878\ : ClkMux
    port map (
            O => \N__50236\,
            I => \N__49856\
        );

    \I__11877\ : ClkMux
    port map (
            O => \N__50235\,
            I => \N__49856\
        );

    \I__11876\ : ClkMux
    port map (
            O => \N__50234\,
            I => \N__49856\
        );

    \I__11875\ : ClkMux
    port map (
            O => \N__50233\,
            I => \N__49856\
        );

    \I__11874\ : ClkMux
    port map (
            O => \N__50232\,
            I => \N__49856\
        );

    \I__11873\ : ClkMux
    port map (
            O => \N__50231\,
            I => \N__49856\
        );

    \I__11872\ : ClkMux
    port map (
            O => \N__50230\,
            I => \N__49856\
        );

    \I__11871\ : ClkMux
    port map (
            O => \N__50229\,
            I => \N__49856\
        );

    \I__11870\ : ClkMux
    port map (
            O => \N__50228\,
            I => \N__49856\
        );

    \I__11869\ : ClkMux
    port map (
            O => \N__50227\,
            I => \N__49856\
        );

    \I__11868\ : ClkMux
    port map (
            O => \N__50226\,
            I => \N__49856\
        );

    \I__11867\ : ClkMux
    port map (
            O => \N__50225\,
            I => \N__49856\
        );

    \I__11866\ : ClkMux
    port map (
            O => \N__50224\,
            I => \N__49856\
        );

    \I__11865\ : ClkMux
    port map (
            O => \N__50223\,
            I => \N__49856\
        );

    \I__11864\ : ClkMux
    port map (
            O => \N__50222\,
            I => \N__49856\
        );

    \I__11863\ : ClkMux
    port map (
            O => \N__50221\,
            I => \N__49856\
        );

    \I__11862\ : ClkMux
    port map (
            O => \N__50220\,
            I => \N__49856\
        );

    \I__11861\ : ClkMux
    port map (
            O => \N__50219\,
            I => \N__49856\
        );

    \I__11860\ : ClkMux
    port map (
            O => \N__50218\,
            I => \N__49856\
        );

    \I__11859\ : ClkMux
    port map (
            O => \N__50217\,
            I => \N__49856\
        );

    \I__11858\ : ClkMux
    port map (
            O => \N__50216\,
            I => \N__49856\
        );

    \I__11857\ : ClkMux
    port map (
            O => \N__50215\,
            I => \N__49856\
        );

    \I__11856\ : ClkMux
    port map (
            O => \N__50214\,
            I => \N__49856\
        );

    \I__11855\ : ClkMux
    port map (
            O => \N__50213\,
            I => \N__49856\
        );

    \I__11854\ : ClkMux
    port map (
            O => \N__50212\,
            I => \N__49856\
        );

    \I__11853\ : ClkMux
    port map (
            O => \N__50211\,
            I => \N__49856\
        );

    \I__11852\ : ClkMux
    port map (
            O => \N__50210\,
            I => \N__49856\
        );

    \I__11851\ : ClkMux
    port map (
            O => \N__50209\,
            I => \N__49856\
        );

    \I__11850\ : ClkMux
    port map (
            O => \N__50208\,
            I => \N__49856\
        );

    \I__11849\ : ClkMux
    port map (
            O => \N__50207\,
            I => \N__49856\
        );

    \I__11848\ : ClkMux
    port map (
            O => \N__50206\,
            I => \N__49856\
        );

    \I__11847\ : ClkMux
    port map (
            O => \N__50205\,
            I => \N__49856\
        );

    \I__11846\ : ClkMux
    port map (
            O => \N__50204\,
            I => \N__49856\
        );

    \I__11845\ : ClkMux
    port map (
            O => \N__50203\,
            I => \N__49856\
        );

    \I__11844\ : ClkMux
    port map (
            O => \N__50202\,
            I => \N__49856\
        );

    \I__11843\ : ClkMux
    port map (
            O => \N__50201\,
            I => \N__49856\
        );

    \I__11842\ : ClkMux
    port map (
            O => \N__50200\,
            I => \N__49856\
        );

    \I__11841\ : ClkMux
    port map (
            O => \N__50199\,
            I => \N__49856\
        );

    \I__11840\ : ClkMux
    port map (
            O => \N__50198\,
            I => \N__49856\
        );

    \I__11839\ : ClkMux
    port map (
            O => \N__50197\,
            I => \N__49856\
        );

    \I__11838\ : ClkMux
    port map (
            O => \N__50196\,
            I => \N__49856\
        );

    \I__11837\ : ClkMux
    port map (
            O => \N__50195\,
            I => \N__49856\
        );

    \I__11836\ : ClkMux
    port map (
            O => \N__50194\,
            I => \N__49856\
        );

    \I__11835\ : ClkMux
    port map (
            O => \N__50193\,
            I => \N__49856\
        );

    \I__11834\ : ClkMux
    port map (
            O => \N__50192\,
            I => \N__49856\
        );

    \I__11833\ : ClkMux
    port map (
            O => \N__50191\,
            I => \N__49856\
        );

    \I__11832\ : ClkMux
    port map (
            O => \N__50190\,
            I => \N__49856\
        );

    \I__11831\ : ClkMux
    port map (
            O => \N__50189\,
            I => \N__49856\
        );

    \I__11830\ : ClkMux
    port map (
            O => \N__50188\,
            I => \N__49856\
        );

    \I__11829\ : ClkMux
    port map (
            O => \N__50187\,
            I => \N__49856\
        );

    \I__11828\ : ClkMux
    port map (
            O => \N__50186\,
            I => \N__49856\
        );

    \I__11827\ : ClkMux
    port map (
            O => \N__50185\,
            I => \N__49856\
        );

    \I__11826\ : ClkMux
    port map (
            O => \N__50184\,
            I => \N__49856\
        );

    \I__11825\ : ClkMux
    port map (
            O => \N__50183\,
            I => \N__49856\
        );

    \I__11824\ : ClkMux
    port map (
            O => \N__50182\,
            I => \N__49856\
        );

    \I__11823\ : ClkMux
    port map (
            O => \N__50181\,
            I => \N__49856\
        );

    \I__11822\ : ClkMux
    port map (
            O => \N__50180\,
            I => \N__49856\
        );

    \I__11821\ : ClkMux
    port map (
            O => \N__50179\,
            I => \N__49856\
        );

    \I__11820\ : ClkMux
    port map (
            O => \N__50178\,
            I => \N__49856\
        );

    \I__11819\ : ClkMux
    port map (
            O => \N__50177\,
            I => \N__49856\
        );

    \I__11818\ : ClkMux
    port map (
            O => \N__50176\,
            I => \N__49856\
        );

    \I__11817\ : ClkMux
    port map (
            O => \N__50175\,
            I => \N__49856\
        );

    \I__11816\ : ClkMux
    port map (
            O => \N__50174\,
            I => \N__49856\
        );

    \I__11815\ : ClkMux
    port map (
            O => \N__50173\,
            I => \N__49856\
        );

    \I__11814\ : ClkMux
    port map (
            O => \N__50172\,
            I => \N__49856\
        );

    \I__11813\ : ClkMux
    port map (
            O => \N__50171\,
            I => \N__49856\
        );

    \I__11812\ : ClkMux
    port map (
            O => \N__50170\,
            I => \N__49856\
        );

    \I__11811\ : ClkMux
    port map (
            O => \N__50169\,
            I => \N__49856\
        );

    \I__11810\ : Glb2LocalMux
    port map (
            O => \N__50166\,
            I => \N__49856\
        );

    \I__11809\ : ClkMux
    port map (
            O => \N__50165\,
            I => \N__49856\
        );

    \I__11808\ : GlobalMux
    port map (
            O => \N__49856\,
            I => clock_output_0
        );

    \I__11807\ : InMux
    port map (
            O => \N__49853\,
            I => \N__49840\
        );

    \I__11806\ : InMux
    port map (
            O => \N__49852\,
            I => \N__49840\
        );

    \I__11805\ : InMux
    port map (
            O => \N__49851\,
            I => \N__49840\
        );

    \I__11804\ : InMux
    port map (
            O => \N__49850\,
            I => \N__49823\
        );

    \I__11803\ : InMux
    port map (
            O => \N__49849\,
            I => \N__49823\
        );

    \I__11802\ : InMux
    port map (
            O => \N__49848\,
            I => \N__49823\
        );

    \I__11801\ : InMux
    port map (
            O => \N__49847\,
            I => \N__49823\
        );

    \I__11800\ : LocalMux
    port map (
            O => \N__49840\,
            I => \N__49820\
        );

    \I__11799\ : InMux
    port map (
            O => \N__49839\,
            I => \N__49811\
        );

    \I__11798\ : InMux
    port map (
            O => \N__49838\,
            I => \N__49811\
        );

    \I__11797\ : InMux
    port map (
            O => \N__49837\,
            I => \N__49811\
        );

    \I__11796\ : InMux
    port map (
            O => \N__49836\,
            I => \N__49811\
        );

    \I__11795\ : CEMux
    port map (
            O => \N__49835\,
            I => \N__49808\
        );

    \I__11794\ : CEMux
    port map (
            O => \N__49834\,
            I => \N__49800\
        );

    \I__11793\ : InMux
    port map (
            O => \N__49833\,
            I => \N__49796\
        );

    \I__11792\ : CEMux
    port map (
            O => \N__49832\,
            I => \N__49793\
        );

    \I__11791\ : LocalMux
    port map (
            O => \N__49823\,
            I => \N__49781\
        );

    \I__11790\ : Span4Mux_h
    port map (
            O => \N__49820\,
            I => \N__49781\
        );

    \I__11789\ : LocalMux
    port map (
            O => \N__49811\,
            I => \N__49781\
        );

    \I__11788\ : LocalMux
    port map (
            O => \N__49808\,
            I => \N__49778\
        );

    \I__11787\ : CEMux
    port map (
            O => \N__49807\,
            I => \N__49763\
        );

    \I__11786\ : CEMux
    port map (
            O => \N__49806\,
            I => \N__49760\
        );

    \I__11785\ : CEMux
    port map (
            O => \N__49805\,
            I => \N__49757\
        );

    \I__11784\ : CEMux
    port map (
            O => \N__49804\,
            I => \N__49754\
        );

    \I__11783\ : CEMux
    port map (
            O => \N__49803\,
            I => \N__49751\
        );

    \I__11782\ : LocalMux
    port map (
            O => \N__49800\,
            I => \N__49748\
        );

    \I__11781\ : CEMux
    port map (
            O => \N__49799\,
            I => \N__49741\
        );

    \I__11780\ : LocalMux
    port map (
            O => \N__49796\,
            I => \N__49736\
        );

    \I__11779\ : LocalMux
    port map (
            O => \N__49793\,
            I => \N__49736\
        );

    \I__11778\ : CEMux
    port map (
            O => \N__49792\,
            I => \N__49730\
        );

    \I__11777\ : CEMux
    port map (
            O => \N__49791\,
            I => \N__49727\
        );

    \I__11776\ : InMux
    port map (
            O => \N__49790\,
            I => \N__49720\
        );

    \I__11775\ : InMux
    port map (
            O => \N__49789\,
            I => \N__49720\
        );

    \I__11774\ : InMux
    port map (
            O => \N__49788\,
            I => \N__49720\
        );

    \I__11773\ : Span4Mux_v
    port map (
            O => \N__49781\,
            I => \N__49715\
        );

    \I__11772\ : Span4Mux_v
    port map (
            O => \N__49778\,
            I => \N__49715\
        );

    \I__11771\ : InMux
    port map (
            O => \N__49777\,
            I => \N__49706\
        );

    \I__11770\ : InMux
    port map (
            O => \N__49776\,
            I => \N__49706\
        );

    \I__11769\ : InMux
    port map (
            O => \N__49775\,
            I => \N__49706\
        );

    \I__11768\ : InMux
    port map (
            O => \N__49774\,
            I => \N__49706\
        );

    \I__11767\ : InMux
    port map (
            O => \N__49773\,
            I => \N__49697\
        );

    \I__11766\ : InMux
    port map (
            O => \N__49772\,
            I => \N__49697\
        );

    \I__11765\ : InMux
    port map (
            O => \N__49771\,
            I => \N__49697\
        );

    \I__11764\ : InMux
    port map (
            O => \N__49770\,
            I => \N__49697\
        );

    \I__11763\ : InMux
    port map (
            O => \N__49769\,
            I => \N__49688\
        );

    \I__11762\ : InMux
    port map (
            O => \N__49768\,
            I => \N__49688\
        );

    \I__11761\ : InMux
    port map (
            O => \N__49767\,
            I => \N__49688\
        );

    \I__11760\ : InMux
    port map (
            O => \N__49766\,
            I => \N__49688\
        );

    \I__11759\ : LocalMux
    port map (
            O => \N__49763\,
            I => \N__49685\
        );

    \I__11758\ : LocalMux
    port map (
            O => \N__49760\,
            I => \N__49680\
        );

    \I__11757\ : LocalMux
    port map (
            O => \N__49757\,
            I => \N__49680\
        );

    \I__11756\ : LocalMux
    port map (
            O => \N__49754\,
            I => \N__49677\
        );

    \I__11755\ : LocalMux
    port map (
            O => \N__49751\,
            I => \N__49672\
        );

    \I__11754\ : Span4Mux_h
    port map (
            O => \N__49748\,
            I => \N__49672\
        );

    \I__11753\ : InMux
    port map (
            O => \N__49747\,
            I => \N__49663\
        );

    \I__11752\ : InMux
    port map (
            O => \N__49746\,
            I => \N__49663\
        );

    \I__11751\ : InMux
    port map (
            O => \N__49745\,
            I => \N__49663\
        );

    \I__11750\ : InMux
    port map (
            O => \N__49744\,
            I => \N__49663\
        );

    \I__11749\ : LocalMux
    port map (
            O => \N__49741\,
            I => \N__49660\
        );

    \I__11748\ : Span4Mux_v
    port map (
            O => \N__49736\,
            I => \N__49657\
        );

    \I__11747\ : CEMux
    port map (
            O => \N__49735\,
            I => \N__49654\
        );

    \I__11746\ : CEMux
    port map (
            O => \N__49734\,
            I => \N__49651\
        );

    \I__11745\ : CEMux
    port map (
            O => \N__49733\,
            I => \N__49648\
        );

    \I__11744\ : LocalMux
    port map (
            O => \N__49730\,
            I => \N__49645\
        );

    \I__11743\ : LocalMux
    port map (
            O => \N__49727\,
            I => \N__49642\
        );

    \I__11742\ : LocalMux
    port map (
            O => \N__49720\,
            I => \N__49631\
        );

    \I__11741\ : Span4Mux_h
    port map (
            O => \N__49715\,
            I => \N__49631\
        );

    \I__11740\ : LocalMux
    port map (
            O => \N__49706\,
            I => \N__49631\
        );

    \I__11739\ : LocalMux
    port map (
            O => \N__49697\,
            I => \N__49631\
        );

    \I__11738\ : LocalMux
    port map (
            O => \N__49688\,
            I => \N__49631\
        );

    \I__11737\ : Span4Mux_h
    port map (
            O => \N__49685\,
            I => \N__49628\
        );

    \I__11736\ : Sp12to4
    port map (
            O => \N__49680\,
            I => \N__49625\
        );

    \I__11735\ : Span4Mux_v
    port map (
            O => \N__49677\,
            I => \N__49614\
        );

    \I__11734\ : Span4Mux_v
    port map (
            O => \N__49672\,
            I => \N__49614\
        );

    \I__11733\ : LocalMux
    port map (
            O => \N__49663\,
            I => \N__49614\
        );

    \I__11732\ : Span4Mux_v
    port map (
            O => \N__49660\,
            I => \N__49614\
        );

    \I__11731\ : Span4Mux_h
    port map (
            O => \N__49657\,
            I => \N__49614\
        );

    \I__11730\ : LocalMux
    port map (
            O => \N__49654\,
            I => \N__49611\
        );

    \I__11729\ : LocalMux
    port map (
            O => \N__49651\,
            I => \N__49608\
        );

    \I__11728\ : LocalMux
    port map (
            O => \N__49648\,
            I => \N__49603\
        );

    \I__11727\ : Span4Mux_h
    port map (
            O => \N__49645\,
            I => \N__49603\
        );

    \I__11726\ : Span4Mux_h
    port map (
            O => \N__49642\,
            I => \N__49598\
        );

    \I__11725\ : Span4Mux_v
    port map (
            O => \N__49631\,
            I => \N__49598\
        );

    \I__11724\ : Span4Mux_h
    port map (
            O => \N__49628\,
            I => \N__49595\
        );

    \I__11723\ : Span12Mux_s9_v
    port map (
            O => \N__49625\,
            I => \N__49592\
        );

    \I__11722\ : Span4Mux_h
    port map (
            O => \N__49614\,
            I => \N__49589\
        );

    \I__11721\ : Odrv4
    port map (
            O => \N__49611\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__11720\ : Odrv12
    port map (
            O => \N__49608\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__11719\ : Odrv4
    port map (
            O => \N__49603\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__11718\ : Odrv4
    port map (
            O => \N__49598\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__11717\ : Odrv4
    port map (
            O => \N__49595\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__11716\ : Odrv12
    port map (
            O => \N__49592\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__11715\ : Odrv4
    port map (
            O => \N__49589\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__11714\ : InMux
    port map (
            O => \N__49574\,
            I => \N__49568\
        );

    \I__11713\ : InMux
    port map (
            O => \N__49573\,
            I => \N__49565\
        );

    \I__11712\ : InMux
    port map (
            O => \N__49572\,
            I => \N__49562\
        );

    \I__11711\ : InMux
    port map (
            O => \N__49571\,
            I => \N__49559\
        );

    \I__11710\ : LocalMux
    port map (
            O => \N__49568\,
            I => \N__49556\
        );

    \I__11709\ : LocalMux
    port map (
            O => \N__49565\,
            I => \N__49553\
        );

    \I__11708\ : LocalMux
    port map (
            O => \N__49562\,
            I => \N__49545\
        );

    \I__11707\ : LocalMux
    port map (
            O => \N__49559\,
            I => \N__49541\
        );

    \I__11706\ : Glb2LocalMux
    port map (
            O => \N__49556\,
            I => \N__49076\
        );

    \I__11705\ : Glb2LocalMux
    port map (
            O => \N__49553\,
            I => \N__49076\
        );

    \I__11704\ : SRMux
    port map (
            O => \N__49552\,
            I => \N__49076\
        );

    \I__11703\ : SRMux
    port map (
            O => \N__49551\,
            I => \N__49076\
        );

    \I__11702\ : SRMux
    port map (
            O => \N__49550\,
            I => \N__49076\
        );

    \I__11701\ : SRMux
    port map (
            O => \N__49549\,
            I => \N__49076\
        );

    \I__11700\ : SRMux
    port map (
            O => \N__49548\,
            I => \N__49076\
        );

    \I__11699\ : Glb2LocalMux
    port map (
            O => \N__49545\,
            I => \N__49076\
        );

    \I__11698\ : SRMux
    port map (
            O => \N__49544\,
            I => \N__49076\
        );

    \I__11697\ : Glb2LocalMux
    port map (
            O => \N__49541\,
            I => \N__49076\
        );

    \I__11696\ : SRMux
    port map (
            O => \N__49540\,
            I => \N__49076\
        );

    \I__11695\ : SRMux
    port map (
            O => \N__49539\,
            I => \N__49076\
        );

    \I__11694\ : SRMux
    port map (
            O => \N__49538\,
            I => \N__49076\
        );

    \I__11693\ : SRMux
    port map (
            O => \N__49537\,
            I => \N__49076\
        );

    \I__11692\ : SRMux
    port map (
            O => \N__49536\,
            I => \N__49076\
        );

    \I__11691\ : SRMux
    port map (
            O => \N__49535\,
            I => \N__49076\
        );

    \I__11690\ : SRMux
    port map (
            O => \N__49534\,
            I => \N__49076\
        );

    \I__11689\ : SRMux
    port map (
            O => \N__49533\,
            I => \N__49076\
        );

    \I__11688\ : SRMux
    port map (
            O => \N__49532\,
            I => \N__49076\
        );

    \I__11687\ : SRMux
    port map (
            O => \N__49531\,
            I => \N__49076\
        );

    \I__11686\ : SRMux
    port map (
            O => \N__49530\,
            I => \N__49076\
        );

    \I__11685\ : SRMux
    port map (
            O => \N__49529\,
            I => \N__49076\
        );

    \I__11684\ : SRMux
    port map (
            O => \N__49528\,
            I => \N__49076\
        );

    \I__11683\ : SRMux
    port map (
            O => \N__49527\,
            I => \N__49076\
        );

    \I__11682\ : SRMux
    port map (
            O => \N__49526\,
            I => \N__49076\
        );

    \I__11681\ : SRMux
    port map (
            O => \N__49525\,
            I => \N__49076\
        );

    \I__11680\ : SRMux
    port map (
            O => \N__49524\,
            I => \N__49076\
        );

    \I__11679\ : SRMux
    port map (
            O => \N__49523\,
            I => \N__49076\
        );

    \I__11678\ : SRMux
    port map (
            O => \N__49522\,
            I => \N__49076\
        );

    \I__11677\ : SRMux
    port map (
            O => \N__49521\,
            I => \N__49076\
        );

    \I__11676\ : SRMux
    port map (
            O => \N__49520\,
            I => \N__49076\
        );

    \I__11675\ : SRMux
    port map (
            O => \N__49519\,
            I => \N__49076\
        );

    \I__11674\ : SRMux
    port map (
            O => \N__49518\,
            I => \N__49076\
        );

    \I__11673\ : SRMux
    port map (
            O => \N__49517\,
            I => \N__49076\
        );

    \I__11672\ : SRMux
    port map (
            O => \N__49516\,
            I => \N__49076\
        );

    \I__11671\ : SRMux
    port map (
            O => \N__49515\,
            I => \N__49076\
        );

    \I__11670\ : SRMux
    port map (
            O => \N__49514\,
            I => \N__49076\
        );

    \I__11669\ : SRMux
    port map (
            O => \N__49513\,
            I => \N__49076\
        );

    \I__11668\ : SRMux
    port map (
            O => \N__49512\,
            I => \N__49076\
        );

    \I__11667\ : SRMux
    port map (
            O => \N__49511\,
            I => \N__49076\
        );

    \I__11666\ : SRMux
    port map (
            O => \N__49510\,
            I => \N__49076\
        );

    \I__11665\ : SRMux
    port map (
            O => \N__49509\,
            I => \N__49076\
        );

    \I__11664\ : SRMux
    port map (
            O => \N__49508\,
            I => \N__49076\
        );

    \I__11663\ : SRMux
    port map (
            O => \N__49507\,
            I => \N__49076\
        );

    \I__11662\ : SRMux
    port map (
            O => \N__49506\,
            I => \N__49076\
        );

    \I__11661\ : SRMux
    port map (
            O => \N__49505\,
            I => \N__49076\
        );

    \I__11660\ : SRMux
    port map (
            O => \N__49504\,
            I => \N__49076\
        );

    \I__11659\ : SRMux
    port map (
            O => \N__49503\,
            I => \N__49076\
        );

    \I__11658\ : SRMux
    port map (
            O => \N__49502\,
            I => \N__49076\
        );

    \I__11657\ : SRMux
    port map (
            O => \N__49501\,
            I => \N__49076\
        );

    \I__11656\ : SRMux
    port map (
            O => \N__49500\,
            I => \N__49076\
        );

    \I__11655\ : SRMux
    port map (
            O => \N__49499\,
            I => \N__49076\
        );

    \I__11654\ : SRMux
    port map (
            O => \N__49498\,
            I => \N__49076\
        );

    \I__11653\ : SRMux
    port map (
            O => \N__49497\,
            I => \N__49076\
        );

    \I__11652\ : SRMux
    port map (
            O => \N__49496\,
            I => \N__49076\
        );

    \I__11651\ : SRMux
    port map (
            O => \N__49495\,
            I => \N__49076\
        );

    \I__11650\ : SRMux
    port map (
            O => \N__49494\,
            I => \N__49076\
        );

    \I__11649\ : SRMux
    port map (
            O => \N__49493\,
            I => \N__49076\
        );

    \I__11648\ : SRMux
    port map (
            O => \N__49492\,
            I => \N__49076\
        );

    \I__11647\ : SRMux
    port map (
            O => \N__49491\,
            I => \N__49076\
        );

    \I__11646\ : SRMux
    port map (
            O => \N__49490\,
            I => \N__49076\
        );

    \I__11645\ : SRMux
    port map (
            O => \N__49489\,
            I => \N__49076\
        );

    \I__11644\ : SRMux
    port map (
            O => \N__49488\,
            I => \N__49076\
        );

    \I__11643\ : SRMux
    port map (
            O => \N__49487\,
            I => \N__49076\
        );

    \I__11642\ : SRMux
    port map (
            O => \N__49486\,
            I => \N__49076\
        );

    \I__11641\ : SRMux
    port map (
            O => \N__49485\,
            I => \N__49076\
        );

    \I__11640\ : SRMux
    port map (
            O => \N__49484\,
            I => \N__49076\
        );

    \I__11639\ : SRMux
    port map (
            O => \N__49483\,
            I => \N__49076\
        );

    \I__11638\ : SRMux
    port map (
            O => \N__49482\,
            I => \N__49076\
        );

    \I__11637\ : SRMux
    port map (
            O => \N__49481\,
            I => \N__49076\
        );

    \I__11636\ : SRMux
    port map (
            O => \N__49480\,
            I => \N__49076\
        );

    \I__11635\ : SRMux
    port map (
            O => \N__49479\,
            I => \N__49076\
        );

    \I__11634\ : SRMux
    port map (
            O => \N__49478\,
            I => \N__49076\
        );

    \I__11633\ : SRMux
    port map (
            O => \N__49477\,
            I => \N__49076\
        );

    \I__11632\ : SRMux
    port map (
            O => \N__49476\,
            I => \N__49076\
        );

    \I__11631\ : SRMux
    port map (
            O => \N__49475\,
            I => \N__49076\
        );

    \I__11630\ : SRMux
    port map (
            O => \N__49474\,
            I => \N__49076\
        );

    \I__11629\ : SRMux
    port map (
            O => \N__49473\,
            I => \N__49076\
        );

    \I__11628\ : SRMux
    port map (
            O => \N__49472\,
            I => \N__49076\
        );

    \I__11627\ : SRMux
    port map (
            O => \N__49471\,
            I => \N__49076\
        );

    \I__11626\ : SRMux
    port map (
            O => \N__49470\,
            I => \N__49076\
        );

    \I__11625\ : SRMux
    port map (
            O => \N__49469\,
            I => \N__49076\
        );

    \I__11624\ : SRMux
    port map (
            O => \N__49468\,
            I => \N__49076\
        );

    \I__11623\ : SRMux
    port map (
            O => \N__49467\,
            I => \N__49076\
        );

    \I__11622\ : SRMux
    port map (
            O => \N__49466\,
            I => \N__49076\
        );

    \I__11621\ : SRMux
    port map (
            O => \N__49465\,
            I => \N__49076\
        );

    \I__11620\ : SRMux
    port map (
            O => \N__49464\,
            I => \N__49076\
        );

    \I__11619\ : SRMux
    port map (
            O => \N__49463\,
            I => \N__49076\
        );

    \I__11618\ : SRMux
    port map (
            O => \N__49462\,
            I => \N__49076\
        );

    \I__11617\ : SRMux
    port map (
            O => \N__49461\,
            I => \N__49076\
        );

    \I__11616\ : SRMux
    port map (
            O => \N__49460\,
            I => \N__49076\
        );

    \I__11615\ : SRMux
    port map (
            O => \N__49459\,
            I => \N__49076\
        );

    \I__11614\ : SRMux
    port map (
            O => \N__49458\,
            I => \N__49076\
        );

    \I__11613\ : SRMux
    port map (
            O => \N__49457\,
            I => \N__49076\
        );

    \I__11612\ : SRMux
    port map (
            O => \N__49456\,
            I => \N__49076\
        );

    \I__11611\ : SRMux
    port map (
            O => \N__49455\,
            I => \N__49076\
        );

    \I__11610\ : SRMux
    port map (
            O => \N__49454\,
            I => \N__49076\
        );

    \I__11609\ : SRMux
    port map (
            O => \N__49453\,
            I => \N__49076\
        );

    \I__11608\ : SRMux
    port map (
            O => \N__49452\,
            I => \N__49076\
        );

    \I__11607\ : SRMux
    port map (
            O => \N__49451\,
            I => \N__49076\
        );

    \I__11606\ : SRMux
    port map (
            O => \N__49450\,
            I => \N__49076\
        );

    \I__11605\ : SRMux
    port map (
            O => \N__49449\,
            I => \N__49076\
        );

    \I__11604\ : SRMux
    port map (
            O => \N__49448\,
            I => \N__49076\
        );

    \I__11603\ : SRMux
    port map (
            O => \N__49447\,
            I => \N__49076\
        );

    \I__11602\ : SRMux
    port map (
            O => \N__49446\,
            I => \N__49076\
        );

    \I__11601\ : SRMux
    port map (
            O => \N__49445\,
            I => \N__49076\
        );

    \I__11600\ : SRMux
    port map (
            O => \N__49444\,
            I => \N__49076\
        );

    \I__11599\ : SRMux
    port map (
            O => \N__49443\,
            I => \N__49076\
        );

    \I__11598\ : SRMux
    port map (
            O => \N__49442\,
            I => \N__49076\
        );

    \I__11597\ : SRMux
    port map (
            O => \N__49441\,
            I => \N__49076\
        );

    \I__11596\ : SRMux
    port map (
            O => \N__49440\,
            I => \N__49076\
        );

    \I__11595\ : SRMux
    port map (
            O => \N__49439\,
            I => \N__49076\
        );

    \I__11594\ : SRMux
    port map (
            O => \N__49438\,
            I => \N__49076\
        );

    \I__11593\ : SRMux
    port map (
            O => \N__49437\,
            I => \N__49076\
        );

    \I__11592\ : SRMux
    port map (
            O => \N__49436\,
            I => \N__49076\
        );

    \I__11591\ : SRMux
    port map (
            O => \N__49435\,
            I => \N__49076\
        );

    \I__11590\ : SRMux
    port map (
            O => \N__49434\,
            I => \N__49076\
        );

    \I__11589\ : SRMux
    port map (
            O => \N__49433\,
            I => \N__49076\
        );

    \I__11588\ : SRMux
    port map (
            O => \N__49432\,
            I => \N__49076\
        );

    \I__11587\ : SRMux
    port map (
            O => \N__49431\,
            I => \N__49076\
        );

    \I__11586\ : SRMux
    port map (
            O => \N__49430\,
            I => \N__49076\
        );

    \I__11585\ : SRMux
    port map (
            O => \N__49429\,
            I => \N__49076\
        );

    \I__11584\ : SRMux
    port map (
            O => \N__49428\,
            I => \N__49076\
        );

    \I__11583\ : SRMux
    port map (
            O => \N__49427\,
            I => \N__49076\
        );

    \I__11582\ : SRMux
    port map (
            O => \N__49426\,
            I => \N__49076\
        );

    \I__11581\ : SRMux
    port map (
            O => \N__49425\,
            I => \N__49076\
        );

    \I__11580\ : SRMux
    port map (
            O => \N__49424\,
            I => \N__49076\
        );

    \I__11579\ : SRMux
    port map (
            O => \N__49423\,
            I => \N__49076\
        );

    \I__11578\ : SRMux
    port map (
            O => \N__49422\,
            I => \N__49076\
        );

    \I__11577\ : SRMux
    port map (
            O => \N__49421\,
            I => \N__49076\
        );

    \I__11576\ : SRMux
    port map (
            O => \N__49420\,
            I => \N__49076\
        );

    \I__11575\ : SRMux
    port map (
            O => \N__49419\,
            I => \N__49076\
        );

    \I__11574\ : SRMux
    port map (
            O => \N__49418\,
            I => \N__49076\
        );

    \I__11573\ : SRMux
    port map (
            O => \N__49417\,
            I => \N__49076\
        );

    \I__11572\ : SRMux
    port map (
            O => \N__49416\,
            I => \N__49076\
        );

    \I__11571\ : SRMux
    port map (
            O => \N__49415\,
            I => \N__49076\
        );

    \I__11570\ : SRMux
    port map (
            O => \N__49414\,
            I => \N__49076\
        );

    \I__11569\ : SRMux
    port map (
            O => \N__49413\,
            I => \N__49076\
        );

    \I__11568\ : SRMux
    port map (
            O => \N__49412\,
            I => \N__49076\
        );

    \I__11567\ : SRMux
    port map (
            O => \N__49411\,
            I => \N__49076\
        );

    \I__11566\ : SRMux
    port map (
            O => \N__49410\,
            I => \N__49076\
        );

    \I__11565\ : SRMux
    port map (
            O => \N__49409\,
            I => \N__49076\
        );

    \I__11564\ : SRMux
    port map (
            O => \N__49408\,
            I => \N__49076\
        );

    \I__11563\ : SRMux
    port map (
            O => \N__49407\,
            I => \N__49076\
        );

    \I__11562\ : SRMux
    port map (
            O => \N__49406\,
            I => \N__49076\
        );

    \I__11561\ : SRMux
    port map (
            O => \N__49405\,
            I => \N__49076\
        );

    \I__11560\ : SRMux
    port map (
            O => \N__49404\,
            I => \N__49076\
        );

    \I__11559\ : SRMux
    port map (
            O => \N__49403\,
            I => \N__49076\
        );

    \I__11558\ : SRMux
    port map (
            O => \N__49402\,
            I => \N__49076\
        );

    \I__11557\ : SRMux
    port map (
            O => \N__49401\,
            I => \N__49076\
        );

    \I__11556\ : SRMux
    port map (
            O => \N__49400\,
            I => \N__49076\
        );

    \I__11555\ : SRMux
    port map (
            O => \N__49399\,
            I => \N__49076\
        );

    \I__11554\ : SRMux
    port map (
            O => \N__49398\,
            I => \N__49076\
        );

    \I__11553\ : SRMux
    port map (
            O => \N__49397\,
            I => \N__49076\
        );

    \I__11552\ : SRMux
    port map (
            O => \N__49396\,
            I => \N__49076\
        );

    \I__11551\ : SRMux
    port map (
            O => \N__49395\,
            I => \N__49076\
        );

    \I__11550\ : SRMux
    port map (
            O => \N__49394\,
            I => \N__49076\
        );

    \I__11549\ : SRMux
    port map (
            O => \N__49393\,
            I => \N__49076\
        );

    \I__11548\ : GlobalMux
    port map (
            O => \N__49076\,
            I => \N__49073\
        );

    \I__11547\ : gio2CtrlBuf
    port map (
            O => \N__49073\,
            I => red_c_g
        );

    \I__11546\ : CascadeMux
    port map (
            O => \N__49070\,
            I => \N__49067\
        );

    \I__11545\ : InMux
    port map (
            O => \N__49067\,
            I => \N__49064\
        );

    \I__11544\ : LocalMux
    port map (
            O => \N__49064\,
            I => \N__49061\
        );

    \I__11543\ : Span4Mux_h
    port map (
            O => \N__49061\,
            I => \N__49058\
        );

    \I__11542\ : Odrv4
    port map (
            O => \N__49058\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt26\
        );

    \I__11541\ : InMux
    port map (
            O => \N__49055\,
            I => \N__49049\
        );

    \I__11540\ : InMux
    port map (
            O => \N__49054\,
            I => \N__49049\
        );

    \I__11539\ : LocalMux
    port map (
            O => \N__49049\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_26\
        );

    \I__11538\ : InMux
    port map (
            O => \N__49046\,
            I => \N__49039\
        );

    \I__11537\ : InMux
    port map (
            O => \N__49045\,
            I => \N__49039\
        );

    \I__11536\ : InMux
    port map (
            O => \N__49044\,
            I => \N__49036\
        );

    \I__11535\ : LocalMux
    port map (
            O => \N__49039\,
            I => \N__49033\
        );

    \I__11534\ : LocalMux
    port map (
            O => \N__49036\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__11533\ : Odrv4
    port map (
            O => \N__49033\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__11532\ : CascadeMux
    port map (
            O => \N__49028\,
            I => \N__49024\
        );

    \I__11531\ : CascadeMux
    port map (
            O => \N__49027\,
            I => \N__49021\
        );

    \I__11530\ : InMux
    port map (
            O => \N__49024\,
            I => \N__49015\
        );

    \I__11529\ : InMux
    port map (
            O => \N__49021\,
            I => \N__49015\
        );

    \I__11528\ : InMux
    port map (
            O => \N__49020\,
            I => \N__49012\
        );

    \I__11527\ : LocalMux
    port map (
            O => \N__49015\,
            I => \N__49009\
        );

    \I__11526\ : LocalMux
    port map (
            O => \N__49012\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__11525\ : Odrv4
    port map (
            O => \N__49009\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__11524\ : InMux
    port map (
            O => \N__49004\,
            I => \N__48998\
        );

    \I__11523\ : InMux
    port map (
            O => \N__49003\,
            I => \N__48998\
        );

    \I__11522\ : LocalMux
    port map (
            O => \N__48998\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_27\
        );

    \I__11521\ : InMux
    port map (
            O => \N__48995\,
            I => \N__48992\
        );

    \I__11520\ : LocalMux
    port map (
            O => \N__48992\,
            I => \N__48989\
        );

    \I__11519\ : Span4Mux_h
    port map (
            O => \N__48989\,
            I => \N__48986\
        );

    \I__11518\ : Odrv4
    port map (
            O => \N__48986\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26\
        );

    \I__11517\ : InMux
    port map (
            O => \N__48983\,
            I => \N__48979\
        );

    \I__11516\ : InMux
    port map (
            O => \N__48982\,
            I => \N__48975\
        );

    \I__11515\ : LocalMux
    port map (
            O => \N__48979\,
            I => \N__48972\
        );

    \I__11514\ : InMux
    port map (
            O => \N__48978\,
            I => \N__48969\
        );

    \I__11513\ : LocalMux
    port map (
            O => \N__48975\,
            I => \N__48965\
        );

    \I__11512\ : Span4Mux_v
    port map (
            O => \N__48972\,
            I => \N__48960\
        );

    \I__11511\ : LocalMux
    port map (
            O => \N__48969\,
            I => \N__48960\
        );

    \I__11510\ : InMux
    port map (
            O => \N__48968\,
            I => \N__48957\
        );

    \I__11509\ : Span4Mux_v
    port map (
            O => \N__48965\,
            I => \N__48954\
        );

    \I__11508\ : Span4Mux_v
    port map (
            O => \N__48960\,
            I => \N__48949\
        );

    \I__11507\ : LocalMux
    port map (
            O => \N__48957\,
            I => \N__48949\
        );

    \I__11506\ : Span4Mux_h
    port map (
            O => \N__48954\,
            I => \N__48946\
        );

    \I__11505\ : Span4Mux_h
    port map (
            O => \N__48949\,
            I => \N__48943\
        );

    \I__11504\ : Odrv4
    port map (
            O => \N__48946\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__11503\ : Odrv4
    port map (
            O => \N__48943\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__11502\ : CascadeMux
    port map (
            O => \N__48938\,
            I => \N__48932\
        );

    \I__11501\ : CascadeMux
    port map (
            O => \N__48937\,
            I => \N__48927\
        );

    \I__11500\ : InMux
    port map (
            O => \N__48936\,
            I => \N__48911\
        );

    \I__11499\ : InMux
    port map (
            O => \N__48935\,
            I => \N__48911\
        );

    \I__11498\ : InMux
    port map (
            O => \N__48932\,
            I => \N__48911\
        );

    \I__11497\ : InMux
    port map (
            O => \N__48931\,
            I => \N__48911\
        );

    \I__11496\ : InMux
    port map (
            O => \N__48930\,
            I => \N__48894\
        );

    \I__11495\ : InMux
    port map (
            O => \N__48927\,
            I => \N__48894\
        );

    \I__11494\ : InMux
    port map (
            O => \N__48926\,
            I => \N__48894\
        );

    \I__11493\ : InMux
    port map (
            O => \N__48925\,
            I => \N__48881\
        );

    \I__11492\ : InMux
    port map (
            O => \N__48924\,
            I => \N__48864\
        );

    \I__11491\ : InMux
    port map (
            O => \N__48923\,
            I => \N__48864\
        );

    \I__11490\ : InMux
    port map (
            O => \N__48922\,
            I => \N__48851\
        );

    \I__11489\ : InMux
    port map (
            O => \N__48921\,
            I => \N__48846\
        );

    \I__11488\ : InMux
    port map (
            O => \N__48920\,
            I => \N__48846\
        );

    \I__11487\ : LocalMux
    port map (
            O => \N__48911\,
            I => \N__48843\
        );

    \I__11486\ : InMux
    port map (
            O => \N__48910\,
            I => \N__48840\
        );

    \I__11485\ : InMux
    port map (
            O => \N__48909\,
            I => \N__48836\
        );

    \I__11484\ : InMux
    port map (
            O => \N__48908\,
            I => \N__48823\
        );

    \I__11483\ : InMux
    port map (
            O => \N__48907\,
            I => \N__48820\
        );

    \I__11482\ : InMux
    port map (
            O => \N__48906\,
            I => \N__48817\
        );

    \I__11481\ : InMux
    port map (
            O => \N__48905\,
            I => \N__48814\
        );

    \I__11480\ : InMux
    port map (
            O => \N__48904\,
            I => \N__48805\
        );

    \I__11479\ : InMux
    port map (
            O => \N__48903\,
            I => \N__48805\
        );

    \I__11478\ : InMux
    port map (
            O => \N__48902\,
            I => \N__48805\
        );

    \I__11477\ : InMux
    port map (
            O => \N__48901\,
            I => \N__48805\
        );

    \I__11476\ : LocalMux
    port map (
            O => \N__48894\,
            I => \N__48802\
        );

    \I__11475\ : InMux
    port map (
            O => \N__48893\,
            I => \N__48795\
        );

    \I__11474\ : InMux
    port map (
            O => \N__48892\,
            I => \N__48795\
        );

    \I__11473\ : InMux
    port map (
            O => \N__48891\,
            I => \N__48795\
        );

    \I__11472\ : InMux
    port map (
            O => \N__48890\,
            I => \N__48788\
        );

    \I__11471\ : InMux
    port map (
            O => \N__48889\,
            I => \N__48788\
        );

    \I__11470\ : InMux
    port map (
            O => \N__48888\,
            I => \N__48788\
        );

    \I__11469\ : InMux
    port map (
            O => \N__48887\,
            I => \N__48779\
        );

    \I__11468\ : InMux
    port map (
            O => \N__48886\,
            I => \N__48779\
        );

    \I__11467\ : InMux
    port map (
            O => \N__48885\,
            I => \N__48779\
        );

    \I__11466\ : InMux
    port map (
            O => \N__48884\,
            I => \N__48779\
        );

    \I__11465\ : LocalMux
    port map (
            O => \N__48881\,
            I => \N__48773\
        );

    \I__11464\ : InMux
    port map (
            O => \N__48880\,
            I => \N__48770\
        );

    \I__11463\ : InMux
    port map (
            O => \N__48879\,
            I => \N__48765\
        );

    \I__11462\ : InMux
    port map (
            O => \N__48878\,
            I => \N__48765\
        );

    \I__11461\ : InMux
    port map (
            O => \N__48877\,
            I => \N__48760\
        );

    \I__11460\ : InMux
    port map (
            O => \N__48876\,
            I => \N__48760\
        );

    \I__11459\ : InMux
    port map (
            O => \N__48875\,
            I => \N__48752\
        );

    \I__11458\ : InMux
    port map (
            O => \N__48874\,
            I => \N__48752\
        );

    \I__11457\ : InMux
    port map (
            O => \N__48873\,
            I => \N__48749\
        );

    \I__11456\ : InMux
    port map (
            O => \N__48872\,
            I => \N__48744\
        );

    \I__11455\ : InMux
    port map (
            O => \N__48871\,
            I => \N__48744\
        );

    \I__11454\ : InMux
    port map (
            O => \N__48870\,
            I => \N__48739\
        );

    \I__11453\ : InMux
    port map (
            O => \N__48869\,
            I => \N__48739\
        );

    \I__11452\ : LocalMux
    port map (
            O => \N__48864\,
            I => \N__48736\
        );

    \I__11451\ : InMux
    port map (
            O => \N__48863\,
            I => \N__48727\
        );

    \I__11450\ : InMux
    port map (
            O => \N__48862\,
            I => \N__48727\
        );

    \I__11449\ : InMux
    port map (
            O => \N__48861\,
            I => \N__48727\
        );

    \I__11448\ : InMux
    port map (
            O => \N__48860\,
            I => \N__48727\
        );

    \I__11447\ : InMux
    port map (
            O => \N__48859\,
            I => \N__48724\
        );

    \I__11446\ : InMux
    port map (
            O => \N__48858\,
            I => \N__48719\
        );

    \I__11445\ : InMux
    port map (
            O => \N__48857\,
            I => \N__48719\
        );

    \I__11444\ : InMux
    port map (
            O => \N__48856\,
            I => \N__48716\
        );

    \I__11443\ : InMux
    port map (
            O => \N__48855\,
            I => \N__48711\
        );

    \I__11442\ : InMux
    port map (
            O => \N__48854\,
            I => \N__48711\
        );

    \I__11441\ : LocalMux
    port map (
            O => \N__48851\,
            I => \N__48702\
        );

    \I__11440\ : LocalMux
    port map (
            O => \N__48846\,
            I => \N__48702\
        );

    \I__11439\ : Span4Mux_v
    port map (
            O => \N__48843\,
            I => \N__48702\
        );

    \I__11438\ : LocalMux
    port map (
            O => \N__48840\,
            I => \N__48702\
        );

    \I__11437\ : InMux
    port map (
            O => \N__48839\,
            I => \N__48699\
        );

    \I__11436\ : LocalMux
    port map (
            O => \N__48836\,
            I => \N__48696\
        );

    \I__11435\ : InMux
    port map (
            O => \N__48835\,
            I => \N__48693\
        );

    \I__11434\ : InMux
    port map (
            O => \N__48834\,
            I => \N__48678\
        );

    \I__11433\ : InMux
    port map (
            O => \N__48833\,
            I => \N__48678\
        );

    \I__11432\ : InMux
    port map (
            O => \N__48832\,
            I => \N__48678\
        );

    \I__11431\ : InMux
    port map (
            O => \N__48831\,
            I => \N__48678\
        );

    \I__11430\ : InMux
    port map (
            O => \N__48830\,
            I => \N__48678\
        );

    \I__11429\ : InMux
    port map (
            O => \N__48829\,
            I => \N__48662\
        );

    \I__11428\ : InMux
    port map (
            O => \N__48828\,
            I => \N__48657\
        );

    \I__11427\ : InMux
    port map (
            O => \N__48827\,
            I => \N__48657\
        );

    \I__11426\ : InMux
    port map (
            O => \N__48826\,
            I => \N__48654\
        );

    \I__11425\ : LocalMux
    port map (
            O => \N__48823\,
            I => \N__48644\
        );

    \I__11424\ : LocalMux
    port map (
            O => \N__48820\,
            I => \N__48644\
        );

    \I__11423\ : LocalMux
    port map (
            O => \N__48817\,
            I => \N__48644\
        );

    \I__11422\ : LocalMux
    port map (
            O => \N__48814\,
            I => \N__48631\
        );

    \I__11421\ : LocalMux
    port map (
            O => \N__48805\,
            I => \N__48631\
        );

    \I__11420\ : Span4Mux_h
    port map (
            O => \N__48802\,
            I => \N__48631\
        );

    \I__11419\ : LocalMux
    port map (
            O => \N__48795\,
            I => \N__48631\
        );

    \I__11418\ : LocalMux
    port map (
            O => \N__48788\,
            I => \N__48631\
        );

    \I__11417\ : LocalMux
    port map (
            O => \N__48779\,
            I => \N__48631\
        );

    \I__11416\ : InMux
    port map (
            O => \N__48778\,
            I => \N__48624\
        );

    \I__11415\ : InMux
    port map (
            O => \N__48777\,
            I => \N__48624\
        );

    \I__11414\ : InMux
    port map (
            O => \N__48776\,
            I => \N__48624\
        );

    \I__11413\ : Span4Mux_h
    port map (
            O => \N__48773\,
            I => \N__48619\
        );

    \I__11412\ : LocalMux
    port map (
            O => \N__48770\,
            I => \N__48619\
        );

    \I__11411\ : LocalMux
    port map (
            O => \N__48765\,
            I => \N__48614\
        );

    \I__11410\ : LocalMux
    port map (
            O => \N__48760\,
            I => \N__48614\
        );

    \I__11409\ : InMux
    port map (
            O => \N__48759\,
            I => \N__48607\
        );

    \I__11408\ : InMux
    port map (
            O => \N__48758\,
            I => \N__48607\
        );

    \I__11407\ : InMux
    port map (
            O => \N__48757\,
            I => \N__48607\
        );

    \I__11406\ : LocalMux
    port map (
            O => \N__48752\,
            I => \N__48590\
        );

    \I__11405\ : LocalMux
    port map (
            O => \N__48749\,
            I => \N__48590\
        );

    \I__11404\ : LocalMux
    port map (
            O => \N__48744\,
            I => \N__48590\
        );

    \I__11403\ : LocalMux
    port map (
            O => \N__48739\,
            I => \N__48590\
        );

    \I__11402\ : Span4Mux_v
    port map (
            O => \N__48736\,
            I => \N__48590\
        );

    \I__11401\ : LocalMux
    port map (
            O => \N__48727\,
            I => \N__48590\
        );

    \I__11400\ : LocalMux
    port map (
            O => \N__48724\,
            I => \N__48590\
        );

    \I__11399\ : LocalMux
    port map (
            O => \N__48719\,
            I => \N__48590\
        );

    \I__11398\ : LocalMux
    port map (
            O => \N__48716\,
            I => \N__48583\
        );

    \I__11397\ : LocalMux
    port map (
            O => \N__48711\,
            I => \N__48583\
        );

    \I__11396\ : Span4Mux_v
    port map (
            O => \N__48702\,
            I => \N__48583\
        );

    \I__11395\ : LocalMux
    port map (
            O => \N__48699\,
            I => \N__48580\
        );

    \I__11394\ : Span4Mux_v
    port map (
            O => \N__48696\,
            I => \N__48575\
        );

    \I__11393\ : LocalMux
    port map (
            O => \N__48693\,
            I => \N__48575\
        );

    \I__11392\ : InMux
    port map (
            O => \N__48692\,
            I => \N__48568\
        );

    \I__11391\ : InMux
    port map (
            O => \N__48691\,
            I => \N__48568\
        );

    \I__11390\ : InMux
    port map (
            O => \N__48690\,
            I => \N__48568\
        );

    \I__11389\ : InMux
    port map (
            O => \N__48689\,
            I => \N__48565\
        );

    \I__11388\ : LocalMux
    port map (
            O => \N__48678\,
            I => \N__48562\
        );

    \I__11387\ : InMux
    port map (
            O => \N__48677\,
            I => \N__48549\
        );

    \I__11386\ : InMux
    port map (
            O => \N__48676\,
            I => \N__48549\
        );

    \I__11385\ : InMux
    port map (
            O => \N__48675\,
            I => \N__48549\
        );

    \I__11384\ : InMux
    port map (
            O => \N__48674\,
            I => \N__48549\
        );

    \I__11383\ : InMux
    port map (
            O => \N__48673\,
            I => \N__48549\
        );

    \I__11382\ : InMux
    port map (
            O => \N__48672\,
            I => \N__48549\
        );

    \I__11381\ : InMux
    port map (
            O => \N__48671\,
            I => \N__48540\
        );

    \I__11380\ : InMux
    port map (
            O => \N__48670\,
            I => \N__48540\
        );

    \I__11379\ : InMux
    port map (
            O => \N__48669\,
            I => \N__48540\
        );

    \I__11378\ : InMux
    port map (
            O => \N__48668\,
            I => \N__48540\
        );

    \I__11377\ : InMux
    port map (
            O => \N__48667\,
            I => \N__48533\
        );

    \I__11376\ : InMux
    port map (
            O => \N__48666\,
            I => \N__48533\
        );

    \I__11375\ : InMux
    port map (
            O => \N__48665\,
            I => \N__48533\
        );

    \I__11374\ : LocalMux
    port map (
            O => \N__48662\,
            I => \N__48526\
        );

    \I__11373\ : LocalMux
    port map (
            O => \N__48657\,
            I => \N__48526\
        );

    \I__11372\ : LocalMux
    port map (
            O => \N__48654\,
            I => \N__48526\
        );

    \I__11371\ : InMux
    port map (
            O => \N__48653\,
            I => \N__48519\
        );

    \I__11370\ : InMux
    port map (
            O => \N__48652\,
            I => \N__48519\
        );

    \I__11369\ : InMux
    port map (
            O => \N__48651\,
            I => \N__48519\
        );

    \I__11368\ : Span4Mux_v
    port map (
            O => \N__48644\,
            I => \N__48512\
        );

    \I__11367\ : Span4Mux_v
    port map (
            O => \N__48631\,
            I => \N__48512\
        );

    \I__11366\ : LocalMux
    port map (
            O => \N__48624\,
            I => \N__48512\
        );

    \I__11365\ : Span4Mux_h
    port map (
            O => \N__48619\,
            I => \N__48507\
        );

    \I__11364\ : Span4Mux_h
    port map (
            O => \N__48614\,
            I => \N__48507\
        );

    \I__11363\ : LocalMux
    port map (
            O => \N__48607\,
            I => \N__48500\
        );

    \I__11362\ : Span4Mux_v
    port map (
            O => \N__48590\,
            I => \N__48500\
        );

    \I__11361\ : Span4Mux_h
    port map (
            O => \N__48583\,
            I => \N__48500\
        );

    \I__11360\ : Span4Mux_v
    port map (
            O => \N__48580\,
            I => \N__48495\
        );

    \I__11359\ : Span4Mux_h
    port map (
            O => \N__48575\,
            I => \N__48495\
        );

    \I__11358\ : LocalMux
    port map (
            O => \N__48568\,
            I => \N__48488\
        );

    \I__11357\ : LocalMux
    port map (
            O => \N__48565\,
            I => \N__48488\
        );

    \I__11356\ : Span12Mux_s8_h
    port map (
            O => \N__48562\,
            I => \N__48488\
        );

    \I__11355\ : LocalMux
    port map (
            O => \N__48549\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11354\ : LocalMux
    port map (
            O => \N__48540\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11353\ : LocalMux
    port map (
            O => \N__48533\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11352\ : Odrv4
    port map (
            O => \N__48526\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11351\ : LocalMux
    port map (
            O => \N__48519\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11350\ : Odrv4
    port map (
            O => \N__48512\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11349\ : Odrv4
    port map (
            O => \N__48507\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11348\ : Odrv4
    port map (
            O => \N__48500\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11347\ : Odrv4
    port map (
            O => \N__48495\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11346\ : Odrv12
    port map (
            O => \N__48488\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11345\ : InMux
    port map (
            O => \N__48467\,
            I => \N__48464\
        );

    \I__11344\ : LocalMux
    port map (
            O => \N__48464\,
            I => \N__48459\
        );

    \I__11343\ : InMux
    port map (
            O => \N__48463\,
            I => \N__48456\
        );

    \I__11342\ : InMux
    port map (
            O => \N__48462\,
            I => \N__48453\
        );

    \I__11341\ : Span4Mux_v
    port map (
            O => \N__48459\,
            I => \N__48450\
        );

    \I__11340\ : LocalMux
    port map (
            O => \N__48456\,
            I => \N__48447\
        );

    \I__11339\ : LocalMux
    port map (
            O => \N__48453\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27\
        );

    \I__11338\ : Odrv4
    port map (
            O => \N__48450\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27\
        );

    \I__11337\ : Odrv4
    port map (
            O => \N__48447\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27\
        );

    \I__11336\ : CascadeMux
    port map (
            O => \N__48440\,
            I => \N__48432\
        );

    \I__11335\ : InMux
    port map (
            O => \N__48439\,
            I => \N__48428\
        );

    \I__11334\ : InMux
    port map (
            O => \N__48438\,
            I => \N__48425\
        );

    \I__11333\ : InMux
    port map (
            O => \N__48437\,
            I => \N__48422\
        );

    \I__11332\ : InMux
    port map (
            O => \N__48436\,
            I => \N__48419\
        );

    \I__11331\ : InMux
    port map (
            O => \N__48435\,
            I => \N__48397\
        );

    \I__11330\ : InMux
    port map (
            O => \N__48432\,
            I => \N__48397\
        );

    \I__11329\ : InMux
    port map (
            O => \N__48431\,
            I => \N__48397\
        );

    \I__11328\ : LocalMux
    port map (
            O => \N__48428\,
            I => \N__48388\
        );

    \I__11327\ : LocalMux
    port map (
            O => \N__48425\,
            I => \N__48388\
        );

    \I__11326\ : LocalMux
    port map (
            O => \N__48422\,
            I => \N__48388\
        );

    \I__11325\ : LocalMux
    port map (
            O => \N__48419\,
            I => \N__48388\
        );

    \I__11324\ : InMux
    port map (
            O => \N__48418\,
            I => \N__48381\
        );

    \I__11323\ : InMux
    port map (
            O => \N__48417\,
            I => \N__48381\
        );

    \I__11322\ : InMux
    port map (
            O => \N__48416\,
            I => \N__48381\
        );

    \I__11321\ : InMux
    port map (
            O => \N__48415\,
            I => \N__48372\
        );

    \I__11320\ : InMux
    port map (
            O => \N__48414\,
            I => \N__48372\
        );

    \I__11319\ : InMux
    port map (
            O => \N__48413\,
            I => \N__48372\
        );

    \I__11318\ : InMux
    port map (
            O => \N__48412\,
            I => \N__48372\
        );

    \I__11317\ : InMux
    port map (
            O => \N__48411\,
            I => \N__48368\
        );

    \I__11316\ : InMux
    port map (
            O => \N__48410\,
            I => \N__48363\
        );

    \I__11315\ : InMux
    port map (
            O => \N__48409\,
            I => \N__48363\
        );

    \I__11314\ : InMux
    port map (
            O => \N__48408\,
            I => \N__48360\
        );

    \I__11313\ : InMux
    port map (
            O => \N__48407\,
            I => \N__48355\
        );

    \I__11312\ : InMux
    port map (
            O => \N__48406\,
            I => \N__48355\
        );

    \I__11311\ : InMux
    port map (
            O => \N__48405\,
            I => \N__48352\
        );

    \I__11310\ : InMux
    port map (
            O => \N__48404\,
            I => \N__48349\
        );

    \I__11309\ : LocalMux
    port map (
            O => \N__48397\,
            I => \N__48345\
        );

    \I__11308\ : Span12Mux_s6_v
    port map (
            O => \N__48388\,
            I => \N__48326\
        );

    \I__11307\ : LocalMux
    port map (
            O => \N__48381\,
            I => \N__48326\
        );

    \I__11306\ : LocalMux
    port map (
            O => \N__48372\,
            I => \N__48326\
        );

    \I__11305\ : InMux
    port map (
            O => \N__48371\,
            I => \N__48323\
        );

    \I__11304\ : LocalMux
    port map (
            O => \N__48368\,
            I => \N__48312\
        );

    \I__11303\ : LocalMux
    port map (
            O => \N__48363\,
            I => \N__48312\
        );

    \I__11302\ : LocalMux
    port map (
            O => \N__48360\,
            I => \N__48312\
        );

    \I__11301\ : LocalMux
    port map (
            O => \N__48355\,
            I => \N__48312\
        );

    \I__11300\ : LocalMux
    port map (
            O => \N__48352\,
            I => \N__48312\
        );

    \I__11299\ : LocalMux
    port map (
            O => \N__48349\,
            I => \N__48309\
        );

    \I__11298\ : InMux
    port map (
            O => \N__48348\,
            I => \N__48306\
        );

    \I__11297\ : Span4Mux_h
    port map (
            O => \N__48345\,
            I => \N__48296\
        );

    \I__11296\ : CascadeMux
    port map (
            O => \N__48344\,
            I => \N__48292\
        );

    \I__11295\ : CascadeMux
    port map (
            O => \N__48343\,
            I => \N__48288\
        );

    \I__11294\ : CascadeMux
    port map (
            O => \N__48342\,
            I => \N__48284\
        );

    \I__11293\ : CascadeMux
    port map (
            O => \N__48341\,
            I => \N__48280\
        );

    \I__11292\ : CascadeMux
    port map (
            O => \N__48340\,
            I => \N__48276\
        );

    \I__11291\ : CascadeMux
    port map (
            O => \N__48339\,
            I => \N__48272\
        );

    \I__11290\ : CascadeMux
    port map (
            O => \N__48338\,
            I => \N__48268\
        );

    \I__11289\ : CascadeMux
    port map (
            O => \N__48337\,
            I => \N__48264\
        );

    \I__11288\ : CascadeMux
    port map (
            O => \N__48336\,
            I => \N__48260\
        );

    \I__11287\ : CascadeMux
    port map (
            O => \N__48335\,
            I => \N__48256\
        );

    \I__11286\ : CascadeMux
    port map (
            O => \N__48334\,
            I => \N__48252\
        );

    \I__11285\ : InMux
    port map (
            O => \N__48333\,
            I => \N__48245\
        );

    \I__11284\ : Span12Mux_v
    port map (
            O => \N__48326\,
            I => \N__48238\
        );

    \I__11283\ : LocalMux
    port map (
            O => \N__48323\,
            I => \N__48238\
        );

    \I__11282\ : Span12Mux_s11_v
    port map (
            O => \N__48312\,
            I => \N__48238\
        );

    \I__11281\ : Span4Mux_s1_h
    port map (
            O => \N__48309\,
            I => \N__48235\
        );

    \I__11280\ : LocalMux
    port map (
            O => \N__48306\,
            I => \N__48232\
        );

    \I__11279\ : InMux
    port map (
            O => \N__48305\,
            I => \N__48225\
        );

    \I__11278\ : InMux
    port map (
            O => \N__48304\,
            I => \N__48225\
        );

    \I__11277\ : InMux
    port map (
            O => \N__48303\,
            I => \N__48225\
        );

    \I__11276\ : InMux
    port map (
            O => \N__48302\,
            I => \N__48216\
        );

    \I__11275\ : InMux
    port map (
            O => \N__48301\,
            I => \N__48216\
        );

    \I__11274\ : InMux
    port map (
            O => \N__48300\,
            I => \N__48216\
        );

    \I__11273\ : InMux
    port map (
            O => \N__48299\,
            I => \N__48216\
        );

    \I__11272\ : Span4Mux_h
    port map (
            O => \N__48296\,
            I => \N__48213\
        );

    \I__11271\ : InMux
    port map (
            O => \N__48295\,
            I => \N__48198\
        );

    \I__11270\ : InMux
    port map (
            O => \N__48292\,
            I => \N__48198\
        );

    \I__11269\ : InMux
    port map (
            O => \N__48291\,
            I => \N__48198\
        );

    \I__11268\ : InMux
    port map (
            O => \N__48288\,
            I => \N__48198\
        );

    \I__11267\ : InMux
    port map (
            O => \N__48287\,
            I => \N__48198\
        );

    \I__11266\ : InMux
    port map (
            O => \N__48284\,
            I => \N__48198\
        );

    \I__11265\ : InMux
    port map (
            O => \N__48283\,
            I => \N__48198\
        );

    \I__11264\ : InMux
    port map (
            O => \N__48280\,
            I => \N__48181\
        );

    \I__11263\ : InMux
    port map (
            O => \N__48279\,
            I => \N__48181\
        );

    \I__11262\ : InMux
    port map (
            O => \N__48276\,
            I => \N__48181\
        );

    \I__11261\ : InMux
    port map (
            O => \N__48275\,
            I => \N__48181\
        );

    \I__11260\ : InMux
    port map (
            O => \N__48272\,
            I => \N__48181\
        );

    \I__11259\ : InMux
    port map (
            O => \N__48271\,
            I => \N__48181\
        );

    \I__11258\ : InMux
    port map (
            O => \N__48268\,
            I => \N__48181\
        );

    \I__11257\ : InMux
    port map (
            O => \N__48267\,
            I => \N__48181\
        );

    \I__11256\ : InMux
    port map (
            O => \N__48264\,
            I => \N__48164\
        );

    \I__11255\ : InMux
    port map (
            O => \N__48263\,
            I => \N__48164\
        );

    \I__11254\ : InMux
    port map (
            O => \N__48260\,
            I => \N__48164\
        );

    \I__11253\ : InMux
    port map (
            O => \N__48259\,
            I => \N__48164\
        );

    \I__11252\ : InMux
    port map (
            O => \N__48256\,
            I => \N__48164\
        );

    \I__11251\ : InMux
    port map (
            O => \N__48255\,
            I => \N__48164\
        );

    \I__11250\ : InMux
    port map (
            O => \N__48252\,
            I => \N__48164\
        );

    \I__11249\ : InMux
    port map (
            O => \N__48251\,
            I => \N__48164\
        );

    \I__11248\ : CascadeMux
    port map (
            O => \N__48250\,
            I => \N__48160\
        );

    \I__11247\ : CascadeMux
    port map (
            O => \N__48249\,
            I => \N__48156\
        );

    \I__11246\ : CascadeMux
    port map (
            O => \N__48248\,
            I => \N__48152\
        );

    \I__11245\ : LocalMux
    port map (
            O => \N__48245\,
            I => \N__48147\
        );

    \I__11244\ : Span12Mux_h
    port map (
            O => \N__48238\,
            I => \N__48144\
        );

    \I__11243\ : Span4Mux_v
    port map (
            O => \N__48235\,
            I => \N__48139\
        );

    \I__11242\ : Span4Mux_s1_h
    port map (
            O => \N__48232\,
            I => \N__48139\
        );

    \I__11241\ : LocalMux
    port map (
            O => \N__48225\,
            I => \N__48134\
        );

    \I__11240\ : LocalMux
    port map (
            O => \N__48216\,
            I => \N__48134\
        );

    \I__11239\ : Sp12to4
    port map (
            O => \N__48213\,
            I => \N__48129\
        );

    \I__11238\ : LocalMux
    port map (
            O => \N__48198\,
            I => \N__48129\
        );

    \I__11237\ : LocalMux
    port map (
            O => \N__48181\,
            I => \N__48126\
        );

    \I__11236\ : LocalMux
    port map (
            O => \N__48164\,
            I => \N__48123\
        );

    \I__11235\ : InMux
    port map (
            O => \N__48163\,
            I => \N__48108\
        );

    \I__11234\ : InMux
    port map (
            O => \N__48160\,
            I => \N__48108\
        );

    \I__11233\ : InMux
    port map (
            O => \N__48159\,
            I => \N__48108\
        );

    \I__11232\ : InMux
    port map (
            O => \N__48156\,
            I => \N__48108\
        );

    \I__11231\ : InMux
    port map (
            O => \N__48155\,
            I => \N__48108\
        );

    \I__11230\ : InMux
    port map (
            O => \N__48152\,
            I => \N__48108\
        );

    \I__11229\ : InMux
    port map (
            O => \N__48151\,
            I => \N__48108\
        );

    \I__11228\ : InMux
    port map (
            O => \N__48150\,
            I => \N__48105\
        );

    \I__11227\ : Span4Mux_v
    port map (
            O => \N__48147\,
            I => \N__48102\
        );

    \I__11226\ : Span12Mux_h
    port map (
            O => \N__48144\,
            I => \N__48095\
        );

    \I__11225\ : Sp12to4
    port map (
            O => \N__48139\,
            I => \N__48095\
        );

    \I__11224\ : Span12Mux_s1_h
    port map (
            O => \N__48134\,
            I => \N__48095\
        );

    \I__11223\ : Span12Mux_s9_v
    port map (
            O => \N__48129\,
            I => \N__48084\
        );

    \I__11222\ : Sp12to4
    port map (
            O => \N__48126\,
            I => \N__48084\
        );

    \I__11221\ : Span12Mux_s8_h
    port map (
            O => \N__48123\,
            I => \N__48084\
        );

    \I__11220\ : LocalMux
    port map (
            O => \N__48108\,
            I => \N__48084\
        );

    \I__11219\ : LocalMux
    port map (
            O => \N__48105\,
            I => \N__48084\
        );

    \I__11218\ : Span4Mux_v
    port map (
            O => \N__48102\,
            I => \N__48081\
        );

    \I__11217\ : Span12Mux_v
    port map (
            O => \N__48095\,
            I => \N__48078\
        );

    \I__11216\ : Span12Mux_v
    port map (
            O => \N__48084\,
            I => \N__48075\
        );

    \I__11215\ : Span4Mux_h
    port map (
            O => \N__48081\,
            I => \N__48072\
        );

    \I__11214\ : Odrv12
    port map (
            O => \N__48078\,
            I => \CONSTANT_ONE_NET\
        );

    \I__11213\ : Odrv12
    port map (
            O => \N__48075\,
            I => \CONSTANT_ONE_NET\
        );

    \I__11212\ : Odrv4
    port map (
            O => \N__48072\,
            I => \CONSTANT_ONE_NET\
        );

    \I__11211\ : CascadeMux
    port map (
            O => \N__48065\,
            I => \N__48060\
        );

    \I__11210\ : InMux
    port map (
            O => \N__48064\,
            I => \N__48057\
        );

    \I__11209\ : InMux
    port map (
            O => \N__48063\,
            I => \N__48054\
        );

    \I__11208\ : InMux
    port map (
            O => \N__48060\,
            I => \N__48051\
        );

    \I__11207\ : LocalMux
    port map (
            O => \N__48057\,
            I => \N__48048\
        );

    \I__11206\ : LocalMux
    port map (
            O => \N__48054\,
            I => \N__48044\
        );

    \I__11205\ : LocalMux
    port map (
            O => \N__48051\,
            I => \N__48041\
        );

    \I__11204\ : Span4Mux_h
    port map (
            O => \N__48048\,
            I => \N__48038\
        );

    \I__11203\ : InMux
    port map (
            O => \N__48047\,
            I => \N__48035\
        );

    \I__11202\ : Span12Mux_h
    port map (
            O => \N__48044\,
            I => \N__48032\
        );

    \I__11201\ : Span4Mux_v
    port map (
            O => \N__48041\,
            I => \N__48027\
        );

    \I__11200\ : Span4Mux_h
    port map (
            O => \N__48038\,
            I => \N__48027\
        );

    \I__11199\ : LocalMux
    port map (
            O => \N__48035\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__11198\ : Odrv12
    port map (
            O => \N__48032\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__11197\ : Odrv4
    port map (
            O => \N__48027\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__11196\ : InMux
    port map (
            O => \N__48020\,
            I => \N__48017\
        );

    \I__11195\ : LocalMux
    port map (
            O => \N__48017\,
            I => \N__48014\
        );

    \I__11194\ : Span4Mux_h
    port map (
            O => \N__48014\,
            I => \N__48010\
        );

    \I__11193\ : InMux
    port map (
            O => \N__48013\,
            I => \N__48007\
        );

    \I__11192\ : Span4Mux_h
    port map (
            O => \N__48010\,
            I => \N__48004\
        );

    \I__11191\ : LocalMux
    port map (
            O => \N__48007\,
            I => \N__48001\
        );

    \I__11190\ : Span4Mux_v
    port map (
            O => \N__48004\,
            I => \N__47997\
        );

    \I__11189\ : Span4Mux_h
    port map (
            O => \N__48001\,
            I => \N__47993\
        );

    \I__11188\ : InMux
    port map (
            O => \N__48000\,
            I => \N__47990\
        );

    \I__11187\ : Span4Mux_v
    port map (
            O => \N__47997\,
            I => \N__47987\
        );

    \I__11186\ : InMux
    port map (
            O => \N__47996\,
            I => \N__47984\
        );

    \I__11185\ : Span4Mux_h
    port map (
            O => \N__47993\,
            I => \N__47981\
        );

    \I__11184\ : LocalMux
    port map (
            O => \N__47990\,
            I => \N__47978\
        );

    \I__11183\ : Odrv4
    port map (
            O => \N__47987\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__11182\ : LocalMux
    port map (
            O => \N__47984\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__11181\ : Odrv4
    port map (
            O => \N__47981\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__11180\ : Odrv12
    port map (
            O => \N__47978\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__11179\ : InMux
    port map (
            O => \N__47969\,
            I => \N__47966\
        );

    \I__11178\ : LocalMux
    port map (
            O => \N__47966\,
            I => \N__47963\
        );

    \I__11177\ : Span4Mux_v
    port map (
            O => \N__47963\,
            I => \N__47959\
        );

    \I__11176\ : InMux
    port map (
            O => \N__47962\,
            I => \N__47956\
        );

    \I__11175\ : Span4Mux_h
    port map (
            O => \N__47959\,
            I => \N__47953\
        );

    \I__11174\ : LocalMux
    port map (
            O => \N__47956\,
            I => \N__47950\
        );

    \I__11173\ : Odrv4
    port map (
            O => \N__47953\,
            I => \phase_controller_inst1.state_RNIE87FZ0Z_2\
        );

    \I__11172\ : Odrv12
    port map (
            O => \N__47950\,
            I => \phase_controller_inst1.state_RNIE87FZ0Z_2\
        );

    \I__11171\ : InMux
    port map (
            O => \N__47945\,
            I => \N__47940\
        );

    \I__11170\ : InMux
    port map (
            O => \N__47944\,
            I => \N__47937\
        );

    \I__11169\ : InMux
    port map (
            O => \N__47943\,
            I => \N__47934\
        );

    \I__11168\ : LocalMux
    port map (
            O => \N__47940\,
            I => \N__47931\
        );

    \I__11167\ : LocalMux
    port map (
            O => \N__47937\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18\
        );

    \I__11166\ : LocalMux
    port map (
            O => \N__47934\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18\
        );

    \I__11165\ : Odrv4
    port map (
            O => \N__47931\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18\
        );

    \I__11164\ : InMux
    port map (
            O => \N__47924\,
            I => \N__47919\
        );

    \I__11163\ : InMux
    port map (
            O => \N__47923\,
            I => \N__47916\
        );

    \I__11162\ : InMux
    port map (
            O => \N__47922\,
            I => \N__47913\
        );

    \I__11161\ : LocalMux
    port map (
            O => \N__47919\,
            I => \N__47908\
        );

    \I__11160\ : LocalMux
    port map (
            O => \N__47916\,
            I => \N__47908\
        );

    \I__11159\ : LocalMux
    port map (
            O => \N__47913\,
            I => \N__47904\
        );

    \I__11158\ : Span4Mux_h
    port map (
            O => \N__47908\,
            I => \N__47901\
        );

    \I__11157\ : InMux
    port map (
            O => \N__47907\,
            I => \N__47898\
        );

    \I__11156\ : Odrv12
    port map (
            O => \N__47904\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__11155\ : Odrv4
    port map (
            O => \N__47901\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__11154\ : LocalMux
    port map (
            O => \N__47898\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__11153\ : InMux
    port map (
            O => \N__47891\,
            I => \N__47885\
        );

    \I__11152\ : InMux
    port map (
            O => \N__47890\,
            I => \N__47885\
        );

    \I__11151\ : LocalMux
    port map (
            O => \N__47885\,
            I => \N__47882\
        );

    \I__11150\ : Span4Mux_h
    port map (
            O => \N__47882\,
            I => \N__47879\
        );

    \I__11149\ : Span4Mux_h
    port map (
            O => \N__47879\,
            I => \N__47876\
        );

    \I__11148\ : Odrv4
    port map (
            O => \N__47876\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\
        );

    \I__11147\ : CEMux
    port map (
            O => \N__47873\,
            I => \N__47831\
        );

    \I__11146\ : CEMux
    port map (
            O => \N__47872\,
            I => \N__47831\
        );

    \I__11145\ : CEMux
    port map (
            O => \N__47871\,
            I => \N__47831\
        );

    \I__11144\ : CEMux
    port map (
            O => \N__47870\,
            I => \N__47831\
        );

    \I__11143\ : CEMux
    port map (
            O => \N__47869\,
            I => \N__47831\
        );

    \I__11142\ : CEMux
    port map (
            O => \N__47868\,
            I => \N__47831\
        );

    \I__11141\ : CEMux
    port map (
            O => \N__47867\,
            I => \N__47831\
        );

    \I__11140\ : CEMux
    port map (
            O => \N__47866\,
            I => \N__47831\
        );

    \I__11139\ : CEMux
    port map (
            O => \N__47865\,
            I => \N__47831\
        );

    \I__11138\ : CEMux
    port map (
            O => \N__47864\,
            I => \N__47831\
        );

    \I__11137\ : CEMux
    port map (
            O => \N__47863\,
            I => \N__47831\
        );

    \I__11136\ : CEMux
    port map (
            O => \N__47862\,
            I => \N__47831\
        );

    \I__11135\ : CEMux
    port map (
            O => \N__47861\,
            I => \N__47831\
        );

    \I__11134\ : CEMux
    port map (
            O => \N__47860\,
            I => \N__47831\
        );

    \I__11133\ : GlobalMux
    port map (
            O => \N__47831\,
            I => \N__47828\
        );

    \I__11132\ : gio2CtrlBuf
    port map (
            O => \N__47828\,
            I => \phase_controller_inst2.stoper_hc.un1_start_g\
        );

    \I__11131\ : InMux
    port map (
            O => \N__47825\,
            I => \N__47820\
        );

    \I__11130\ : InMux
    port map (
            O => \N__47824\,
            I => \N__47817\
        );

    \I__11129\ : InMux
    port map (
            O => \N__47823\,
            I => \N__47814\
        );

    \I__11128\ : LocalMux
    port map (
            O => \N__47820\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16\
        );

    \I__11127\ : LocalMux
    port map (
            O => \N__47817\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16\
        );

    \I__11126\ : LocalMux
    port map (
            O => \N__47814\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16\
        );

    \I__11125\ : InMux
    port map (
            O => \N__47807\,
            I => \N__47804\
        );

    \I__11124\ : LocalMux
    port map (
            O => \N__47804\,
            I => \N__47799\
        );

    \I__11123\ : InMux
    port map (
            O => \N__47803\,
            I => \N__47796\
        );

    \I__11122\ : InMux
    port map (
            O => \N__47802\,
            I => \N__47793\
        );

    \I__11121\ : Span4Mux_v
    port map (
            O => \N__47799\,
            I => \N__47789\
        );

    \I__11120\ : LocalMux
    port map (
            O => \N__47796\,
            I => \N__47784\
        );

    \I__11119\ : LocalMux
    port map (
            O => \N__47793\,
            I => \N__47784\
        );

    \I__11118\ : CascadeMux
    port map (
            O => \N__47792\,
            I => \N__47781\
        );

    \I__11117\ : Span4Mux_h
    port map (
            O => \N__47789\,
            I => \N__47778\
        );

    \I__11116\ : Span4Mux_v
    port map (
            O => \N__47784\,
            I => \N__47775\
        );

    \I__11115\ : InMux
    port map (
            O => \N__47781\,
            I => \N__47772\
        );

    \I__11114\ : Odrv4
    port map (
            O => \N__47778\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__11113\ : Odrv4
    port map (
            O => \N__47775\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__11112\ : LocalMux
    port map (
            O => \N__47772\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__11111\ : InMux
    port map (
            O => \N__47765\,
            I => \N__47759\
        );

    \I__11110\ : InMux
    port map (
            O => \N__47764\,
            I => \N__47759\
        );

    \I__11109\ : LocalMux
    port map (
            O => \N__47759\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\
        );

    \I__11108\ : InMux
    port map (
            O => \N__47756\,
            I => \N__47753\
        );

    \I__11107\ : LocalMux
    port map (
            O => \N__47753\,
            I => \N__47750\
        );

    \I__11106\ : Span4Mux_h
    port map (
            O => \N__47750\,
            I => \N__47745\
        );

    \I__11105\ : InMux
    port map (
            O => \N__47749\,
            I => \N__47742\
        );

    \I__11104\ : InMux
    port map (
            O => \N__47748\,
            I => \N__47739\
        );

    \I__11103\ : Span4Mux_h
    port map (
            O => \N__47745\,
            I => \N__47734\
        );

    \I__11102\ : LocalMux
    port map (
            O => \N__47742\,
            I => \N__47734\
        );

    \I__11101\ : LocalMux
    port map (
            O => \N__47739\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22\
        );

    \I__11100\ : Odrv4
    port map (
            O => \N__47734\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22\
        );

    \I__11099\ : InMux
    port map (
            O => \N__47729\,
            I => \N__47724\
        );

    \I__11098\ : InMux
    port map (
            O => \N__47728\,
            I => \N__47721\
        );

    \I__11097\ : InMux
    port map (
            O => \N__47727\,
            I => \N__47717\
        );

    \I__11096\ : LocalMux
    port map (
            O => \N__47724\,
            I => \N__47714\
        );

    \I__11095\ : LocalMux
    port map (
            O => \N__47721\,
            I => \N__47711\
        );

    \I__11094\ : InMux
    port map (
            O => \N__47720\,
            I => \N__47708\
        );

    \I__11093\ : LocalMux
    port map (
            O => \N__47717\,
            I => \N__47705\
        );

    \I__11092\ : Span4Mux_h
    port map (
            O => \N__47714\,
            I => \N__47700\
        );

    \I__11091\ : Span4Mux_v
    port map (
            O => \N__47711\,
            I => \N__47700\
        );

    \I__11090\ : LocalMux
    port map (
            O => \N__47708\,
            I => \N__47697\
        );

    \I__11089\ : Odrv12
    port map (
            O => \N__47705\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__11088\ : Odrv4
    port map (
            O => \N__47700\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__11087\ : Odrv4
    port map (
            O => \N__47697\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__11086\ : CascadeMux
    port map (
            O => \N__47690\,
            I => \N__47687\
        );

    \I__11085\ : InMux
    port map (
            O => \N__47687\,
            I => \N__47684\
        );

    \I__11084\ : LocalMux
    port map (
            O => \N__47684\,
            I => \N__47681\
        );

    \I__11083\ : Span4Mux_h
    port map (
            O => \N__47681\,
            I => \N__47678\
        );

    \I__11082\ : Odrv4
    port map (
            O => \N__47678\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt22\
        );

    \I__11081\ : InMux
    port map (
            O => \N__47675\,
            I => \N__47672\
        );

    \I__11080\ : LocalMux
    port map (
            O => \N__47672\,
            I => \N__47669\
        );

    \I__11079\ : Span12Mux_h
    port map (
            O => \N__47669\,
            I => \N__47665\
        );

    \I__11078\ : InMux
    port map (
            O => \N__47668\,
            I => \N__47662\
        );

    \I__11077\ : Odrv12
    port map (
            O => \N__47665\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23\
        );

    \I__11076\ : LocalMux
    port map (
            O => \N__47662\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23\
        );

    \I__11075\ : InMux
    port map (
            O => \N__47657\,
            I => \N__47650\
        );

    \I__11074\ : InMux
    port map (
            O => \N__47656\,
            I => \N__47650\
        );

    \I__11073\ : InMux
    port map (
            O => \N__47655\,
            I => \N__47647\
        );

    \I__11072\ : LocalMux
    port map (
            O => \N__47650\,
            I => \N__47644\
        );

    \I__11071\ : LocalMux
    port map (
            O => \N__47647\,
            I => \N__47640\
        );

    \I__11070\ : Span4Mux_v
    port map (
            O => \N__47644\,
            I => \N__47637\
        );

    \I__11069\ : InMux
    port map (
            O => \N__47643\,
            I => \N__47634\
        );

    \I__11068\ : Span4Mux_v
    port map (
            O => \N__47640\,
            I => \N__47629\
        );

    \I__11067\ : Span4Mux_h
    port map (
            O => \N__47637\,
            I => \N__47629\
        );

    \I__11066\ : LocalMux
    port map (
            O => \N__47634\,
            I => \N__47626\
        );

    \I__11065\ : Odrv4
    port map (
            O => \N__47629\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__11064\ : Odrv4
    port map (
            O => \N__47626\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__11063\ : CascadeMux
    port map (
            O => \N__47621\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23_cascade_\
        );

    \I__11062\ : InMux
    port map (
            O => \N__47618\,
            I => \N__47612\
        );

    \I__11061\ : InMux
    port map (
            O => \N__47617\,
            I => \N__47612\
        );

    \I__11060\ : LocalMux
    port map (
            O => \N__47612\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_22\
        );

    \I__11059\ : InMux
    port map (
            O => \N__47609\,
            I => \N__47603\
        );

    \I__11058\ : InMux
    port map (
            O => \N__47608\,
            I => \N__47603\
        );

    \I__11057\ : LocalMux
    port map (
            O => \N__47603\,
            I => \N__47599\
        );

    \I__11056\ : InMux
    port map (
            O => \N__47602\,
            I => \N__47596\
        );

    \I__11055\ : Span4Mux_h
    port map (
            O => \N__47599\,
            I => \N__47593\
        );

    \I__11054\ : LocalMux
    port map (
            O => \N__47596\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__11053\ : Odrv4
    port map (
            O => \N__47593\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__11052\ : CascadeMux
    port map (
            O => \N__47588\,
            I => \N__47584\
        );

    \I__11051\ : CascadeMux
    port map (
            O => \N__47587\,
            I => \N__47581\
        );

    \I__11050\ : InMux
    port map (
            O => \N__47584\,
            I => \N__47576\
        );

    \I__11049\ : InMux
    port map (
            O => \N__47581\,
            I => \N__47576\
        );

    \I__11048\ : LocalMux
    port map (
            O => \N__47576\,
            I => \N__47572\
        );

    \I__11047\ : InMux
    port map (
            O => \N__47575\,
            I => \N__47569\
        );

    \I__11046\ : Span4Mux_h
    port map (
            O => \N__47572\,
            I => \N__47566\
        );

    \I__11045\ : LocalMux
    port map (
            O => \N__47569\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__11044\ : Odrv4
    port map (
            O => \N__47566\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__11043\ : InMux
    port map (
            O => \N__47561\,
            I => \N__47555\
        );

    \I__11042\ : InMux
    port map (
            O => \N__47560\,
            I => \N__47555\
        );

    \I__11041\ : LocalMux
    port map (
            O => \N__47555\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_23\
        );

    \I__11040\ : InMux
    port map (
            O => \N__47552\,
            I => \N__47549\
        );

    \I__11039\ : LocalMux
    port map (
            O => \N__47549\,
            I => \N__47546\
        );

    \I__11038\ : Odrv12
    port map (
            O => \N__47546\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22\
        );

    \I__11037\ : InMux
    port map (
            O => \N__47543\,
            I => \N__47540\
        );

    \I__11036\ : LocalMux
    port map (
            O => \N__47540\,
            I => \N__47537\
        );

    \I__11035\ : Span4Mux_h
    port map (
            O => \N__47537\,
            I => \N__47534\
        );

    \I__11034\ : Span4Mux_h
    port map (
            O => \N__47534\,
            I => \N__47530\
        );

    \I__11033\ : InMux
    port map (
            O => \N__47533\,
            I => \N__47527\
        );

    \I__11032\ : Odrv4
    port map (
            O => \N__47530\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7\
        );

    \I__11031\ : LocalMux
    port map (
            O => \N__47527\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7\
        );

    \I__11030\ : InMux
    port map (
            O => \N__47522\,
            I => \N__47515\
        );

    \I__11029\ : InMux
    port map (
            O => \N__47521\,
            I => \N__47515\
        );

    \I__11028\ : InMux
    port map (
            O => \N__47520\,
            I => \N__47512\
        );

    \I__11027\ : LocalMux
    port map (
            O => \N__47515\,
            I => \N__47509\
        );

    \I__11026\ : LocalMux
    port map (
            O => \N__47512\,
            I => \N__47505\
        );

    \I__11025\ : Span12Mux_v
    port map (
            O => \N__47509\,
            I => \N__47502\
        );

    \I__11024\ : InMux
    port map (
            O => \N__47508\,
            I => \N__47499\
        );

    \I__11023\ : Odrv4
    port map (
            O => \N__47505\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__11022\ : Odrv12
    port map (
            O => \N__47502\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__11021\ : LocalMux
    port map (
            O => \N__47499\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__11020\ : CascadeMux
    port map (
            O => \N__47492\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7_cascade_\
        );

    \I__11019\ : InMux
    port map (
            O => \N__47489\,
            I => \N__47486\
        );

    \I__11018\ : LocalMux
    port map (
            O => \N__47486\,
            I => \N__47483\
        );

    \I__11017\ : Span4Mux_h
    port map (
            O => \N__47483\,
            I => \N__47480\
        );

    \I__11016\ : Odrv4
    port map (
            O => \N__47480\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\
        );

    \I__11015\ : InMux
    port map (
            O => \N__47477\,
            I => \N__47472\
        );

    \I__11014\ : InMux
    port map (
            O => \N__47476\,
            I => \N__47469\
        );

    \I__11013\ : InMux
    port map (
            O => \N__47475\,
            I => \N__47466\
        );

    \I__11012\ : LocalMux
    port map (
            O => \N__47472\,
            I => \N__47461\
        );

    \I__11011\ : LocalMux
    port map (
            O => \N__47469\,
            I => \N__47461\
        );

    \I__11010\ : LocalMux
    port map (
            O => \N__47466\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29\
        );

    \I__11009\ : Odrv12
    port map (
            O => \N__47461\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29\
        );

    \I__11008\ : InMux
    port map (
            O => \N__47456\,
            I => \N__47452\
        );

    \I__11007\ : InMux
    port map (
            O => \N__47455\,
            I => \N__47449\
        );

    \I__11006\ : LocalMux
    port map (
            O => \N__47452\,
            I => \N__47444\
        );

    \I__11005\ : LocalMux
    port map (
            O => \N__47449\,
            I => \N__47441\
        );

    \I__11004\ : InMux
    port map (
            O => \N__47448\,
            I => \N__47438\
        );

    \I__11003\ : InMux
    port map (
            O => \N__47447\,
            I => \N__47435\
        );

    \I__11002\ : Span4Mux_v
    port map (
            O => \N__47444\,
            I => \N__47430\
        );

    \I__11001\ : Span4Mux_v
    port map (
            O => \N__47441\,
            I => \N__47430\
        );

    \I__11000\ : LocalMux
    port map (
            O => \N__47438\,
            I => \N__47427\
        );

    \I__10999\ : LocalMux
    port map (
            O => \N__47435\,
            I => \N__47424\
        );

    \I__10998\ : Span4Mux_h
    port map (
            O => \N__47430\,
            I => \N__47419\
        );

    \I__10997\ : Span4Mux_h
    port map (
            O => \N__47427\,
            I => \N__47419\
        );

    \I__10996\ : Span4Mux_h
    port map (
            O => \N__47424\,
            I => \N__47416\
        );

    \I__10995\ : Sp12to4
    port map (
            O => \N__47419\,
            I => \N__47413\
        );

    \I__10994\ : Odrv4
    port map (
            O => \N__47416\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__10993\ : Odrv12
    port map (
            O => \N__47413\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__10992\ : InMux
    port map (
            O => \N__47408\,
            I => \N__47405\
        );

    \I__10991\ : LocalMux
    port map (
            O => \N__47405\,
            I => \N__47402\
        );

    \I__10990\ : Span4Mux_h
    port map (
            O => \N__47402\,
            I => \N__47399\
        );

    \I__10989\ : Odrv4
    port map (
            O => \N__47399\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28\
        );

    \I__10988\ : InMux
    port map (
            O => \N__47396\,
            I => \N__47389\
        );

    \I__10987\ : InMux
    port map (
            O => \N__47395\,
            I => \N__47389\
        );

    \I__10986\ : InMux
    port map (
            O => \N__47394\,
            I => \N__47386\
        );

    \I__10985\ : LocalMux
    port map (
            O => \N__47389\,
            I => \N__47383\
        );

    \I__10984\ : LocalMux
    port map (
            O => \N__47386\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__10983\ : Odrv4
    port map (
            O => \N__47383\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__10982\ : CascadeMux
    port map (
            O => \N__47378\,
            I => \N__47375\
        );

    \I__10981\ : InMux
    port map (
            O => \N__47375\,
            I => \N__47368\
        );

    \I__10980\ : InMux
    port map (
            O => \N__47374\,
            I => \N__47368\
        );

    \I__10979\ : InMux
    port map (
            O => \N__47373\,
            I => \N__47365\
        );

    \I__10978\ : LocalMux
    port map (
            O => \N__47368\,
            I => \N__47362\
        );

    \I__10977\ : LocalMux
    port map (
            O => \N__47365\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__10976\ : Odrv4
    port map (
            O => \N__47362\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__10975\ : CascadeMux
    port map (
            O => \N__47357\,
            I => \N__47354\
        );

    \I__10974\ : InMux
    port map (
            O => \N__47354\,
            I => \N__47348\
        );

    \I__10973\ : InMux
    port map (
            O => \N__47353\,
            I => \N__47348\
        );

    \I__10972\ : LocalMux
    port map (
            O => \N__47348\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_29\
        );

    \I__10971\ : CascadeMux
    port map (
            O => \N__47345\,
            I => \N__47342\
        );

    \I__10970\ : InMux
    port map (
            O => \N__47342\,
            I => \N__47339\
        );

    \I__10969\ : LocalMux
    port map (
            O => \N__47339\,
            I => \N__47336\
        );

    \I__10968\ : Span4Mux_h
    port map (
            O => \N__47336\,
            I => \N__47333\
        );

    \I__10967\ : Odrv4
    port map (
            O => \N__47333\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt28\
        );

    \I__10966\ : InMux
    port map (
            O => \N__47330\,
            I => \N__47327\
        );

    \I__10965\ : LocalMux
    port map (
            O => \N__47327\,
            I => \N__47324\
        );

    \I__10964\ : Span4Mux_h
    port map (
            O => \N__47324\,
            I => \N__47320\
        );

    \I__10963\ : InMux
    port map (
            O => \N__47323\,
            I => \N__47317\
        );

    \I__10962\ : Odrv4
    port map (
            O => \N__47320\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28\
        );

    \I__10961\ : LocalMux
    port map (
            O => \N__47317\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28\
        );

    \I__10960\ : InMux
    port map (
            O => \N__47312\,
            I => \N__47306\
        );

    \I__10959\ : InMux
    port map (
            O => \N__47311\,
            I => \N__47306\
        );

    \I__10958\ : LocalMux
    port map (
            O => \N__47306\,
            I => \N__47302\
        );

    \I__10957\ : InMux
    port map (
            O => \N__47305\,
            I => \N__47298\
        );

    \I__10956\ : Span4Mux_v
    port map (
            O => \N__47302\,
            I => \N__47295\
        );

    \I__10955\ : InMux
    port map (
            O => \N__47301\,
            I => \N__47292\
        );

    \I__10954\ : LocalMux
    port map (
            O => \N__47298\,
            I => \N__47289\
        );

    \I__10953\ : Span4Mux_v
    port map (
            O => \N__47295\,
            I => \N__47284\
        );

    \I__10952\ : LocalMux
    port map (
            O => \N__47292\,
            I => \N__47284\
        );

    \I__10951\ : Span4Mux_v
    port map (
            O => \N__47289\,
            I => \N__47281\
        );

    \I__10950\ : Span4Mux_h
    port map (
            O => \N__47284\,
            I => \N__47278\
        );

    \I__10949\ : Odrv4
    port map (
            O => \N__47281\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__10948\ : Odrv4
    port map (
            O => \N__47278\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__10947\ : CascadeMux
    port map (
            O => \N__47273\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28_cascade_\
        );

    \I__10946\ : InMux
    port map (
            O => \N__47270\,
            I => \N__47264\
        );

    \I__10945\ : InMux
    port map (
            O => \N__47269\,
            I => \N__47264\
        );

    \I__10944\ : LocalMux
    port map (
            O => \N__47264\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_28\
        );

    \I__10943\ : InMux
    port map (
            O => \N__47261\,
            I => \N__47255\
        );

    \I__10942\ : InMux
    port map (
            O => \N__47260\,
            I => \N__47255\
        );

    \I__10941\ : LocalMux
    port map (
            O => \N__47255\,
            I => \N__47252\
        );

    \I__10940\ : Odrv4
    port map (
            O => \N__47252\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\
        );

    \I__10939\ : InMux
    port map (
            O => \N__47249\,
            I => \N__47245\
        );

    \I__10938\ : InMux
    port map (
            O => \N__47248\,
            I => \N__47242\
        );

    \I__10937\ : LocalMux
    port map (
            O => \N__47245\,
            I => \N__47237\
        );

    \I__10936\ : LocalMux
    port map (
            O => \N__47242\,
            I => \N__47237\
        );

    \I__10935\ : Odrv4
    port map (
            O => \N__47237\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\
        );

    \I__10934\ : InMux
    port map (
            O => \N__47234\,
            I => \N__47231\
        );

    \I__10933\ : LocalMux
    port map (
            O => \N__47231\,
            I => \N__47228\
        );

    \I__10932\ : Span4Mux_h
    port map (
            O => \N__47228\,
            I => \N__47224\
        );

    \I__10931\ : InMux
    port map (
            O => \N__47227\,
            I => \N__47221\
        );

    \I__10930\ : Odrv4
    port map (
            O => \N__47224\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17\
        );

    \I__10929\ : LocalMux
    port map (
            O => \N__47221\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17\
        );

    \I__10928\ : InMux
    port map (
            O => \N__47216\,
            I => \N__47210\
        );

    \I__10927\ : InMux
    port map (
            O => \N__47215\,
            I => \N__47210\
        );

    \I__10926\ : LocalMux
    port map (
            O => \N__47210\,
            I => \N__47206\
        );

    \I__10925\ : InMux
    port map (
            O => \N__47209\,
            I => \N__47203\
        );

    \I__10924\ : Span4Mux_h
    port map (
            O => \N__47206\,
            I => \N__47200\
        );

    \I__10923\ : LocalMux
    port map (
            O => \N__47203\,
            I => \N__47196\
        );

    \I__10922\ : Span4Mux_h
    port map (
            O => \N__47200\,
            I => \N__47193\
        );

    \I__10921\ : InMux
    port map (
            O => \N__47199\,
            I => \N__47190\
        );

    \I__10920\ : Odrv4
    port map (
            O => \N__47196\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__10919\ : Odrv4
    port map (
            O => \N__47193\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__10918\ : LocalMux
    port map (
            O => \N__47190\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__10917\ : CascadeMux
    port map (
            O => \N__47183\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17_cascade_\
        );

    \I__10916\ : InMux
    port map (
            O => \N__47180\,
            I => \N__47175\
        );

    \I__10915\ : InMux
    port map (
            O => \N__47179\,
            I => \N__47170\
        );

    \I__10914\ : InMux
    port map (
            O => \N__47178\,
            I => \N__47170\
        );

    \I__10913\ : LocalMux
    port map (
            O => \N__47175\,
            I => \N__47165\
        );

    \I__10912\ : LocalMux
    port map (
            O => \N__47170\,
            I => \N__47165\
        );

    \I__10911\ : Odrv4
    port map (
            O => \N__47165\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__10910\ : CascadeMux
    port map (
            O => \N__47162\,
            I => \N__47158\
        );

    \I__10909\ : CascadeMux
    port map (
            O => \N__47161\,
            I => \N__47155\
        );

    \I__10908\ : InMux
    port map (
            O => \N__47158\,
            I => \N__47150\
        );

    \I__10907\ : InMux
    port map (
            O => \N__47155\,
            I => \N__47150\
        );

    \I__10906\ : LocalMux
    port map (
            O => \N__47150\,
            I => \N__47146\
        );

    \I__10905\ : InMux
    port map (
            O => \N__47149\,
            I => \N__47143\
        );

    \I__10904\ : Span4Mux_v
    port map (
            O => \N__47146\,
            I => \N__47140\
        );

    \I__10903\ : LocalMux
    port map (
            O => \N__47143\,
            I => \N__47135\
        );

    \I__10902\ : Span4Mux_h
    port map (
            O => \N__47140\,
            I => \N__47135\
        );

    \I__10901\ : Odrv4
    port map (
            O => \N__47135\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__10900\ : InMux
    port map (
            O => \N__47132\,
            I => \N__47126\
        );

    \I__10899\ : InMux
    port map (
            O => \N__47131\,
            I => \N__47126\
        );

    \I__10898\ : LocalMux
    port map (
            O => \N__47126\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\
        );

    \I__10897\ : InMux
    port map (
            O => \N__47123\,
            I => \N__47120\
        );

    \I__10896\ : LocalMux
    port map (
            O => \N__47120\,
            I => \N__47117\
        );

    \I__10895\ : Span4Mux_h
    port map (
            O => \N__47117\,
            I => \N__47114\
        );

    \I__10894\ : Odrv4
    port map (
            O => \N__47114\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\
        );

    \I__10893\ : InMux
    port map (
            O => \N__47111\,
            I => \N__47108\
        );

    \I__10892\ : LocalMux
    port map (
            O => \N__47108\,
            I => \N__47104\
        );

    \I__10891\ : InMux
    port map (
            O => \N__47107\,
            I => \N__47101\
        );

    \I__10890\ : Span4Mux_v
    port map (
            O => \N__47104\,
            I => \N__47098\
        );

    \I__10889\ : LocalMux
    port map (
            O => \N__47101\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14\
        );

    \I__10888\ : Odrv4
    port map (
            O => \N__47098\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14\
        );

    \I__10887\ : InMux
    port map (
            O => \N__47093\,
            I => \N__47086\
        );

    \I__10886\ : InMux
    port map (
            O => \N__47092\,
            I => \N__47086\
        );

    \I__10885\ : InMux
    port map (
            O => \N__47091\,
            I => \N__47083\
        );

    \I__10884\ : LocalMux
    port map (
            O => \N__47086\,
            I => \N__47080\
        );

    \I__10883\ : LocalMux
    port map (
            O => \N__47083\,
            I => \N__47076\
        );

    \I__10882\ : Span4Mux_v
    port map (
            O => \N__47080\,
            I => \N__47073\
        );

    \I__10881\ : InMux
    port map (
            O => \N__47079\,
            I => \N__47070\
        );

    \I__10880\ : Odrv4
    port map (
            O => \N__47076\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__10879\ : Odrv4
    port map (
            O => \N__47073\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__10878\ : LocalMux
    port map (
            O => \N__47070\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__10877\ : CascadeMux
    port map (
            O => \N__47063\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14_cascade_\
        );

    \I__10876\ : InMux
    port map (
            O => \N__47060\,
            I => \N__47057\
        );

    \I__10875\ : LocalMux
    port map (
            O => \N__47057\,
            I => \N__47054\
        );

    \I__10874\ : Span4Mux_h
    port map (
            O => \N__47054\,
            I => \N__47051\
        );

    \I__10873\ : Odrv4
    port map (
            O => \N__47051\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\
        );

    \I__10872\ : InMux
    port map (
            O => \N__47048\,
            I => \N__47042\
        );

    \I__10871\ : InMux
    port map (
            O => \N__47047\,
            I => \N__47042\
        );

    \I__10870\ : LocalMux
    port map (
            O => \N__47042\,
            I => \N__47039\
        );

    \I__10869\ : Odrv12
    port map (
            O => \N__47039\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\
        );

    \I__10868\ : CascadeMux
    port map (
            O => \N__47036\,
            I => \N__47033\
        );

    \I__10867\ : InMux
    port map (
            O => \N__47033\,
            I => \N__47027\
        );

    \I__10866\ : InMux
    port map (
            O => \N__47032\,
            I => \N__47027\
        );

    \I__10865\ : LocalMux
    port map (
            O => \N__47027\,
            I => \N__47024\
        );

    \I__10864\ : Span4Mux_h
    port map (
            O => \N__47024\,
            I => \N__47021\
        );

    \I__10863\ : Odrv4
    port map (
            O => \N__47021\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_29\
        );

    \I__10862\ : InMux
    port map (
            O => \N__47018\,
            I => \N__47015\
        );

    \I__10861\ : LocalMux
    port map (
            O => \N__47015\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15\
        );

    \I__10860\ : InMux
    port map (
            O => \N__47012\,
            I => \N__47009\
        );

    \I__10859\ : LocalMux
    port map (
            O => \N__47009\,
            I => \N__47006\
        );

    \I__10858\ : Odrv12
    port map (
            O => \N__47006\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\
        );

    \I__10857\ : InMux
    port map (
            O => \N__47003\,
            I => \N__46999\
        );

    \I__10856\ : InMux
    port map (
            O => \N__47002\,
            I => \N__46996\
        );

    \I__10855\ : LocalMux
    port map (
            O => \N__46999\,
            I => \N__46993\
        );

    \I__10854\ : LocalMux
    port map (
            O => \N__46996\,
            I => \phase_controller_inst1.stoper_hc.runningZ0\
        );

    \I__10853\ : Odrv4
    port map (
            O => \N__46993\,
            I => \phase_controller_inst1.stoper_hc.runningZ0\
        );

    \I__10852\ : InMux
    port map (
            O => \N__46988\,
            I => \N__46982\
        );

    \I__10851\ : InMux
    port map (
            O => \N__46987\,
            I => \N__46974\
        );

    \I__10850\ : InMux
    port map (
            O => \N__46986\,
            I => \N__46974\
        );

    \I__10849\ : InMux
    port map (
            O => \N__46985\,
            I => \N__46974\
        );

    \I__10848\ : LocalMux
    port map (
            O => \N__46982\,
            I => \N__46971\
        );

    \I__10847\ : InMux
    port map (
            O => \N__46981\,
            I => \N__46968\
        );

    \I__10846\ : LocalMux
    port map (
            O => \N__46974\,
            I => \N__46965\
        );

    \I__10845\ : Odrv12
    port map (
            O => \N__46971\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__10844\ : LocalMux
    port map (
            O => \N__46968\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__10843\ : Odrv4
    port map (
            O => \N__46965\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__10842\ : InMux
    port map (
            O => \N__46958\,
            I => \N__46954\
        );

    \I__10841\ : CascadeMux
    port map (
            O => \N__46957\,
            I => \N__46951\
        );

    \I__10840\ : LocalMux
    port map (
            O => \N__46954\,
            I => \N__46947\
        );

    \I__10839\ : InMux
    port map (
            O => \N__46951\,
            I => \N__46942\
        );

    \I__10838\ : InMux
    port map (
            O => \N__46950\,
            I => \N__46942\
        );

    \I__10837\ : Span4Mux_h
    port map (
            O => \N__46947\,
            I => \N__46939\
        );

    \I__10836\ : LocalMux
    port map (
            O => \N__46942\,
            I => \N__46936\
        );

    \I__10835\ : Odrv4
    port map (
            O => \N__46939\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__10834\ : Odrv4
    port map (
            O => \N__46936\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__10833\ : CascadeMux
    port map (
            O => \N__46931\,
            I => \N__46927\
        );

    \I__10832\ : InMux
    port map (
            O => \N__46930\,
            I => \N__46923\
        );

    \I__10831\ : InMux
    port map (
            O => \N__46927\,
            I => \N__46920\
        );

    \I__10830\ : InMux
    port map (
            O => \N__46926\,
            I => \N__46917\
        );

    \I__10829\ : LocalMux
    port map (
            O => \N__46923\,
            I => \N__46913\
        );

    \I__10828\ : LocalMux
    port map (
            O => \N__46920\,
            I => \N__46910\
        );

    \I__10827\ : LocalMux
    port map (
            O => \N__46917\,
            I => \N__46907\
        );

    \I__10826\ : CascadeMux
    port map (
            O => \N__46916\,
            I => \N__46904\
        );

    \I__10825\ : Span4Mux_h
    port map (
            O => \N__46913\,
            I => \N__46901\
        );

    \I__10824\ : Span4Mux_v
    port map (
            O => \N__46910\,
            I => \N__46896\
        );

    \I__10823\ : Span4Mux_h
    port map (
            O => \N__46907\,
            I => \N__46896\
        );

    \I__10822\ : InMux
    port map (
            O => \N__46904\,
            I => \N__46891\
        );

    \I__10821\ : Span4Mux_h
    port map (
            O => \N__46901\,
            I => \N__46888\
        );

    \I__10820\ : Span4Mux_h
    port map (
            O => \N__46896\,
            I => \N__46885\
        );

    \I__10819\ : InMux
    port map (
            O => \N__46895\,
            I => \N__46880\
        );

    \I__10818\ : InMux
    port map (
            O => \N__46894\,
            I => \N__46880\
        );

    \I__10817\ : LocalMux
    port map (
            O => \N__46891\,
            I => phase_controller_inst1_state_4
        );

    \I__10816\ : Odrv4
    port map (
            O => \N__46888\,
            I => phase_controller_inst1_state_4
        );

    \I__10815\ : Odrv4
    port map (
            O => \N__46885\,
            I => phase_controller_inst1_state_4
        );

    \I__10814\ : LocalMux
    port map (
            O => \N__46880\,
            I => phase_controller_inst1_state_4
        );

    \I__10813\ : InMux
    port map (
            O => \N__46871\,
            I => \N__46868\
        );

    \I__10812\ : LocalMux
    port map (
            O => \N__46868\,
            I => \N__46865\
        );

    \I__10811\ : Span4Mux_v
    port map (
            O => \N__46865\,
            I => \N__46862\
        );

    \I__10810\ : Span4Mux_h
    port map (
            O => \N__46862\,
            I => \N__46859\
        );

    \I__10809\ : Odrv4
    port map (
            O => \N__46859\,
            I => \phase_controller_inst1.start_timer_hc_0_sqmuxa\
        );

    \I__10808\ : CascadeMux
    port map (
            O => \N__46856\,
            I => \N__46853\
        );

    \I__10807\ : InMux
    port map (
            O => \N__46853\,
            I => \N__46845\
        );

    \I__10806\ : InMux
    port map (
            O => \N__46852\,
            I => \N__46845\
        );

    \I__10805\ : InMux
    port map (
            O => \N__46851\,
            I => \N__46840\
        );

    \I__10804\ : InMux
    port map (
            O => \N__46850\,
            I => \N__46840\
        );

    \I__10803\ : LocalMux
    port map (
            O => \N__46845\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__10802\ : LocalMux
    port map (
            O => \N__46840\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__10801\ : InMux
    port map (
            O => \N__46835\,
            I => \N__46828\
        );

    \I__10800\ : InMux
    port map (
            O => \N__46834\,
            I => \N__46828\
        );

    \I__10799\ : CascadeMux
    port map (
            O => \N__46833\,
            I => \N__46825\
        );

    \I__10798\ : LocalMux
    port map (
            O => \N__46828\,
            I => \N__46822\
        );

    \I__10797\ : InMux
    port map (
            O => \N__46825\,
            I => \N__46817\
        );

    \I__10796\ : Span4Mux_h
    port map (
            O => \N__46822\,
            I => \N__46814\
        );

    \I__10795\ : InMux
    port map (
            O => \N__46821\,
            I => \N__46809\
        );

    \I__10794\ : InMux
    port map (
            O => \N__46820\,
            I => \N__46809\
        );

    \I__10793\ : LocalMux
    port map (
            O => \N__46817\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__10792\ : Odrv4
    port map (
            O => \N__46814\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__10791\ : LocalMux
    port map (
            O => \N__46809\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__10790\ : CascadeMux
    port map (
            O => \N__46802\,
            I => \N__46799\
        );

    \I__10789\ : InMux
    port map (
            O => \N__46799\,
            I => \N__46796\
        );

    \I__10788\ : LocalMux
    port map (
            O => \N__46796\,
            I => \N__46793\
        );

    \I__10787\ : Span4Mux_v
    port map (
            O => \N__46793\,
            I => \N__46790\
        );

    \I__10786\ : Span4Mux_h
    port map (
            O => \N__46790\,
            I => \N__46787\
        );

    \I__10785\ : Span4Mux_s3_h
    port map (
            O => \N__46787\,
            I => \N__46784\
        );

    \I__10784\ : Odrv4
    port map (
            O => \N__46784\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt16\
        );

    \I__10783\ : CascadeMux
    port map (
            O => \N__46781\,
            I => \N__46778\
        );

    \I__10782\ : InMux
    port map (
            O => \N__46778\,
            I => \N__46773\
        );

    \I__10781\ : InMux
    port map (
            O => \N__46777\,
            I => \N__46770\
        );

    \I__10780\ : InMux
    port map (
            O => \N__46776\,
            I => \N__46767\
        );

    \I__10779\ : LocalMux
    port map (
            O => \N__46773\,
            I => \N__46762\
        );

    \I__10778\ : LocalMux
    port map (
            O => \N__46770\,
            I => \N__46762\
        );

    \I__10777\ : LocalMux
    port map (
            O => \N__46767\,
            I => \N__46757\
        );

    \I__10776\ : Span4Mux_v
    port map (
            O => \N__46762\,
            I => \N__46757\
        );

    \I__10775\ : Odrv4
    port map (
            O => \N__46757\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__10774\ : InMux
    port map (
            O => \N__46754\,
            I => \current_shift_inst.timer_s1.counter_cry_25\
        );

    \I__10773\ : CascadeMux
    port map (
            O => \N__46751\,
            I => \N__46748\
        );

    \I__10772\ : InMux
    port map (
            O => \N__46748\,
            I => \N__46744\
        );

    \I__10771\ : InMux
    port map (
            O => \N__46747\,
            I => \N__46741\
        );

    \I__10770\ : LocalMux
    port map (
            O => \N__46744\,
            I => \N__46735\
        );

    \I__10769\ : LocalMux
    port map (
            O => \N__46741\,
            I => \N__46735\
        );

    \I__10768\ : InMux
    port map (
            O => \N__46740\,
            I => \N__46732\
        );

    \I__10767\ : Span4Mux_v
    port map (
            O => \N__46735\,
            I => \N__46729\
        );

    \I__10766\ : LocalMux
    port map (
            O => \N__46732\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__10765\ : Odrv4
    port map (
            O => \N__46729\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__10764\ : InMux
    port map (
            O => \N__46724\,
            I => \current_shift_inst.timer_s1.counter_cry_26\
        );

    \I__10763\ : InMux
    port map (
            O => \N__46721\,
            I => \N__46718\
        );

    \I__10762\ : LocalMux
    port map (
            O => \N__46718\,
            I => \N__46714\
        );

    \I__10761\ : InMux
    port map (
            O => \N__46717\,
            I => \N__46711\
        );

    \I__10760\ : Span4Mux_h
    port map (
            O => \N__46714\,
            I => \N__46708\
        );

    \I__10759\ : LocalMux
    port map (
            O => \N__46711\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__10758\ : Odrv4
    port map (
            O => \N__46708\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__10757\ : InMux
    port map (
            O => \N__46703\,
            I => \current_shift_inst.timer_s1.counter_cry_27\
        );

    \I__10756\ : InMux
    port map (
            O => \N__46700\,
            I => \N__46684\
        );

    \I__10755\ : InMux
    port map (
            O => \N__46699\,
            I => \N__46684\
        );

    \I__10754\ : InMux
    port map (
            O => \N__46698\,
            I => \N__46684\
        );

    \I__10753\ : InMux
    port map (
            O => \N__46697\,
            I => \N__46684\
        );

    \I__10752\ : InMux
    port map (
            O => \N__46696\,
            I => \N__46675\
        );

    \I__10751\ : InMux
    port map (
            O => \N__46695\,
            I => \N__46675\
        );

    \I__10750\ : InMux
    port map (
            O => \N__46694\,
            I => \N__46675\
        );

    \I__10749\ : InMux
    port map (
            O => \N__46693\,
            I => \N__46675\
        );

    \I__10748\ : LocalMux
    port map (
            O => \N__46684\,
            I => \N__46648\
        );

    \I__10747\ : LocalMux
    port map (
            O => \N__46675\,
            I => \N__46648\
        );

    \I__10746\ : InMux
    port map (
            O => \N__46674\,
            I => \N__46639\
        );

    \I__10745\ : InMux
    port map (
            O => \N__46673\,
            I => \N__46639\
        );

    \I__10744\ : InMux
    port map (
            O => \N__46672\,
            I => \N__46639\
        );

    \I__10743\ : InMux
    port map (
            O => \N__46671\,
            I => \N__46639\
        );

    \I__10742\ : InMux
    port map (
            O => \N__46670\,
            I => \N__46634\
        );

    \I__10741\ : InMux
    port map (
            O => \N__46669\,
            I => \N__46634\
        );

    \I__10740\ : InMux
    port map (
            O => \N__46668\,
            I => \N__46625\
        );

    \I__10739\ : InMux
    port map (
            O => \N__46667\,
            I => \N__46625\
        );

    \I__10738\ : InMux
    port map (
            O => \N__46666\,
            I => \N__46625\
        );

    \I__10737\ : InMux
    port map (
            O => \N__46665\,
            I => \N__46625\
        );

    \I__10736\ : InMux
    port map (
            O => \N__46664\,
            I => \N__46616\
        );

    \I__10735\ : InMux
    port map (
            O => \N__46663\,
            I => \N__46616\
        );

    \I__10734\ : InMux
    port map (
            O => \N__46662\,
            I => \N__46616\
        );

    \I__10733\ : InMux
    port map (
            O => \N__46661\,
            I => \N__46616\
        );

    \I__10732\ : InMux
    port map (
            O => \N__46660\,
            I => \N__46607\
        );

    \I__10731\ : InMux
    port map (
            O => \N__46659\,
            I => \N__46607\
        );

    \I__10730\ : InMux
    port map (
            O => \N__46658\,
            I => \N__46607\
        );

    \I__10729\ : InMux
    port map (
            O => \N__46657\,
            I => \N__46607\
        );

    \I__10728\ : InMux
    port map (
            O => \N__46656\,
            I => \N__46598\
        );

    \I__10727\ : InMux
    port map (
            O => \N__46655\,
            I => \N__46598\
        );

    \I__10726\ : InMux
    port map (
            O => \N__46654\,
            I => \N__46598\
        );

    \I__10725\ : InMux
    port map (
            O => \N__46653\,
            I => \N__46598\
        );

    \I__10724\ : Span4Mux_h
    port map (
            O => \N__46648\,
            I => \N__46591\
        );

    \I__10723\ : LocalMux
    port map (
            O => \N__46639\,
            I => \N__46591\
        );

    \I__10722\ : LocalMux
    port map (
            O => \N__46634\,
            I => \N__46591\
        );

    \I__10721\ : LocalMux
    port map (
            O => \N__46625\,
            I => \N__46582\
        );

    \I__10720\ : LocalMux
    port map (
            O => \N__46616\,
            I => \N__46582\
        );

    \I__10719\ : LocalMux
    port map (
            O => \N__46607\,
            I => \N__46582\
        );

    \I__10718\ : LocalMux
    port map (
            O => \N__46598\,
            I => \N__46582\
        );

    \I__10717\ : Span4Mux_v
    port map (
            O => \N__46591\,
            I => \N__46577\
        );

    \I__10716\ : Span4Mux_v
    port map (
            O => \N__46582\,
            I => \N__46577\
        );

    \I__10715\ : Odrv4
    port map (
            O => \N__46577\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__10714\ : InMux
    port map (
            O => \N__46574\,
            I => \current_shift_inst.timer_s1.counter_cry_28\
        );

    \I__10713\ : InMux
    port map (
            O => \N__46571\,
            I => \N__46568\
        );

    \I__10712\ : LocalMux
    port map (
            O => \N__46568\,
            I => \N__46564\
        );

    \I__10711\ : InMux
    port map (
            O => \N__46567\,
            I => \N__46561\
        );

    \I__10710\ : Span4Mux_h
    port map (
            O => \N__46564\,
            I => \N__46558\
        );

    \I__10709\ : LocalMux
    port map (
            O => \N__46561\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__10708\ : Odrv4
    port map (
            O => \N__46558\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__10707\ : CEMux
    port map (
            O => \N__46553\,
            I => \N__46548\
        );

    \I__10706\ : CEMux
    port map (
            O => \N__46552\,
            I => \N__46545\
        );

    \I__10705\ : CEMux
    port map (
            O => \N__46551\,
            I => \N__46541\
        );

    \I__10704\ : LocalMux
    port map (
            O => \N__46548\,
            I => \N__46538\
        );

    \I__10703\ : LocalMux
    port map (
            O => \N__46545\,
            I => \N__46535\
        );

    \I__10702\ : CEMux
    port map (
            O => \N__46544\,
            I => \N__46532\
        );

    \I__10701\ : LocalMux
    port map (
            O => \N__46541\,
            I => \N__46529\
        );

    \I__10700\ : Span4Mux_v
    port map (
            O => \N__46538\,
            I => \N__46526\
        );

    \I__10699\ : Span4Mux_v
    port map (
            O => \N__46535\,
            I => \N__46523\
        );

    \I__10698\ : LocalMux
    port map (
            O => \N__46532\,
            I => \N__46520\
        );

    \I__10697\ : Span4Mux_h
    port map (
            O => \N__46529\,
            I => \N__46517\
        );

    \I__10696\ : Span4Mux_h
    port map (
            O => \N__46526\,
            I => \N__46514\
        );

    \I__10695\ : Span4Mux_h
    port map (
            O => \N__46523\,
            I => \N__46509\
        );

    \I__10694\ : Span4Mux_h
    port map (
            O => \N__46520\,
            I => \N__46509\
        );

    \I__10693\ : Odrv4
    port map (
            O => \N__46517\,
            I => \current_shift_inst.timer_s1.N_163_i\
        );

    \I__10692\ : Odrv4
    port map (
            O => \N__46514\,
            I => \current_shift_inst.timer_s1.N_163_i\
        );

    \I__10691\ : Odrv4
    port map (
            O => \N__46509\,
            I => \current_shift_inst.timer_s1.N_163_i\
        );

    \I__10690\ : IoInMux
    port map (
            O => \N__46502\,
            I => \N__46499\
        );

    \I__10689\ : LocalMux
    port map (
            O => \N__46499\,
            I => \N__46495\
        );

    \I__10688\ : InMux
    port map (
            O => \N__46498\,
            I => \N__46492\
        );

    \I__10687\ : Odrv12
    port map (
            O => \N__46495\,
            I => \T12_c\
        );

    \I__10686\ : LocalMux
    port map (
            O => \N__46492\,
            I => \T12_c\
        );

    \I__10685\ : InMux
    port map (
            O => \N__46487\,
            I => \N__46484\
        );

    \I__10684\ : LocalMux
    port map (
            O => \N__46484\,
            I => \N__46480\
        );

    \I__10683\ : InMux
    port map (
            O => \N__46483\,
            I => \N__46477\
        );

    \I__10682\ : Span4Mux_v
    port map (
            O => \N__46480\,
            I => \N__46471\
        );

    \I__10681\ : LocalMux
    port map (
            O => \N__46477\,
            I => \N__46471\
        );

    \I__10680\ : InMux
    port map (
            O => \N__46476\,
            I => \N__46468\
        );

    \I__10679\ : Span4Mux_h
    port map (
            O => \N__46471\,
            I => \N__46465\
        );

    \I__10678\ : LocalMux
    port map (
            O => \N__46468\,
            I => \elapsed_time_ns_1_RNIDV2T9_0_1\
        );

    \I__10677\ : Odrv4
    port map (
            O => \N__46465\,
            I => \elapsed_time_ns_1_RNIDV2T9_0_1\
        );

    \I__10676\ : InMux
    port map (
            O => \N__46460\,
            I => \N__46455\
        );

    \I__10675\ : InMux
    port map (
            O => \N__46459\,
            I => \N__46452\
        );

    \I__10674\ : InMux
    port map (
            O => \N__46458\,
            I => \N__46449\
        );

    \I__10673\ : LocalMux
    port map (
            O => \N__46455\,
            I => \N__46445\
        );

    \I__10672\ : LocalMux
    port map (
            O => \N__46452\,
            I => \N__46442\
        );

    \I__10671\ : LocalMux
    port map (
            O => \N__46449\,
            I => \N__46439\
        );

    \I__10670\ : InMux
    port map (
            O => \N__46448\,
            I => \N__46436\
        );

    \I__10669\ : Span4Mux_v
    port map (
            O => \N__46445\,
            I => \N__46431\
        );

    \I__10668\ : Span4Mux_v
    port map (
            O => \N__46442\,
            I => \N__46431\
        );

    \I__10667\ : Span4Mux_v
    port map (
            O => \N__46439\,
            I => \N__46428\
        );

    \I__10666\ : LocalMux
    port map (
            O => \N__46436\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__10665\ : Odrv4
    port map (
            O => \N__46431\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__10664\ : Odrv4
    port map (
            O => \N__46428\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__10663\ : InMux
    port map (
            O => \N__46421\,
            I => \N__46418\
        );

    \I__10662\ : LocalMux
    port map (
            O => \N__46418\,
            I => \N__46415\
        );

    \I__10661\ : Span4Mux_h
    port map (
            O => \N__46415\,
            I => \N__46410\
        );

    \I__10660\ : InMux
    port map (
            O => \N__46414\,
            I => \N__46406\
        );

    \I__10659\ : InMux
    port map (
            O => \N__46413\,
            I => \N__46403\
        );

    \I__10658\ : Span4Mux_v
    port map (
            O => \N__46410\,
            I => \N__46400\
        );

    \I__10657\ : InMux
    port map (
            O => \N__46409\,
            I => \N__46397\
        );

    \I__10656\ : LocalMux
    port map (
            O => \N__46406\,
            I => \N__46394\
        );

    \I__10655\ : LocalMux
    port map (
            O => \N__46403\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__10654\ : Odrv4
    port map (
            O => \N__46400\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__10653\ : LocalMux
    port map (
            O => \N__46397\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__10652\ : Odrv4
    port map (
            O => \N__46394\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__10651\ : CascadeMux
    port map (
            O => \N__46385\,
            I => \N__46380\
        );

    \I__10650\ : InMux
    port map (
            O => \N__46384\,
            I => \N__46376\
        );

    \I__10649\ : InMux
    port map (
            O => \N__46383\,
            I => \N__46373\
        );

    \I__10648\ : InMux
    port map (
            O => \N__46380\,
            I => \N__46370\
        );

    \I__10647\ : InMux
    port map (
            O => \N__46379\,
            I => \N__46367\
        );

    \I__10646\ : LocalMux
    port map (
            O => \N__46376\,
            I => \N__46364\
        );

    \I__10645\ : LocalMux
    port map (
            O => \N__46373\,
            I => \N__46361\
        );

    \I__10644\ : LocalMux
    port map (
            O => \N__46370\,
            I => \N__46358\
        );

    \I__10643\ : LocalMux
    port map (
            O => \N__46367\,
            I => \N__46355\
        );

    \I__10642\ : Span4Mux_v
    port map (
            O => \N__46364\,
            I => \N__46350\
        );

    \I__10641\ : Span4Mux_v
    port map (
            O => \N__46361\,
            I => \N__46350\
        );

    \I__10640\ : Span4Mux_v
    port map (
            O => \N__46358\,
            I => \N__46347\
        );

    \I__10639\ : Odrv4
    port map (
            O => \N__46355\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__10638\ : Odrv4
    port map (
            O => \N__46350\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__10637\ : Odrv4
    port map (
            O => \N__46347\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__10636\ : InMux
    port map (
            O => \N__46340\,
            I => \N__46336\
        );

    \I__10635\ : InMux
    port map (
            O => \N__46339\,
            I => \N__46332\
        );

    \I__10634\ : LocalMux
    port map (
            O => \N__46336\,
            I => \N__46328\
        );

    \I__10633\ : InMux
    port map (
            O => \N__46335\,
            I => \N__46325\
        );

    \I__10632\ : LocalMux
    port map (
            O => \N__46332\,
            I => \N__46322\
        );

    \I__10631\ : InMux
    port map (
            O => \N__46331\,
            I => \N__46319\
        );

    \I__10630\ : Span4Mux_h
    port map (
            O => \N__46328\,
            I => \N__46316\
        );

    \I__10629\ : LocalMux
    port map (
            O => \N__46325\,
            I => \N__46309\
        );

    \I__10628\ : Span4Mux_v
    port map (
            O => \N__46322\,
            I => \N__46309\
        );

    \I__10627\ : LocalMux
    port map (
            O => \N__46319\,
            I => \N__46309\
        );

    \I__10626\ : Odrv4
    port map (
            O => \N__46316\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__10625\ : Odrv4
    port map (
            O => \N__46309\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__10624\ : InMux
    port map (
            O => \N__46304\,
            I => \current_shift_inst.timer_s1.counter_cry_16\
        );

    \I__10623\ : CascadeMux
    port map (
            O => \N__46301\,
            I => \N__46298\
        );

    \I__10622\ : InMux
    port map (
            O => \N__46298\,
            I => \N__46293\
        );

    \I__10621\ : InMux
    port map (
            O => \N__46297\,
            I => \N__46290\
        );

    \I__10620\ : InMux
    port map (
            O => \N__46296\,
            I => \N__46287\
        );

    \I__10619\ : LocalMux
    port map (
            O => \N__46293\,
            I => \N__46282\
        );

    \I__10618\ : LocalMux
    port map (
            O => \N__46290\,
            I => \N__46282\
        );

    \I__10617\ : LocalMux
    port map (
            O => \N__46287\,
            I => \N__46277\
        );

    \I__10616\ : Span4Mux_v
    port map (
            O => \N__46282\,
            I => \N__46277\
        );

    \I__10615\ : Odrv4
    port map (
            O => \N__46277\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__10614\ : InMux
    port map (
            O => \N__46274\,
            I => \current_shift_inst.timer_s1.counter_cry_17\
        );

    \I__10613\ : InMux
    port map (
            O => \N__46271\,
            I => \N__46265\
        );

    \I__10612\ : InMux
    port map (
            O => \N__46270\,
            I => \N__46265\
        );

    \I__10611\ : LocalMux
    port map (
            O => \N__46265\,
            I => \N__46261\
        );

    \I__10610\ : InMux
    port map (
            O => \N__46264\,
            I => \N__46258\
        );

    \I__10609\ : Span4Mux_v
    port map (
            O => \N__46261\,
            I => \N__46255\
        );

    \I__10608\ : LocalMux
    port map (
            O => \N__46258\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__10607\ : Odrv4
    port map (
            O => \N__46255\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__10606\ : InMux
    port map (
            O => \N__46250\,
            I => \current_shift_inst.timer_s1.counter_cry_18\
        );

    \I__10605\ : CascadeMux
    port map (
            O => \N__46247\,
            I => \N__46244\
        );

    \I__10604\ : InMux
    port map (
            O => \N__46244\,
            I => \N__46240\
        );

    \I__10603\ : InMux
    port map (
            O => \N__46243\,
            I => \N__46237\
        );

    \I__10602\ : LocalMux
    port map (
            O => \N__46240\,
            I => \N__46231\
        );

    \I__10601\ : LocalMux
    port map (
            O => \N__46237\,
            I => \N__46231\
        );

    \I__10600\ : InMux
    port map (
            O => \N__46236\,
            I => \N__46228\
        );

    \I__10599\ : Span4Mux_h
    port map (
            O => \N__46231\,
            I => \N__46225\
        );

    \I__10598\ : LocalMux
    port map (
            O => \N__46228\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__10597\ : Odrv4
    port map (
            O => \N__46225\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__10596\ : InMux
    port map (
            O => \N__46220\,
            I => \current_shift_inst.timer_s1.counter_cry_19\
        );

    \I__10595\ : CascadeMux
    port map (
            O => \N__46217\,
            I => \N__46213\
        );

    \I__10594\ : CascadeMux
    port map (
            O => \N__46216\,
            I => \N__46210\
        );

    \I__10593\ : InMux
    port map (
            O => \N__46213\,
            I => \N__46205\
        );

    \I__10592\ : InMux
    port map (
            O => \N__46210\,
            I => \N__46205\
        );

    \I__10591\ : LocalMux
    port map (
            O => \N__46205\,
            I => \N__46201\
        );

    \I__10590\ : InMux
    port map (
            O => \N__46204\,
            I => \N__46198\
        );

    \I__10589\ : Span4Mux_h
    port map (
            O => \N__46201\,
            I => \N__46195\
        );

    \I__10588\ : LocalMux
    port map (
            O => \N__46198\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__10587\ : Odrv4
    port map (
            O => \N__46195\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__10586\ : InMux
    port map (
            O => \N__46190\,
            I => \current_shift_inst.timer_s1.counter_cry_20\
        );

    \I__10585\ : InMux
    port map (
            O => \N__46187\,
            I => \N__46181\
        );

    \I__10584\ : InMux
    port map (
            O => \N__46186\,
            I => \N__46181\
        );

    \I__10583\ : LocalMux
    port map (
            O => \N__46181\,
            I => \N__46177\
        );

    \I__10582\ : InMux
    port map (
            O => \N__46180\,
            I => \N__46174\
        );

    \I__10581\ : Span4Mux_h
    port map (
            O => \N__46177\,
            I => \N__46171\
        );

    \I__10580\ : LocalMux
    port map (
            O => \N__46174\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__10579\ : Odrv4
    port map (
            O => \N__46171\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__10578\ : InMux
    port map (
            O => \N__46166\,
            I => \current_shift_inst.timer_s1.counter_cry_21\
        );

    \I__10577\ : InMux
    port map (
            O => \N__46163\,
            I => \N__46157\
        );

    \I__10576\ : InMux
    port map (
            O => \N__46162\,
            I => \N__46157\
        );

    \I__10575\ : LocalMux
    port map (
            O => \N__46157\,
            I => \N__46153\
        );

    \I__10574\ : InMux
    port map (
            O => \N__46156\,
            I => \N__46150\
        );

    \I__10573\ : Span4Mux_h
    port map (
            O => \N__46153\,
            I => \N__46147\
        );

    \I__10572\ : LocalMux
    port map (
            O => \N__46150\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__10571\ : Odrv4
    port map (
            O => \N__46147\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__10570\ : InMux
    port map (
            O => \N__46142\,
            I => \current_shift_inst.timer_s1.counter_cry_22\
        );

    \I__10569\ : CascadeMux
    port map (
            O => \N__46139\,
            I => \N__46135\
        );

    \I__10568\ : CascadeMux
    port map (
            O => \N__46138\,
            I => \N__46132\
        );

    \I__10567\ : InMux
    port map (
            O => \N__46135\,
            I => \N__46129\
        );

    \I__10566\ : InMux
    port map (
            O => \N__46132\,
            I => \N__46126\
        );

    \I__10565\ : LocalMux
    port map (
            O => \N__46129\,
            I => \N__46122\
        );

    \I__10564\ : LocalMux
    port map (
            O => \N__46126\,
            I => \N__46119\
        );

    \I__10563\ : InMux
    port map (
            O => \N__46125\,
            I => \N__46116\
        );

    \I__10562\ : Span4Mux_h
    port map (
            O => \N__46122\,
            I => \N__46113\
        );

    \I__10561\ : Span4Mux_h
    port map (
            O => \N__46119\,
            I => \N__46110\
        );

    \I__10560\ : LocalMux
    port map (
            O => \N__46116\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__10559\ : Odrv4
    port map (
            O => \N__46113\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__10558\ : Odrv4
    port map (
            O => \N__46110\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__10557\ : InMux
    port map (
            O => \N__46103\,
            I => \bfn_18_20_0_\
        );

    \I__10556\ : CascadeMux
    port map (
            O => \N__46100\,
            I => \N__46096\
        );

    \I__10555\ : CascadeMux
    port map (
            O => \N__46099\,
            I => \N__46093\
        );

    \I__10554\ : InMux
    port map (
            O => \N__46096\,
            I => \N__46090\
        );

    \I__10553\ : InMux
    port map (
            O => \N__46093\,
            I => \N__46087\
        );

    \I__10552\ : LocalMux
    port map (
            O => \N__46090\,
            I => \N__46083\
        );

    \I__10551\ : LocalMux
    port map (
            O => \N__46087\,
            I => \N__46080\
        );

    \I__10550\ : InMux
    port map (
            O => \N__46086\,
            I => \N__46077\
        );

    \I__10549\ : Span4Mux_h
    port map (
            O => \N__46083\,
            I => \N__46074\
        );

    \I__10548\ : Span4Mux_h
    port map (
            O => \N__46080\,
            I => \N__46071\
        );

    \I__10547\ : LocalMux
    port map (
            O => \N__46077\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__10546\ : Odrv4
    port map (
            O => \N__46074\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__10545\ : Odrv4
    port map (
            O => \N__46071\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__10544\ : InMux
    port map (
            O => \N__46064\,
            I => \current_shift_inst.timer_s1.counter_cry_24\
        );

    \I__10543\ : CascadeMux
    port map (
            O => \N__46061\,
            I => \N__46058\
        );

    \I__10542\ : InMux
    port map (
            O => \N__46058\,
            I => \N__46054\
        );

    \I__10541\ : InMux
    port map (
            O => \N__46057\,
            I => \N__46051\
        );

    \I__10540\ : LocalMux
    port map (
            O => \N__46054\,
            I => \N__46047\
        );

    \I__10539\ : LocalMux
    port map (
            O => \N__46051\,
            I => \N__46044\
        );

    \I__10538\ : InMux
    port map (
            O => \N__46050\,
            I => \N__46041\
        );

    \I__10537\ : Span4Mux_h
    port map (
            O => \N__46047\,
            I => \N__46038\
        );

    \I__10536\ : Span4Mux_h
    port map (
            O => \N__46044\,
            I => \N__46035\
        );

    \I__10535\ : LocalMux
    port map (
            O => \N__46041\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__10534\ : Odrv4
    port map (
            O => \N__46038\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__10533\ : Odrv4
    port map (
            O => \N__46035\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__10532\ : InMux
    port map (
            O => \N__46028\,
            I => \current_shift_inst.timer_s1.counter_cry_8\
        );

    \I__10531\ : InMux
    port map (
            O => \N__46025\,
            I => \N__46018\
        );

    \I__10530\ : InMux
    port map (
            O => \N__46024\,
            I => \N__46018\
        );

    \I__10529\ : InMux
    port map (
            O => \N__46023\,
            I => \N__46015\
        );

    \I__10528\ : LocalMux
    port map (
            O => \N__46018\,
            I => \N__46012\
        );

    \I__10527\ : LocalMux
    port map (
            O => \N__46015\,
            I => \N__46007\
        );

    \I__10526\ : Span4Mux_v
    port map (
            O => \N__46012\,
            I => \N__46007\
        );

    \I__10525\ : Odrv4
    port map (
            O => \N__46007\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__10524\ : InMux
    port map (
            O => \N__46004\,
            I => \current_shift_inst.timer_s1.counter_cry_9\
        );

    \I__10523\ : InMux
    port map (
            O => \N__46001\,
            I => \N__45995\
        );

    \I__10522\ : InMux
    port map (
            O => \N__46000\,
            I => \N__45995\
        );

    \I__10521\ : LocalMux
    port map (
            O => \N__45995\,
            I => \N__45991\
        );

    \I__10520\ : InMux
    port map (
            O => \N__45994\,
            I => \N__45988\
        );

    \I__10519\ : Span4Mux_v
    port map (
            O => \N__45991\,
            I => \N__45985\
        );

    \I__10518\ : LocalMux
    port map (
            O => \N__45988\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__10517\ : Odrv4
    port map (
            O => \N__45985\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__10516\ : InMux
    port map (
            O => \N__45980\,
            I => \current_shift_inst.timer_s1.counter_cry_10\
        );

    \I__10515\ : CascadeMux
    port map (
            O => \N__45977\,
            I => \N__45973\
        );

    \I__10514\ : CascadeMux
    port map (
            O => \N__45976\,
            I => \N__45970\
        );

    \I__10513\ : InMux
    port map (
            O => \N__45973\,
            I => \N__45965\
        );

    \I__10512\ : InMux
    port map (
            O => \N__45970\,
            I => \N__45965\
        );

    \I__10511\ : LocalMux
    port map (
            O => \N__45965\,
            I => \N__45961\
        );

    \I__10510\ : InMux
    port map (
            O => \N__45964\,
            I => \N__45958\
        );

    \I__10509\ : Span4Mux_h
    port map (
            O => \N__45961\,
            I => \N__45955\
        );

    \I__10508\ : LocalMux
    port map (
            O => \N__45958\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__10507\ : Odrv4
    port map (
            O => \N__45955\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__10506\ : InMux
    port map (
            O => \N__45950\,
            I => \current_shift_inst.timer_s1.counter_cry_11\
        );

    \I__10505\ : CascadeMux
    port map (
            O => \N__45947\,
            I => \N__45943\
        );

    \I__10504\ : CascadeMux
    port map (
            O => \N__45946\,
            I => \N__45940\
        );

    \I__10503\ : InMux
    port map (
            O => \N__45943\,
            I => \N__45935\
        );

    \I__10502\ : InMux
    port map (
            O => \N__45940\,
            I => \N__45935\
        );

    \I__10501\ : LocalMux
    port map (
            O => \N__45935\,
            I => \N__45931\
        );

    \I__10500\ : InMux
    port map (
            O => \N__45934\,
            I => \N__45928\
        );

    \I__10499\ : Span4Mux_h
    port map (
            O => \N__45931\,
            I => \N__45925\
        );

    \I__10498\ : LocalMux
    port map (
            O => \N__45928\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__10497\ : Odrv4
    port map (
            O => \N__45925\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__10496\ : InMux
    port map (
            O => \N__45920\,
            I => \current_shift_inst.timer_s1.counter_cry_12\
        );

    \I__10495\ : InMux
    port map (
            O => \N__45917\,
            I => \N__45911\
        );

    \I__10494\ : InMux
    port map (
            O => \N__45916\,
            I => \N__45911\
        );

    \I__10493\ : LocalMux
    port map (
            O => \N__45911\,
            I => \N__45907\
        );

    \I__10492\ : InMux
    port map (
            O => \N__45910\,
            I => \N__45904\
        );

    \I__10491\ : Span4Mux_h
    port map (
            O => \N__45907\,
            I => \N__45901\
        );

    \I__10490\ : LocalMux
    port map (
            O => \N__45904\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__10489\ : Odrv4
    port map (
            O => \N__45901\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__10488\ : InMux
    port map (
            O => \N__45896\,
            I => \current_shift_inst.timer_s1.counter_cry_13\
        );

    \I__10487\ : CascadeMux
    port map (
            O => \N__45893\,
            I => \N__45890\
        );

    \I__10486\ : InMux
    port map (
            O => \N__45890\,
            I => \N__45886\
        );

    \I__10485\ : InMux
    port map (
            O => \N__45889\,
            I => \N__45883\
        );

    \I__10484\ : LocalMux
    port map (
            O => \N__45886\,
            I => \N__45877\
        );

    \I__10483\ : LocalMux
    port map (
            O => \N__45883\,
            I => \N__45877\
        );

    \I__10482\ : InMux
    port map (
            O => \N__45882\,
            I => \N__45874\
        );

    \I__10481\ : Span4Mux_h
    port map (
            O => \N__45877\,
            I => \N__45871\
        );

    \I__10480\ : LocalMux
    port map (
            O => \N__45874\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__10479\ : Odrv4
    port map (
            O => \N__45871\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__10478\ : InMux
    port map (
            O => \N__45866\,
            I => \current_shift_inst.timer_s1.counter_cry_14\
        );

    \I__10477\ : CascadeMux
    port map (
            O => \N__45863\,
            I => \N__45859\
        );

    \I__10476\ : CascadeMux
    port map (
            O => \N__45862\,
            I => \N__45856\
        );

    \I__10475\ : InMux
    port map (
            O => \N__45859\,
            I => \N__45853\
        );

    \I__10474\ : InMux
    port map (
            O => \N__45856\,
            I => \N__45850\
        );

    \I__10473\ : LocalMux
    port map (
            O => \N__45853\,
            I => \N__45846\
        );

    \I__10472\ : LocalMux
    port map (
            O => \N__45850\,
            I => \N__45843\
        );

    \I__10471\ : InMux
    port map (
            O => \N__45849\,
            I => \N__45840\
        );

    \I__10470\ : Span4Mux_h
    port map (
            O => \N__45846\,
            I => \N__45837\
        );

    \I__10469\ : Span4Mux_h
    port map (
            O => \N__45843\,
            I => \N__45834\
        );

    \I__10468\ : LocalMux
    port map (
            O => \N__45840\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__10467\ : Odrv4
    port map (
            O => \N__45837\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__10466\ : Odrv4
    port map (
            O => \N__45834\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__10465\ : InMux
    port map (
            O => \N__45827\,
            I => \bfn_18_19_0_\
        );

    \I__10464\ : CascadeMux
    port map (
            O => \N__45824\,
            I => \N__45821\
        );

    \I__10463\ : InMux
    port map (
            O => \N__45821\,
            I => \N__45817\
        );

    \I__10462\ : InMux
    port map (
            O => \N__45820\,
            I => \N__45814\
        );

    \I__10461\ : LocalMux
    port map (
            O => \N__45817\,
            I => \N__45810\
        );

    \I__10460\ : LocalMux
    port map (
            O => \N__45814\,
            I => \N__45807\
        );

    \I__10459\ : InMux
    port map (
            O => \N__45813\,
            I => \N__45804\
        );

    \I__10458\ : Span4Mux_h
    port map (
            O => \N__45810\,
            I => \N__45801\
        );

    \I__10457\ : Span4Mux_h
    port map (
            O => \N__45807\,
            I => \N__45798\
        );

    \I__10456\ : LocalMux
    port map (
            O => \N__45804\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__10455\ : Odrv4
    port map (
            O => \N__45801\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__10454\ : Odrv4
    port map (
            O => \N__45798\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__10453\ : InMux
    port map (
            O => \N__45791\,
            I => \N__45787\
        );

    \I__10452\ : InMux
    port map (
            O => \N__45790\,
            I => \N__45784\
        );

    \I__10451\ : LocalMux
    port map (
            O => \N__45787\,
            I => \N__45780\
        );

    \I__10450\ : LocalMux
    port map (
            O => \N__45784\,
            I => \N__45777\
        );

    \I__10449\ : InMux
    port map (
            O => \N__45783\,
            I => \N__45774\
        );

    \I__10448\ : Span4Mux_h
    port map (
            O => \N__45780\,
            I => \N__45771\
        );

    \I__10447\ : Odrv4
    port map (
            O => \N__45777\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__10446\ : LocalMux
    port map (
            O => \N__45774\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__10445\ : Odrv4
    port map (
            O => \N__45771\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__10444\ : InMux
    port map (
            O => \N__45764\,
            I => \current_shift_inst.timer_s1.counter_cry_0\
        );

    \I__10443\ : CascadeMux
    port map (
            O => \N__45761\,
            I => \N__45757\
        );

    \I__10442\ : CascadeMux
    port map (
            O => \N__45760\,
            I => \N__45754\
        );

    \I__10441\ : InMux
    port map (
            O => \N__45757\,
            I => \N__45748\
        );

    \I__10440\ : InMux
    port map (
            O => \N__45754\,
            I => \N__45748\
        );

    \I__10439\ : InMux
    port map (
            O => \N__45753\,
            I => \N__45745\
        );

    \I__10438\ : LocalMux
    port map (
            O => \N__45748\,
            I => \N__45742\
        );

    \I__10437\ : LocalMux
    port map (
            O => \N__45745\,
            I => \N__45737\
        );

    \I__10436\ : Span4Mux_v
    port map (
            O => \N__45742\,
            I => \N__45737\
        );

    \I__10435\ : Odrv4
    port map (
            O => \N__45737\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__10434\ : InMux
    port map (
            O => \N__45734\,
            I => \current_shift_inst.timer_s1.counter_cry_1\
        );

    \I__10433\ : CascadeMux
    port map (
            O => \N__45731\,
            I => \N__45727\
        );

    \I__10432\ : CascadeMux
    port map (
            O => \N__45730\,
            I => \N__45724\
        );

    \I__10431\ : InMux
    port map (
            O => \N__45727\,
            I => \N__45719\
        );

    \I__10430\ : InMux
    port map (
            O => \N__45724\,
            I => \N__45719\
        );

    \I__10429\ : LocalMux
    port map (
            O => \N__45719\,
            I => \N__45715\
        );

    \I__10428\ : InMux
    port map (
            O => \N__45718\,
            I => \N__45712\
        );

    \I__10427\ : Span4Mux_v
    port map (
            O => \N__45715\,
            I => \N__45709\
        );

    \I__10426\ : LocalMux
    port map (
            O => \N__45712\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__10425\ : Odrv4
    port map (
            O => \N__45709\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__10424\ : InMux
    port map (
            O => \N__45704\,
            I => \current_shift_inst.timer_s1.counter_cry_2\
        );

    \I__10423\ : CascadeMux
    port map (
            O => \N__45701\,
            I => \N__45698\
        );

    \I__10422\ : InMux
    port map (
            O => \N__45698\,
            I => \N__45694\
        );

    \I__10421\ : InMux
    port map (
            O => \N__45697\,
            I => \N__45691\
        );

    \I__10420\ : LocalMux
    port map (
            O => \N__45694\,
            I => \N__45685\
        );

    \I__10419\ : LocalMux
    port map (
            O => \N__45691\,
            I => \N__45685\
        );

    \I__10418\ : InMux
    port map (
            O => \N__45690\,
            I => \N__45682\
        );

    \I__10417\ : Span4Mux_h
    port map (
            O => \N__45685\,
            I => \N__45679\
        );

    \I__10416\ : LocalMux
    port map (
            O => \N__45682\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__10415\ : Odrv4
    port map (
            O => \N__45679\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__10414\ : InMux
    port map (
            O => \N__45674\,
            I => \current_shift_inst.timer_s1.counter_cry_3\
        );

    \I__10413\ : CascadeMux
    port map (
            O => \N__45671\,
            I => \N__45668\
        );

    \I__10412\ : InMux
    port map (
            O => \N__45668\,
            I => \N__45664\
        );

    \I__10411\ : InMux
    port map (
            O => \N__45667\,
            I => \N__45661\
        );

    \I__10410\ : LocalMux
    port map (
            O => \N__45664\,
            I => \N__45655\
        );

    \I__10409\ : LocalMux
    port map (
            O => \N__45661\,
            I => \N__45655\
        );

    \I__10408\ : InMux
    port map (
            O => \N__45660\,
            I => \N__45652\
        );

    \I__10407\ : Span4Mux_h
    port map (
            O => \N__45655\,
            I => \N__45649\
        );

    \I__10406\ : LocalMux
    port map (
            O => \N__45652\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__10405\ : Odrv4
    port map (
            O => \N__45649\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__10404\ : InMux
    port map (
            O => \N__45644\,
            I => \current_shift_inst.timer_s1.counter_cry_4\
        );

    \I__10403\ : CascadeMux
    port map (
            O => \N__45641\,
            I => \N__45638\
        );

    \I__10402\ : InMux
    port map (
            O => \N__45638\,
            I => \N__45634\
        );

    \I__10401\ : InMux
    port map (
            O => \N__45637\,
            I => \N__45631\
        );

    \I__10400\ : LocalMux
    port map (
            O => \N__45634\,
            I => \N__45625\
        );

    \I__10399\ : LocalMux
    port map (
            O => \N__45631\,
            I => \N__45625\
        );

    \I__10398\ : InMux
    port map (
            O => \N__45630\,
            I => \N__45622\
        );

    \I__10397\ : Span4Mux_h
    port map (
            O => \N__45625\,
            I => \N__45619\
        );

    \I__10396\ : LocalMux
    port map (
            O => \N__45622\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__10395\ : Odrv4
    port map (
            O => \N__45619\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__10394\ : InMux
    port map (
            O => \N__45614\,
            I => \current_shift_inst.timer_s1.counter_cry_5\
        );

    \I__10393\ : CascadeMux
    port map (
            O => \N__45611\,
            I => \N__45608\
        );

    \I__10392\ : InMux
    port map (
            O => \N__45608\,
            I => \N__45604\
        );

    \I__10391\ : InMux
    port map (
            O => \N__45607\,
            I => \N__45601\
        );

    \I__10390\ : LocalMux
    port map (
            O => \N__45604\,
            I => \N__45595\
        );

    \I__10389\ : LocalMux
    port map (
            O => \N__45601\,
            I => \N__45595\
        );

    \I__10388\ : InMux
    port map (
            O => \N__45600\,
            I => \N__45592\
        );

    \I__10387\ : Span4Mux_h
    port map (
            O => \N__45595\,
            I => \N__45589\
        );

    \I__10386\ : LocalMux
    port map (
            O => \N__45592\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__10385\ : Odrv4
    port map (
            O => \N__45589\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__10384\ : InMux
    port map (
            O => \N__45584\,
            I => \current_shift_inst.timer_s1.counter_cry_6\
        );

    \I__10383\ : CascadeMux
    port map (
            O => \N__45581\,
            I => \N__45578\
        );

    \I__10382\ : InMux
    port map (
            O => \N__45578\,
            I => \N__45574\
        );

    \I__10381\ : InMux
    port map (
            O => \N__45577\,
            I => \N__45571\
        );

    \I__10380\ : LocalMux
    port map (
            O => \N__45574\,
            I => \N__45567\
        );

    \I__10379\ : LocalMux
    port map (
            O => \N__45571\,
            I => \N__45564\
        );

    \I__10378\ : InMux
    port map (
            O => \N__45570\,
            I => \N__45561\
        );

    \I__10377\ : Span4Mux_h
    port map (
            O => \N__45567\,
            I => \N__45558\
        );

    \I__10376\ : Span4Mux_h
    port map (
            O => \N__45564\,
            I => \N__45555\
        );

    \I__10375\ : LocalMux
    port map (
            O => \N__45561\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__10374\ : Odrv4
    port map (
            O => \N__45558\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__10373\ : Odrv4
    port map (
            O => \N__45555\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__10372\ : InMux
    port map (
            O => \N__45548\,
            I => \bfn_18_18_0_\
        );

    \I__10371\ : InMux
    port map (
            O => \N__45545\,
            I => \N__45539\
        );

    \I__10370\ : InMux
    port map (
            O => \N__45544\,
            I => \N__45539\
        );

    \I__10369\ : LocalMux
    port map (
            O => \N__45539\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_28\
        );

    \I__10368\ : CascadeMux
    port map (
            O => \N__45536\,
            I => \N__45533\
        );

    \I__10367\ : InMux
    port map (
            O => \N__45533\,
            I => \N__45527\
        );

    \I__10366\ : InMux
    port map (
            O => \N__45532\,
            I => \N__45527\
        );

    \I__10365\ : LocalMux
    port map (
            O => \N__45527\,
            I => \N__45523\
        );

    \I__10364\ : InMux
    port map (
            O => \N__45526\,
            I => \N__45520\
        );

    \I__10363\ : Span4Mux_h
    port map (
            O => \N__45523\,
            I => \N__45517\
        );

    \I__10362\ : LocalMux
    port map (
            O => \N__45520\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__10361\ : Odrv4
    port map (
            O => \N__45517\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__10360\ : InMux
    port map (
            O => \N__45512\,
            I => \N__45506\
        );

    \I__10359\ : InMux
    port map (
            O => \N__45511\,
            I => \N__45506\
        );

    \I__10358\ : LocalMux
    port map (
            O => \N__45506\,
            I => \N__45502\
        );

    \I__10357\ : InMux
    port map (
            O => \N__45505\,
            I => \N__45499\
        );

    \I__10356\ : Span12Mux_v
    port map (
            O => \N__45502\,
            I => \N__45496\
        );

    \I__10355\ : LocalMux
    port map (
            O => \N__45499\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__10354\ : Odrv12
    port map (
            O => \N__45496\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__10353\ : InMux
    port map (
            O => \N__45491\,
            I => \N__45488\
        );

    \I__10352\ : LocalMux
    port map (
            O => \N__45488\,
            I => \N__45485\
        );

    \I__10351\ : Odrv4
    port map (
            O => \N__45485\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt28\
        );

    \I__10350\ : CascadeMux
    port map (
            O => \N__45482\,
            I => \N__45477\
        );

    \I__10349\ : InMux
    port map (
            O => \N__45481\,
            I => \N__45474\
        );

    \I__10348\ : InMux
    port map (
            O => \N__45480\,
            I => \N__45471\
        );

    \I__10347\ : InMux
    port map (
            O => \N__45477\,
            I => \N__45468\
        );

    \I__10346\ : LocalMux
    port map (
            O => \N__45474\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__10345\ : LocalMux
    port map (
            O => \N__45471\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__10344\ : LocalMux
    port map (
            O => \N__45468\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__10343\ : InMux
    port map (
            O => \N__45461\,
            I => \N__45458\
        );

    \I__10342\ : LocalMux
    port map (
            O => \N__45458\,
            I => \current_shift_inst.un4_control_input1_1\
        );

    \I__10341\ : InMux
    port map (
            O => \N__45455\,
            I => \N__45426\
        );

    \I__10340\ : InMux
    port map (
            O => \N__45454\,
            I => \N__45426\
        );

    \I__10339\ : InMux
    port map (
            O => \N__45453\,
            I => \N__45419\
        );

    \I__10338\ : InMux
    port map (
            O => \N__45452\,
            I => \N__45419\
        );

    \I__10337\ : CascadeMux
    port map (
            O => \N__45451\,
            I => \N__45411\
        );

    \I__10336\ : InMux
    port map (
            O => \N__45450\,
            I => \N__45401\
        );

    \I__10335\ : CascadeMux
    port map (
            O => \N__45449\,
            I => \N__45393\
        );

    \I__10334\ : CascadeMux
    port map (
            O => \N__45448\,
            I => \N__45387\
        );

    \I__10333\ : CascadeMux
    port map (
            O => \N__45447\,
            I => \N__45379\
        );

    \I__10332\ : InMux
    port map (
            O => \N__45446\,
            I => \N__45369\
        );

    \I__10331\ : InMux
    port map (
            O => \N__45445\,
            I => \N__45369\
        );

    \I__10330\ : InMux
    port map (
            O => \N__45444\,
            I => \N__45369\
        );

    \I__10329\ : InMux
    port map (
            O => \N__45443\,
            I => \N__45362\
        );

    \I__10328\ : InMux
    port map (
            O => \N__45442\,
            I => \N__45362\
        );

    \I__10327\ : InMux
    port map (
            O => \N__45441\,
            I => \N__45362\
        );

    \I__10326\ : InMux
    port map (
            O => \N__45440\,
            I => \N__45359\
        );

    \I__10325\ : InMux
    port map (
            O => \N__45439\,
            I => \N__45352\
        );

    \I__10324\ : InMux
    port map (
            O => \N__45438\,
            I => \N__45352\
        );

    \I__10323\ : InMux
    port map (
            O => \N__45437\,
            I => \N__45352\
        );

    \I__10322\ : InMux
    port map (
            O => \N__45436\,
            I => \N__45339\
        );

    \I__10321\ : InMux
    port map (
            O => \N__45435\,
            I => \N__45339\
        );

    \I__10320\ : InMux
    port map (
            O => \N__45434\,
            I => \N__45339\
        );

    \I__10319\ : InMux
    port map (
            O => \N__45433\,
            I => \N__45339\
        );

    \I__10318\ : InMux
    port map (
            O => \N__45432\,
            I => \N__45339\
        );

    \I__10317\ : InMux
    port map (
            O => \N__45431\,
            I => \N__45339\
        );

    \I__10316\ : LocalMux
    port map (
            O => \N__45426\,
            I => \N__45336\
        );

    \I__10315\ : InMux
    port map (
            O => \N__45425\,
            I => \N__45330\
        );

    \I__10314\ : InMux
    port map (
            O => \N__45424\,
            I => \N__45330\
        );

    \I__10313\ : LocalMux
    port map (
            O => \N__45419\,
            I => \N__45327\
        );

    \I__10312\ : InMux
    port map (
            O => \N__45418\,
            I => \N__45324\
        );

    \I__10311\ : InMux
    port map (
            O => \N__45417\,
            I => \N__45319\
        );

    \I__10310\ : InMux
    port map (
            O => \N__45416\,
            I => \N__45319\
        );

    \I__10309\ : InMux
    port map (
            O => \N__45415\,
            I => \N__45304\
        );

    \I__10308\ : InMux
    port map (
            O => \N__45414\,
            I => \N__45304\
        );

    \I__10307\ : InMux
    port map (
            O => \N__45411\,
            I => \N__45304\
        );

    \I__10306\ : InMux
    port map (
            O => \N__45410\,
            I => \N__45304\
        );

    \I__10305\ : InMux
    port map (
            O => \N__45409\,
            I => \N__45304\
        );

    \I__10304\ : InMux
    port map (
            O => \N__45408\,
            I => \N__45304\
        );

    \I__10303\ : InMux
    port map (
            O => \N__45407\,
            I => \N__45304\
        );

    \I__10302\ : InMux
    port map (
            O => \N__45406\,
            I => \N__45297\
        );

    \I__10301\ : InMux
    port map (
            O => \N__45405\,
            I => \N__45297\
        );

    \I__10300\ : InMux
    port map (
            O => \N__45404\,
            I => \N__45297\
        );

    \I__10299\ : LocalMux
    port map (
            O => \N__45401\,
            I => \N__45294\
        );

    \I__10298\ : InMux
    port map (
            O => \N__45400\,
            I => \N__45285\
        );

    \I__10297\ : InMux
    port map (
            O => \N__45399\,
            I => \N__45285\
        );

    \I__10296\ : InMux
    port map (
            O => \N__45398\,
            I => \N__45285\
        );

    \I__10295\ : InMux
    port map (
            O => \N__45397\,
            I => \N__45285\
        );

    \I__10294\ : InMux
    port map (
            O => \N__45396\,
            I => \N__45262\
        );

    \I__10293\ : InMux
    port map (
            O => \N__45393\,
            I => \N__45262\
        );

    \I__10292\ : InMux
    port map (
            O => \N__45392\,
            I => \N__45262\
        );

    \I__10291\ : InMux
    port map (
            O => \N__45391\,
            I => \N__45262\
        );

    \I__10290\ : InMux
    port map (
            O => \N__45390\,
            I => \N__45262\
        );

    \I__10289\ : InMux
    port map (
            O => \N__45387\,
            I => \N__45262\
        );

    \I__10288\ : InMux
    port map (
            O => \N__45386\,
            I => \N__45262\
        );

    \I__10287\ : InMux
    port map (
            O => \N__45385\,
            I => \N__45247\
        );

    \I__10286\ : InMux
    port map (
            O => \N__45384\,
            I => \N__45247\
        );

    \I__10285\ : InMux
    port map (
            O => \N__45383\,
            I => \N__45247\
        );

    \I__10284\ : InMux
    port map (
            O => \N__45382\,
            I => \N__45247\
        );

    \I__10283\ : InMux
    port map (
            O => \N__45379\,
            I => \N__45247\
        );

    \I__10282\ : InMux
    port map (
            O => \N__45378\,
            I => \N__45247\
        );

    \I__10281\ : InMux
    port map (
            O => \N__45377\,
            I => \N__45247\
        );

    \I__10280\ : InMux
    port map (
            O => \N__45376\,
            I => \N__45244\
        );

    \I__10279\ : LocalMux
    port map (
            O => \N__45369\,
            I => \N__45241\
        );

    \I__10278\ : LocalMux
    port map (
            O => \N__45362\,
            I => \N__45236\
        );

    \I__10277\ : LocalMux
    port map (
            O => \N__45359\,
            I => \N__45236\
        );

    \I__10276\ : LocalMux
    port map (
            O => \N__45352\,
            I => \N__45233\
        );

    \I__10275\ : LocalMux
    port map (
            O => \N__45339\,
            I => \N__45228\
        );

    \I__10274\ : Span4Mux_h
    port map (
            O => \N__45336\,
            I => \N__45228\
        );

    \I__10273\ : InMux
    port map (
            O => \N__45335\,
            I => \N__45225\
        );

    \I__10272\ : LocalMux
    port map (
            O => \N__45330\,
            I => \N__45209\
        );

    \I__10271\ : Span4Mux_v
    port map (
            O => \N__45327\,
            I => \N__45209\
        );

    \I__10270\ : LocalMux
    port map (
            O => \N__45324\,
            I => \N__45209\
        );

    \I__10269\ : LocalMux
    port map (
            O => \N__45319\,
            I => \N__45209\
        );

    \I__10268\ : LocalMux
    port map (
            O => \N__45304\,
            I => \N__45206\
        );

    \I__10267\ : LocalMux
    port map (
            O => \N__45297\,
            I => \N__45203\
        );

    \I__10266\ : Span4Mux_h
    port map (
            O => \N__45294\,
            I => \N__45198\
        );

    \I__10265\ : LocalMux
    port map (
            O => \N__45285\,
            I => \N__45198\
        );

    \I__10264\ : InMux
    port map (
            O => \N__45284\,
            I => \N__45195\
        );

    \I__10263\ : InMux
    port map (
            O => \N__45283\,
            I => \N__45190\
        );

    \I__10262\ : InMux
    port map (
            O => \N__45282\,
            I => \N__45190\
        );

    \I__10261\ : InMux
    port map (
            O => \N__45281\,
            I => \N__45185\
        );

    \I__10260\ : InMux
    port map (
            O => \N__45280\,
            I => \N__45185\
        );

    \I__10259\ : InMux
    port map (
            O => \N__45279\,
            I => \N__45178\
        );

    \I__10258\ : InMux
    port map (
            O => \N__45278\,
            I => \N__45178\
        );

    \I__10257\ : InMux
    port map (
            O => \N__45277\,
            I => \N__45178\
        );

    \I__10256\ : LocalMux
    port map (
            O => \N__45262\,
            I => \N__45173\
        );

    \I__10255\ : LocalMux
    port map (
            O => \N__45247\,
            I => \N__45173\
        );

    \I__10254\ : LocalMux
    port map (
            O => \N__45244\,
            I => \N__45170\
        );

    \I__10253\ : Span4Mux_h
    port map (
            O => \N__45241\,
            I => \N__45165\
        );

    \I__10252\ : Span4Mux_h
    port map (
            O => \N__45236\,
            I => \N__45165\
        );

    \I__10251\ : Span4Mux_v
    port map (
            O => \N__45233\,
            I => \N__45158\
        );

    \I__10250\ : Span4Mux_v
    port map (
            O => \N__45228\,
            I => \N__45158\
        );

    \I__10249\ : LocalMux
    port map (
            O => \N__45225\,
            I => \N__45158\
        );

    \I__10248\ : InMux
    port map (
            O => \N__45224\,
            I => \N__45151\
        );

    \I__10247\ : InMux
    port map (
            O => \N__45223\,
            I => \N__45151\
        );

    \I__10246\ : InMux
    port map (
            O => \N__45222\,
            I => \N__45151\
        );

    \I__10245\ : InMux
    port map (
            O => \N__45221\,
            I => \N__45142\
        );

    \I__10244\ : InMux
    port map (
            O => \N__45220\,
            I => \N__45142\
        );

    \I__10243\ : InMux
    port map (
            O => \N__45219\,
            I => \N__45142\
        );

    \I__10242\ : InMux
    port map (
            O => \N__45218\,
            I => \N__45142\
        );

    \I__10241\ : Span4Mux_v
    port map (
            O => \N__45209\,
            I => \N__45139\
        );

    \I__10240\ : Span4Mux_v
    port map (
            O => \N__45206\,
            I => \N__45132\
        );

    \I__10239\ : Span4Mux_h
    port map (
            O => \N__45203\,
            I => \N__45132\
        );

    \I__10238\ : Span4Mux_v
    port map (
            O => \N__45198\,
            I => \N__45132\
        );

    \I__10237\ : LocalMux
    port map (
            O => \N__45195\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10236\ : LocalMux
    port map (
            O => \N__45190\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10235\ : LocalMux
    port map (
            O => \N__45185\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10234\ : LocalMux
    port map (
            O => \N__45178\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10233\ : Odrv4
    port map (
            O => \N__45173\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10232\ : Odrv4
    port map (
            O => \N__45170\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10231\ : Odrv4
    port map (
            O => \N__45165\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10230\ : Odrv4
    port map (
            O => \N__45158\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10229\ : LocalMux
    port map (
            O => \N__45151\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10228\ : LocalMux
    port map (
            O => \N__45142\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10227\ : Odrv4
    port map (
            O => \N__45139\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10226\ : Odrv4
    port map (
            O => \N__45132\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10225\ : CascadeMux
    port map (
            O => \N__45107\,
            I => \current_shift_inst.un4_control_input1_1_cascade_\
        );

    \I__10224\ : InMux
    port map (
            O => \N__45104\,
            I => \N__45098\
        );

    \I__10223\ : InMux
    port map (
            O => \N__45103\,
            I => \N__45095\
        );

    \I__10222\ : InMux
    port map (
            O => \N__45102\,
            I => \N__45090\
        );

    \I__10221\ : InMux
    port map (
            O => \N__45101\,
            I => \N__45090\
        );

    \I__10220\ : LocalMux
    port map (
            O => \N__45098\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__10219\ : LocalMux
    port map (
            O => \N__45095\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__10218\ : LocalMux
    port map (
            O => \N__45090\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__10217\ : InMux
    port map (
            O => \N__45083\,
            I => \N__45080\
        );

    \I__10216\ : LocalMux
    port map (
            O => \N__45080\,
            I => \N__45077\
        );

    \I__10215\ : Span4Mux_v
    port map (
            O => \N__45077\,
            I => \N__45073\
        );

    \I__10214\ : InMux
    port map (
            O => \N__45076\,
            I => \N__45070\
        );

    \I__10213\ : Span4Mux_h
    port map (
            O => \N__45073\,
            I => \N__45067\
        );

    \I__10212\ : LocalMux
    port map (
            O => \N__45070\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__10211\ : Odrv4
    port map (
            O => \N__45067\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__10210\ : CascadeMux
    port map (
            O => \N__45062\,
            I => \N__45059\
        );

    \I__10209\ : InMux
    port map (
            O => \N__45059\,
            I => \N__45055\
        );

    \I__10208\ : InMux
    port map (
            O => \N__45058\,
            I => \N__45052\
        );

    \I__10207\ : LocalMux
    port map (
            O => \N__45055\,
            I => \N__45049\
        );

    \I__10206\ : LocalMux
    port map (
            O => \N__45052\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__10205\ : Odrv12
    port map (
            O => \N__45049\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__10204\ : InMux
    port map (
            O => \N__45044\,
            I => \N__45038\
        );

    \I__10203\ : InMux
    port map (
            O => \N__45043\,
            I => \N__45035\
        );

    \I__10202\ : InMux
    port map (
            O => \N__45042\,
            I => \N__45028\
        );

    \I__10201\ : InMux
    port map (
            O => \N__45041\,
            I => \N__45028\
        );

    \I__10200\ : LocalMux
    port map (
            O => \N__45038\,
            I => \N__45023\
        );

    \I__10199\ : LocalMux
    port map (
            O => \N__45035\,
            I => \N__45023\
        );

    \I__10198\ : InMux
    port map (
            O => \N__45034\,
            I => \N__45020\
        );

    \I__10197\ : InMux
    port map (
            O => \N__45033\,
            I => \N__45017\
        );

    \I__10196\ : LocalMux
    port map (
            O => \N__45028\,
            I => \N__45014\
        );

    \I__10195\ : Span4Mux_v
    port map (
            O => \N__45023\,
            I => \N__45011\
        );

    \I__10194\ : LocalMux
    port map (
            O => \N__45020\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__10193\ : LocalMux
    port map (
            O => \N__45017\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__10192\ : Odrv12
    port map (
            O => \N__45014\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__10191\ : Odrv4
    port map (
            O => \N__45011\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__10190\ : InMux
    port map (
            O => \N__45002\,
            I => \N__44998\
        );

    \I__10189\ : InMux
    port map (
            O => \N__45001\,
            I => \N__44994\
        );

    \I__10188\ : LocalMux
    port map (
            O => \N__44998\,
            I => \N__44991\
        );

    \I__10187\ : InMux
    port map (
            O => \N__44997\,
            I => \N__44988\
        );

    \I__10186\ : LocalMux
    port map (
            O => \N__44994\,
            I => \N__44985\
        );

    \I__10185\ : Span4Mux_v
    port map (
            O => \N__44991\,
            I => \N__44982\
        );

    \I__10184\ : LocalMux
    port map (
            O => \N__44988\,
            I => \N__44979\
        );

    \I__10183\ : Span4Mux_v
    port map (
            O => \N__44985\,
            I => \N__44976\
        );

    \I__10182\ : Span4Mux_v
    port map (
            O => \N__44982\,
            I => \N__44971\
        );

    \I__10181\ : Span4Mux_v
    port map (
            O => \N__44979\,
            I => \N__44971\
        );

    \I__10180\ : Odrv4
    port map (
            O => \N__44976\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__10179\ : Odrv4
    port map (
            O => \N__44971\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__10178\ : InMux
    port map (
            O => \N__44966\,
            I => \N__44963\
        );

    \I__10177\ : LocalMux
    port map (
            O => \N__44963\,
            I => \current_shift_inst.elapsed_time_ns_s1_fast_31\
        );

    \I__10176\ : CEMux
    port map (
            O => \N__44960\,
            I => \N__44936\
        );

    \I__10175\ : CEMux
    port map (
            O => \N__44959\,
            I => \N__44936\
        );

    \I__10174\ : CEMux
    port map (
            O => \N__44958\,
            I => \N__44936\
        );

    \I__10173\ : CEMux
    port map (
            O => \N__44957\,
            I => \N__44936\
        );

    \I__10172\ : CEMux
    port map (
            O => \N__44956\,
            I => \N__44936\
        );

    \I__10171\ : CEMux
    port map (
            O => \N__44955\,
            I => \N__44936\
        );

    \I__10170\ : CEMux
    port map (
            O => \N__44954\,
            I => \N__44936\
        );

    \I__10169\ : CEMux
    port map (
            O => \N__44953\,
            I => \N__44936\
        );

    \I__10168\ : GlobalMux
    port map (
            O => \N__44936\,
            I => \N__44933\
        );

    \I__10167\ : gio2CtrlBuf
    port map (
            O => \N__44933\,
            I => \current_shift_inst.timer_s1.N_162_i_g\
        );

    \I__10166\ : InMux
    port map (
            O => \N__44930\,
            I => \N__44923\
        );

    \I__10165\ : InMux
    port map (
            O => \N__44929\,
            I => \N__44923\
        );

    \I__10164\ : InMux
    port map (
            O => \N__44928\,
            I => \N__44920\
        );

    \I__10163\ : LocalMux
    port map (
            O => \N__44923\,
            I => \N__44917\
        );

    \I__10162\ : LocalMux
    port map (
            O => \N__44920\,
            I => \N__44893\
        );

    \I__10161\ : Span4Mux_v
    port map (
            O => \N__44917\,
            I => \N__44893\
        );

    \I__10160\ : InMux
    port map (
            O => \N__44916\,
            I => \N__44884\
        );

    \I__10159\ : InMux
    port map (
            O => \N__44915\,
            I => \N__44884\
        );

    \I__10158\ : InMux
    port map (
            O => \N__44914\,
            I => \N__44884\
        );

    \I__10157\ : InMux
    port map (
            O => \N__44913\,
            I => \N__44884\
        );

    \I__10156\ : InMux
    port map (
            O => \N__44912\,
            I => \N__44873\
        );

    \I__10155\ : InMux
    port map (
            O => \N__44911\,
            I => \N__44873\
        );

    \I__10154\ : InMux
    port map (
            O => \N__44910\,
            I => \N__44873\
        );

    \I__10153\ : InMux
    port map (
            O => \N__44909\,
            I => \N__44873\
        );

    \I__10152\ : InMux
    port map (
            O => \N__44908\,
            I => \N__44873\
        );

    \I__10151\ : InMux
    port map (
            O => \N__44907\,
            I => \N__44866\
        );

    \I__10150\ : InMux
    port map (
            O => \N__44906\,
            I => \N__44866\
        );

    \I__10149\ : InMux
    port map (
            O => \N__44905\,
            I => \N__44866\
        );

    \I__10148\ : InMux
    port map (
            O => \N__44904\,
            I => \N__44860\
        );

    \I__10147\ : InMux
    port map (
            O => \N__44903\,
            I => \N__44849\
        );

    \I__10146\ : InMux
    port map (
            O => \N__44902\,
            I => \N__44849\
        );

    \I__10145\ : InMux
    port map (
            O => \N__44901\,
            I => \N__44849\
        );

    \I__10144\ : InMux
    port map (
            O => \N__44900\,
            I => \N__44849\
        );

    \I__10143\ : InMux
    port map (
            O => \N__44899\,
            I => \N__44849\
        );

    \I__10142\ : InMux
    port map (
            O => \N__44898\,
            I => \N__44846\
        );

    \I__10141\ : Sp12to4
    port map (
            O => \N__44893\,
            I => \N__44837\
        );

    \I__10140\ : LocalMux
    port map (
            O => \N__44884\,
            I => \N__44837\
        );

    \I__10139\ : LocalMux
    port map (
            O => \N__44873\,
            I => \N__44837\
        );

    \I__10138\ : LocalMux
    port map (
            O => \N__44866\,
            I => \N__44837\
        );

    \I__10137\ : InMux
    port map (
            O => \N__44865\,
            I => \N__44834\
        );

    \I__10136\ : InMux
    port map (
            O => \N__44864\,
            I => \N__44829\
        );

    \I__10135\ : InMux
    port map (
            O => \N__44863\,
            I => \N__44829\
        );

    \I__10134\ : LocalMux
    port map (
            O => \N__44860\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__10133\ : LocalMux
    port map (
            O => \N__44849\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__10132\ : LocalMux
    port map (
            O => \N__44846\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__10131\ : Odrv12
    port map (
            O => \N__44837\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__10130\ : LocalMux
    port map (
            O => \N__44834\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__10129\ : LocalMux
    port map (
            O => \N__44829\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__10128\ : InMux
    port map (
            O => \N__44816\,
            I => \N__44813\
        );

    \I__10127\ : LocalMux
    port map (
            O => \N__44813\,
            I => \N__44808\
        );

    \I__10126\ : InMux
    port map (
            O => \N__44812\,
            I => \N__44805\
        );

    \I__10125\ : InMux
    port map (
            O => \N__44811\,
            I => \N__44802\
        );

    \I__10124\ : Span4Mux_v
    port map (
            O => \N__44808\,
            I => \N__44799\
        );

    \I__10123\ : LocalMux
    port map (
            O => \N__44805\,
            I => \N__44794\
        );

    \I__10122\ : LocalMux
    port map (
            O => \N__44802\,
            I => \N__44794\
        );

    \I__10121\ : Odrv4
    port map (
            O => \N__44799\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__10120\ : Odrv4
    port map (
            O => \N__44794\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__10119\ : InMux
    port map (
            O => \N__44789\,
            I => \N__44786\
        );

    \I__10118\ : LocalMux
    port map (
            O => \N__44786\,
            I => \N__44783\
        );

    \I__10117\ : Span4Mux_v
    port map (
            O => \N__44783\,
            I => \N__44780\
        );

    \I__10116\ : Odrv4
    port map (
            O => \N__44780\,
            I => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\
        );

    \I__10115\ : InMux
    port map (
            O => \N__44777\,
            I => \N__44771\
        );

    \I__10114\ : InMux
    port map (
            O => \N__44776\,
            I => \N__44768\
        );

    \I__10113\ : InMux
    port map (
            O => \N__44775\,
            I => \N__44763\
        );

    \I__10112\ : InMux
    port map (
            O => \N__44774\,
            I => \N__44763\
        );

    \I__10111\ : LocalMux
    port map (
            O => \N__44771\,
            I => \N__44760\
        );

    \I__10110\ : LocalMux
    port map (
            O => \N__44768\,
            I => \N__44757\
        );

    \I__10109\ : LocalMux
    port map (
            O => \N__44763\,
            I => \N__44754\
        );

    \I__10108\ : Span4Mux_h
    port map (
            O => \N__44760\,
            I => \N__44751\
        );

    \I__10107\ : Span4Mux_v
    port map (
            O => \N__44757\,
            I => \N__44746\
        );

    \I__10106\ : Span4Mux_h
    port map (
            O => \N__44754\,
            I => \N__44746\
        );

    \I__10105\ : Odrv4
    port map (
            O => \N__44751\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__10104\ : Odrv4
    port map (
            O => \N__44746\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__10103\ : InMux
    port map (
            O => \N__44741\,
            I => \N__44738\
        );

    \I__10102\ : LocalMux
    port map (
            O => \N__44738\,
            I => \N__44735\
        );

    \I__10101\ : Odrv4
    port map (
            O => \N__44735\,
            I => \current_shift_inst.un4_control_input_1_axb_11\
        );

    \I__10100\ : InMux
    port map (
            O => \N__44732\,
            I => \N__44728\
        );

    \I__10099\ : InMux
    port map (
            O => \N__44731\,
            I => \N__44725\
        );

    \I__10098\ : LocalMux
    port map (
            O => \N__44728\,
            I => \N__44721\
        );

    \I__10097\ : LocalMux
    port map (
            O => \N__44725\,
            I => \N__44718\
        );

    \I__10096\ : InMux
    port map (
            O => \N__44724\,
            I => \N__44715\
        );

    \I__10095\ : Span4Mux_h
    port map (
            O => \N__44721\,
            I => \N__44712\
        );

    \I__10094\ : Odrv4
    port map (
            O => \N__44718\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__10093\ : LocalMux
    port map (
            O => \N__44715\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__10092\ : Odrv4
    port map (
            O => \N__44712\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__10091\ : InMux
    port map (
            O => \N__44705\,
            I => \bfn_18_17_0_\
        );

    \I__10090\ : InMux
    port map (
            O => \N__44702\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\
        );

    \I__10089\ : InMux
    port map (
            O => \N__44699\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\
        );

    \I__10088\ : InMux
    port map (
            O => \N__44696\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\
        );

    \I__10087\ : CascadeMux
    port map (
            O => \N__44693\,
            I => \N__44689\
        );

    \I__10086\ : CascadeMux
    port map (
            O => \N__44692\,
            I => \N__44686\
        );

    \I__10085\ : InMux
    port map (
            O => \N__44689\,
            I => \N__44681\
        );

    \I__10084\ : InMux
    port map (
            O => \N__44686\,
            I => \N__44681\
        );

    \I__10083\ : LocalMux
    port map (
            O => \N__44681\,
            I => \N__44677\
        );

    \I__10082\ : InMux
    port map (
            O => \N__44680\,
            I => \N__44674\
        );

    \I__10081\ : Span4Mux_v
    port map (
            O => \N__44677\,
            I => \N__44671\
        );

    \I__10080\ : LocalMux
    port map (
            O => \N__44674\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__10079\ : Odrv4
    port map (
            O => \N__44671\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__10078\ : InMux
    port map (
            O => \N__44666\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\
        );

    \I__10077\ : InMux
    port map (
            O => \N__44663\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\
        );

    \I__10076\ : InMux
    port map (
            O => \N__44660\,
            I => \N__44654\
        );

    \I__10075\ : InMux
    port map (
            O => \N__44659\,
            I => \N__44654\
        );

    \I__10074\ : LocalMux
    port map (
            O => \N__44654\,
            I => \N__44650\
        );

    \I__10073\ : InMux
    port map (
            O => \N__44653\,
            I => \N__44647\
        );

    \I__10072\ : Span4Mux_v
    port map (
            O => \N__44650\,
            I => \N__44644\
        );

    \I__10071\ : LocalMux
    port map (
            O => \N__44647\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__10070\ : Odrv4
    port map (
            O => \N__44644\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__10069\ : CascadeMux
    port map (
            O => \N__44639\,
            I => \N__44636\
        );

    \I__10068\ : InMux
    port map (
            O => \N__44636\,
            I => \N__44633\
        );

    \I__10067\ : LocalMux
    port map (
            O => \N__44633\,
            I => \N__44630\
        );

    \I__10066\ : Span4Mux_h
    port map (
            O => \N__44630\,
            I => \N__44627\
        );

    \I__10065\ : Odrv4
    port map (
            O => \N__44627\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt26\
        );

    \I__10064\ : CascadeMux
    port map (
            O => \N__44624\,
            I => \N__44620\
        );

    \I__10063\ : InMux
    port map (
            O => \N__44623\,
            I => \N__44615\
        );

    \I__10062\ : InMux
    port map (
            O => \N__44620\,
            I => \N__44615\
        );

    \I__10061\ : LocalMux
    port map (
            O => \N__44615\,
            I => \N__44611\
        );

    \I__10060\ : InMux
    port map (
            O => \N__44614\,
            I => \N__44608\
        );

    \I__10059\ : Span4Mux_v
    port map (
            O => \N__44611\,
            I => \N__44605\
        );

    \I__10058\ : LocalMux
    port map (
            O => \N__44608\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__10057\ : Odrv4
    port map (
            O => \N__44605\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__10056\ : CascadeMux
    port map (
            O => \N__44600\,
            I => \N__44597\
        );

    \I__10055\ : InMux
    port map (
            O => \N__44597\,
            I => \N__44593\
        );

    \I__10054\ : InMux
    port map (
            O => \N__44596\,
            I => \N__44590\
        );

    \I__10053\ : LocalMux
    port map (
            O => \N__44593\,
            I => \N__44584\
        );

    \I__10052\ : LocalMux
    port map (
            O => \N__44590\,
            I => \N__44584\
        );

    \I__10051\ : InMux
    port map (
            O => \N__44589\,
            I => \N__44581\
        );

    \I__10050\ : Span4Mux_v
    port map (
            O => \N__44584\,
            I => \N__44578\
        );

    \I__10049\ : LocalMux
    port map (
            O => \N__44581\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__10048\ : Odrv4
    port map (
            O => \N__44578\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__10047\ : InMux
    port map (
            O => \N__44573\,
            I => \N__44570\
        );

    \I__10046\ : LocalMux
    port map (
            O => \N__44570\,
            I => \N__44567\
        );

    \I__10045\ : Odrv12
    port map (
            O => \N__44567\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26\
        );

    \I__10044\ : CascadeMux
    port map (
            O => \N__44564\,
            I => \N__44561\
        );

    \I__10043\ : InMux
    port map (
            O => \N__44561\,
            I => \N__44558\
        );

    \I__10042\ : LocalMux
    port map (
            O => \N__44558\,
            I => \N__44555\
        );

    \I__10041\ : Odrv4
    port map (
            O => \N__44555\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28\
        );

    \I__10040\ : CascadeMux
    port map (
            O => \N__44552\,
            I => \N__44549\
        );

    \I__10039\ : InMux
    port map (
            O => \N__44549\,
            I => \N__44542\
        );

    \I__10038\ : InMux
    port map (
            O => \N__44548\,
            I => \N__44542\
        );

    \I__10037\ : InMux
    port map (
            O => \N__44547\,
            I => \N__44539\
        );

    \I__10036\ : LocalMux
    port map (
            O => \N__44542\,
            I => \N__44536\
        );

    \I__10035\ : LocalMux
    port map (
            O => \N__44539\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__10034\ : Odrv12
    port map (
            O => \N__44536\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__10033\ : InMux
    port map (
            O => \N__44531\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\
        );

    \I__10032\ : InMux
    port map (
            O => \N__44528\,
            I => \N__44521\
        );

    \I__10031\ : InMux
    port map (
            O => \N__44527\,
            I => \N__44521\
        );

    \I__10030\ : InMux
    port map (
            O => \N__44526\,
            I => \N__44518\
        );

    \I__10029\ : LocalMux
    port map (
            O => \N__44521\,
            I => \N__44515\
        );

    \I__10028\ : LocalMux
    port map (
            O => \N__44518\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__10027\ : Odrv12
    port map (
            O => \N__44515\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__10026\ : InMux
    port map (
            O => \N__44510\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\
        );

    \I__10025\ : CascadeMux
    port map (
            O => \N__44507\,
            I => \N__44503\
        );

    \I__10024\ : InMux
    port map (
            O => \N__44506\,
            I => \N__44497\
        );

    \I__10023\ : InMux
    port map (
            O => \N__44503\,
            I => \N__44497\
        );

    \I__10022\ : InMux
    port map (
            O => \N__44502\,
            I => \N__44494\
        );

    \I__10021\ : LocalMux
    port map (
            O => \N__44497\,
            I => \N__44491\
        );

    \I__10020\ : LocalMux
    port map (
            O => \N__44494\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__10019\ : Odrv12
    port map (
            O => \N__44491\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__10018\ : InMux
    port map (
            O => \N__44486\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\
        );

    \I__10017\ : CascadeMux
    port map (
            O => \N__44483\,
            I => \N__44480\
        );

    \I__10016\ : InMux
    port map (
            O => \N__44480\,
            I => \N__44475\
        );

    \I__10015\ : InMux
    port map (
            O => \N__44479\,
            I => \N__44472\
        );

    \I__10014\ : InMux
    port map (
            O => \N__44478\,
            I => \N__44469\
        );

    \I__10013\ : LocalMux
    port map (
            O => \N__44475\,
            I => \N__44464\
        );

    \I__10012\ : LocalMux
    port map (
            O => \N__44472\,
            I => \N__44464\
        );

    \I__10011\ : LocalMux
    port map (
            O => \N__44469\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__10010\ : Odrv12
    port map (
            O => \N__44464\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__10009\ : InMux
    port map (
            O => \N__44459\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__10008\ : InMux
    port map (
            O => \N__44456\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\
        );

    \I__10007\ : InMux
    port map (
            O => \N__44453\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\
        );

    \I__10006\ : InMux
    port map (
            O => \N__44450\,
            I => \N__44445\
        );

    \I__10005\ : InMux
    port map (
            O => \N__44449\,
            I => \N__44440\
        );

    \I__10004\ : InMux
    port map (
            O => \N__44448\,
            I => \N__44440\
        );

    \I__10003\ : LocalMux
    port map (
            O => \N__44445\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__10002\ : LocalMux
    port map (
            O => \N__44440\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__10001\ : InMux
    port map (
            O => \N__44435\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\
        );

    \I__10000\ : CascadeMux
    port map (
            O => \N__44432\,
            I => \N__44427\
        );

    \I__9999\ : InMux
    port map (
            O => \N__44431\,
            I => \N__44424\
        );

    \I__9998\ : InMux
    port map (
            O => \N__44430\,
            I => \N__44419\
        );

    \I__9997\ : InMux
    port map (
            O => \N__44427\,
            I => \N__44419\
        );

    \I__9996\ : LocalMux
    port map (
            O => \N__44424\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__9995\ : LocalMux
    port map (
            O => \N__44419\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__9994\ : InMux
    port map (
            O => \N__44414\,
            I => \bfn_18_14_0_\
        );

    \I__9993\ : InMux
    port map (
            O => \N__44411\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\
        );

    \I__9992\ : InMux
    port map (
            O => \N__44408\,
            I => \N__44404\
        );

    \I__9991\ : InMux
    port map (
            O => \N__44407\,
            I => \N__44401\
        );

    \I__9990\ : LocalMux
    port map (
            O => \N__44404\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__9989\ : LocalMux
    port map (
            O => \N__44401\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__9988\ : InMux
    port map (
            O => \N__44396\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\
        );

    \I__9987\ : InMux
    port map (
            O => \N__44393\,
            I => \N__44389\
        );

    \I__9986\ : InMux
    port map (
            O => \N__44392\,
            I => \N__44386\
        );

    \I__9985\ : LocalMux
    port map (
            O => \N__44389\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__9984\ : LocalMux
    port map (
            O => \N__44386\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__9983\ : InMux
    port map (
            O => \N__44381\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\
        );

    \I__9982\ : InMux
    port map (
            O => \N__44378\,
            I => \N__44375\
        );

    \I__9981\ : LocalMux
    port map (
            O => \N__44375\,
            I => \N__44371\
        );

    \I__9980\ : InMux
    port map (
            O => \N__44374\,
            I => \N__44368\
        );

    \I__9979\ : Span4Mux_h
    port map (
            O => \N__44371\,
            I => \N__44365\
        );

    \I__9978\ : LocalMux
    port map (
            O => \N__44368\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__9977\ : Odrv4
    port map (
            O => \N__44365\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__9976\ : InMux
    port map (
            O => \N__44360\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\
        );

    \I__9975\ : InMux
    port map (
            O => \N__44357\,
            I => \N__44353\
        );

    \I__9974\ : InMux
    port map (
            O => \N__44356\,
            I => \N__44350\
        );

    \I__9973\ : LocalMux
    port map (
            O => \N__44353\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__9972\ : LocalMux
    port map (
            O => \N__44350\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__9971\ : InMux
    port map (
            O => \N__44345\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\
        );

    \I__9970\ : InMux
    port map (
            O => \N__44342\,
            I => \N__44338\
        );

    \I__9969\ : InMux
    port map (
            O => \N__44341\,
            I => \N__44335\
        );

    \I__9968\ : LocalMux
    port map (
            O => \N__44338\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__9967\ : LocalMux
    port map (
            O => \N__44335\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__9966\ : InMux
    port map (
            O => \N__44330\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\
        );

    \I__9965\ : InMux
    port map (
            O => \N__44327\,
            I => \N__44323\
        );

    \I__9964\ : InMux
    port map (
            O => \N__44326\,
            I => \N__44320\
        );

    \I__9963\ : LocalMux
    port map (
            O => \N__44323\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__9962\ : LocalMux
    port map (
            O => \N__44320\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__9961\ : InMux
    port map (
            O => \N__44315\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\
        );

    \I__9960\ : InMux
    port map (
            O => \N__44312\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\
        );

    \I__9959\ : InMux
    port map (
            O => \N__44309\,
            I => \bfn_18_13_0_\
        );

    \I__9958\ : InMux
    port map (
            O => \N__44306\,
            I => \N__44303\
        );

    \I__9957\ : LocalMux
    port map (
            O => \N__44303\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\
        );

    \I__9956\ : CascadeMux
    port map (
            O => \N__44300\,
            I => \N__44297\
        );

    \I__9955\ : InMux
    port map (
            O => \N__44297\,
            I => \N__44293\
        );

    \I__9954\ : CascadeMux
    port map (
            O => \N__44296\,
            I => \N__44289\
        );

    \I__9953\ : LocalMux
    port map (
            O => \N__44293\,
            I => \N__44286\
        );

    \I__9952\ : InMux
    port map (
            O => \N__44292\,
            I => \N__44283\
        );

    \I__9951\ : InMux
    port map (
            O => \N__44289\,
            I => \N__44280\
        );

    \I__9950\ : Span12Mux_h
    port map (
            O => \N__44286\,
            I => \N__44277\
        );

    \I__9949\ : LocalMux
    port map (
            O => \N__44283\,
            I => \N__44274\
        );

    \I__9948\ : LocalMux
    port map (
            O => \N__44280\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__9947\ : Odrv12
    port map (
            O => \N__44277\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__9946\ : Odrv12
    port map (
            O => \N__44274\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__9945\ : InMux
    port map (
            O => \N__44267\,
            I => \N__44263\
        );

    \I__9944\ : InMux
    port map (
            O => \N__44266\,
            I => \N__44260\
        );

    \I__9943\ : LocalMux
    port map (
            O => \N__44263\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__9942\ : LocalMux
    port map (
            O => \N__44260\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__9941\ : InMux
    port map (
            O => \N__44255\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\
        );

    \I__9940\ : CascadeMux
    port map (
            O => \N__44252\,
            I => \N__44249\
        );

    \I__9939\ : InMux
    port map (
            O => \N__44249\,
            I => \N__44246\
        );

    \I__9938\ : LocalMux
    port map (
            O => \N__44246\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1Z0Z_30\
        );

    \I__9937\ : InMux
    port map (
            O => \N__44243\,
            I => \N__44239\
        );

    \I__9936\ : InMux
    port map (
            O => \N__44242\,
            I => \N__44236\
        );

    \I__9935\ : LocalMux
    port map (
            O => \N__44239\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__9934\ : LocalMux
    port map (
            O => \N__44236\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__9933\ : InMux
    port map (
            O => \N__44231\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\
        );

    \I__9932\ : InMux
    port map (
            O => \N__44228\,
            I => \N__44224\
        );

    \I__9931\ : InMux
    port map (
            O => \N__44227\,
            I => \N__44221\
        );

    \I__9930\ : LocalMux
    port map (
            O => \N__44224\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__9929\ : LocalMux
    port map (
            O => \N__44221\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__9928\ : InMux
    port map (
            O => \N__44216\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\
        );

    \I__9927\ : InMux
    port map (
            O => \N__44213\,
            I => \N__44209\
        );

    \I__9926\ : InMux
    port map (
            O => \N__44212\,
            I => \N__44206\
        );

    \I__9925\ : LocalMux
    port map (
            O => \N__44209\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__9924\ : LocalMux
    port map (
            O => \N__44206\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__9923\ : InMux
    port map (
            O => \N__44201\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\
        );

    \I__9922\ : InMux
    port map (
            O => \N__44198\,
            I => \N__44194\
        );

    \I__9921\ : InMux
    port map (
            O => \N__44197\,
            I => \N__44191\
        );

    \I__9920\ : LocalMux
    port map (
            O => \N__44194\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__9919\ : LocalMux
    port map (
            O => \N__44191\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__9918\ : InMux
    port map (
            O => \N__44186\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\
        );

    \I__9917\ : InMux
    port map (
            O => \N__44183\,
            I => \N__44179\
        );

    \I__9916\ : InMux
    port map (
            O => \N__44182\,
            I => \N__44176\
        );

    \I__9915\ : LocalMux
    port map (
            O => \N__44179\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__9914\ : LocalMux
    port map (
            O => \N__44176\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__9913\ : InMux
    port map (
            O => \N__44171\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\
        );

    \I__9912\ : InMux
    port map (
            O => \N__44168\,
            I => \N__44164\
        );

    \I__9911\ : InMux
    port map (
            O => \N__44167\,
            I => \N__44161\
        );

    \I__9910\ : LocalMux
    port map (
            O => \N__44164\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__9909\ : LocalMux
    port map (
            O => \N__44161\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__9908\ : InMux
    port map (
            O => \N__44156\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\
        );

    \I__9907\ : InMux
    port map (
            O => \N__44153\,
            I => \N__44149\
        );

    \I__9906\ : InMux
    port map (
            O => \N__44152\,
            I => \N__44146\
        );

    \I__9905\ : LocalMux
    port map (
            O => \N__44149\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__9904\ : LocalMux
    port map (
            O => \N__44146\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__9903\ : InMux
    port map (
            O => \N__44141\,
            I => \bfn_18_12_0_\
        );

    \I__9902\ : InMux
    port map (
            O => \N__44138\,
            I => \N__44135\
        );

    \I__9901\ : LocalMux
    port map (
            O => \N__44135\,
            I => \N__44132\
        );

    \I__9900\ : Span4Mux_v
    port map (
            O => \N__44132\,
            I => \N__44129\
        );

    \I__9899\ : Odrv4
    port map (
            O => \N__44129\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\
        );

    \I__9898\ : InMux
    port map (
            O => \N__44126\,
            I => \N__44123\
        );

    \I__9897\ : LocalMux
    port map (
            O => \N__44123\,
            I => \N__44120\
        );

    \I__9896\ : Span4Mux_h
    port map (
            O => \N__44120\,
            I => \N__44116\
        );

    \I__9895\ : InMux
    port map (
            O => \N__44119\,
            I => \N__44113\
        );

    \I__9894\ : Odrv4
    port map (
            O => \N__44116\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19\
        );

    \I__9893\ : LocalMux
    port map (
            O => \N__44113\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19\
        );

    \I__9892\ : CascadeMux
    port map (
            O => \N__44108\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19_cascade_\
        );

    \I__9891\ : InMux
    port map (
            O => \N__44105\,
            I => \N__44100\
        );

    \I__9890\ : InMux
    port map (
            O => \N__44104\,
            I => \N__44095\
        );

    \I__9889\ : InMux
    port map (
            O => \N__44103\,
            I => \N__44095\
        );

    \I__9888\ : LocalMux
    port map (
            O => \N__44100\,
            I => \N__44091\
        );

    \I__9887\ : LocalMux
    port map (
            O => \N__44095\,
            I => \N__44088\
        );

    \I__9886\ : InMux
    port map (
            O => \N__44094\,
            I => \N__44085\
        );

    \I__9885\ : Span4Mux_v
    port map (
            O => \N__44091\,
            I => \N__44080\
        );

    \I__9884\ : Span4Mux_h
    port map (
            O => \N__44088\,
            I => \N__44080\
        );

    \I__9883\ : LocalMux
    port map (
            O => \N__44085\,
            I => \N__44077\
        );

    \I__9882\ : Odrv4
    port map (
            O => \N__44080\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__9881\ : Odrv4
    port map (
            O => \N__44077\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__9880\ : CascadeMux
    port map (
            O => \N__44072\,
            I => \N__44068\
        );

    \I__9879\ : InMux
    port map (
            O => \N__44071\,
            I => \N__44063\
        );

    \I__9878\ : InMux
    port map (
            O => \N__44068\,
            I => \N__44063\
        );

    \I__9877\ : LocalMux
    port map (
            O => \N__44063\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\
        );

    \I__9876\ : InMux
    port map (
            O => \N__44060\,
            I => \N__44056\
        );

    \I__9875\ : InMux
    port map (
            O => \N__44059\,
            I => \N__44052\
        );

    \I__9874\ : LocalMux
    port map (
            O => \N__44056\,
            I => \N__44049\
        );

    \I__9873\ : InMux
    port map (
            O => \N__44055\,
            I => \N__44046\
        );

    \I__9872\ : LocalMux
    port map (
            O => \N__44052\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15\
        );

    \I__9871\ : Odrv12
    port map (
            O => \N__44049\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15\
        );

    \I__9870\ : LocalMux
    port map (
            O => \N__44046\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15\
        );

    \I__9869\ : InMux
    port map (
            O => \N__44039\,
            I => \N__44036\
        );

    \I__9868\ : LocalMux
    port map (
            O => \N__44036\,
            I => \N__44032\
        );

    \I__9867\ : InMux
    port map (
            O => \N__44035\,
            I => \N__44029\
        );

    \I__9866\ : Span4Mux_v
    port map (
            O => \N__44032\,
            I => \N__44022\
        );

    \I__9865\ : LocalMux
    port map (
            O => \N__44029\,
            I => \N__44022\
        );

    \I__9864\ : InMux
    port map (
            O => \N__44028\,
            I => \N__44017\
        );

    \I__9863\ : InMux
    port map (
            O => \N__44027\,
            I => \N__44017\
        );

    \I__9862\ : Odrv4
    port map (
            O => \N__44022\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__9861\ : LocalMux
    port map (
            O => \N__44017\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__9860\ : InMux
    port map (
            O => \N__44012\,
            I => \N__44009\
        );

    \I__9859\ : LocalMux
    port map (
            O => \N__44009\,
            I => \N__44006\
        );

    \I__9858\ : Odrv4
    port map (
            O => \N__44006\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\
        );

    \I__9857\ : InMux
    port map (
            O => \N__44003\,
            I => \N__43997\
        );

    \I__9856\ : InMux
    port map (
            O => \N__44002\,
            I => \N__43997\
        );

    \I__9855\ : LocalMux
    port map (
            O => \N__43997\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\
        );

    \I__9854\ : CascadeMux
    port map (
            O => \N__43994\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_\
        );

    \I__9853\ : InMux
    port map (
            O => \N__43991\,
            I => \N__43988\
        );

    \I__9852\ : LocalMux
    port map (
            O => \N__43988\,
            I => \N__43985\
        );

    \I__9851\ : Span4Mux_h
    port map (
            O => \N__43985\,
            I => \N__43981\
        );

    \I__9850\ : InMux
    port map (
            O => \N__43984\,
            I => \N__43978\
        );

    \I__9849\ : Odrv4
    port map (
            O => \N__43981\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\
        );

    \I__9848\ : LocalMux
    port map (
            O => \N__43978\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\
        );

    \I__9847\ : InMux
    port map (
            O => \N__43973\,
            I => \N__43967\
        );

    \I__9846\ : InMux
    port map (
            O => \N__43972\,
            I => \N__43967\
        );

    \I__9845\ : LocalMux
    port map (
            O => \N__43967\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_20\
        );

    \I__9844\ : InMux
    port map (
            O => \N__43964\,
            I => \N__43960\
        );

    \I__9843\ : InMux
    port map (
            O => \N__43963\,
            I => \N__43957\
        );

    \I__9842\ : LocalMux
    port map (
            O => \N__43960\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_21\
        );

    \I__9841\ : LocalMux
    port map (
            O => \N__43957\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_21\
        );

    \I__9840\ : InMux
    port map (
            O => \N__43952\,
            I => \N__43949\
        );

    \I__9839\ : LocalMux
    port map (
            O => \N__43949\,
            I => \N__43946\
        );

    \I__9838\ : Span4Mux_v
    port map (
            O => \N__43946\,
            I => \N__43943\
        );

    \I__9837\ : Odrv4
    port map (
            O => \N__43943\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20\
        );

    \I__9836\ : InMux
    port map (
            O => \N__43940\,
            I => \N__43935\
        );

    \I__9835\ : InMux
    port map (
            O => \N__43939\,
            I => \N__43932\
        );

    \I__9834\ : CascadeMux
    port map (
            O => \N__43938\,
            I => \N__43929\
        );

    \I__9833\ : LocalMux
    port map (
            O => \N__43935\,
            I => \N__43926\
        );

    \I__9832\ : LocalMux
    port map (
            O => \N__43932\,
            I => \N__43923\
        );

    \I__9831\ : InMux
    port map (
            O => \N__43929\,
            I => \N__43920\
        );

    \I__9830\ : Span4Mux_v
    port map (
            O => \N__43926\,
            I => \N__43916\
        );

    \I__9829\ : Span4Mux_h
    port map (
            O => \N__43923\,
            I => \N__43913\
        );

    \I__9828\ : LocalMux
    port map (
            O => \N__43920\,
            I => \N__43910\
        );

    \I__9827\ : InMux
    port map (
            O => \N__43919\,
            I => \N__43907\
        );

    \I__9826\ : Span4Mux_v
    port map (
            O => \N__43916\,
            I => \N__43904\
        );

    \I__9825\ : Span4Mux_v
    port map (
            O => \N__43913\,
            I => \N__43901\
        );

    \I__9824\ : Span4Mux_h
    port map (
            O => \N__43910\,
            I => \N__43898\
        );

    \I__9823\ : LocalMux
    port map (
            O => \N__43907\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__9822\ : Odrv4
    port map (
            O => \N__43904\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__9821\ : Odrv4
    port map (
            O => \N__43901\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__9820\ : Odrv4
    port map (
            O => \N__43898\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__9819\ : InMux
    port map (
            O => \N__43889\,
            I => \N__43886\
        );

    \I__9818\ : LocalMux
    port map (
            O => \N__43886\,
            I => \N__43882\
        );

    \I__9817\ : InMux
    port map (
            O => \N__43885\,
            I => \N__43878\
        );

    \I__9816\ : Span4Mux_v
    port map (
            O => \N__43882\,
            I => \N__43875\
        );

    \I__9815\ : InMux
    port map (
            O => \N__43881\,
            I => \N__43872\
        );

    \I__9814\ : LocalMux
    port map (
            O => \N__43878\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20\
        );

    \I__9813\ : Odrv4
    port map (
            O => \N__43875\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20\
        );

    \I__9812\ : LocalMux
    port map (
            O => \N__43872\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20\
        );

    \I__9811\ : InMux
    port map (
            O => \N__43865\,
            I => \N__43862\
        );

    \I__9810\ : LocalMux
    port map (
            O => \N__43862\,
            I => \N__43858\
        );

    \I__9809\ : InMux
    port map (
            O => \N__43861\,
            I => \N__43855\
        );

    \I__9808\ : Span4Mux_v
    port map (
            O => \N__43858\,
            I => \N__43851\
        );

    \I__9807\ : LocalMux
    port map (
            O => \N__43855\,
            I => \N__43848\
        );

    \I__9806\ : InMux
    port map (
            O => \N__43854\,
            I => \N__43845\
        );

    \I__9805\ : Odrv4
    port map (
            O => \N__43851\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__9804\ : Odrv12
    port map (
            O => \N__43848\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__9803\ : LocalMux
    port map (
            O => \N__43845\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__9802\ : CascadeMux
    port map (
            O => \N__43838\,
            I => \N__43834\
        );

    \I__9801\ : InMux
    port map (
            O => \N__43837\,
            I => \N__43831\
        );

    \I__9800\ : InMux
    port map (
            O => \N__43834\,
            I => \N__43828\
        );

    \I__9799\ : LocalMux
    port map (
            O => \N__43831\,
            I => \N__43825\
        );

    \I__9798\ : LocalMux
    port map (
            O => \N__43828\,
            I => \N__43821\
        );

    \I__9797\ : Span4Mux_v
    port map (
            O => \N__43825\,
            I => \N__43818\
        );

    \I__9796\ : InMux
    port map (
            O => \N__43824\,
            I => \N__43815\
        );

    \I__9795\ : Span4Mux_v
    port map (
            O => \N__43821\,
            I => \N__43812\
        );

    \I__9794\ : Odrv4
    port map (
            O => \N__43818\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__9793\ : LocalMux
    port map (
            O => \N__43815\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__9792\ : Odrv4
    port map (
            O => \N__43812\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__9791\ : CEMux
    port map (
            O => \N__43805\,
            I => \N__43802\
        );

    \I__9790\ : LocalMux
    port map (
            O => \N__43802\,
            I => \N__43797\
        );

    \I__9789\ : CEMux
    port map (
            O => \N__43801\,
            I => \N__43794\
        );

    \I__9788\ : CEMux
    port map (
            O => \N__43800\,
            I => \N__43789\
        );

    \I__9787\ : Span4Mux_h
    port map (
            O => \N__43797\,
            I => \N__43784\
        );

    \I__9786\ : LocalMux
    port map (
            O => \N__43794\,
            I => \N__43784\
        );

    \I__9785\ : CEMux
    port map (
            O => \N__43793\,
            I => \N__43781\
        );

    \I__9784\ : CEMux
    port map (
            O => \N__43792\,
            I => \N__43778\
        );

    \I__9783\ : LocalMux
    port map (
            O => \N__43789\,
            I => \N__43775\
        );

    \I__9782\ : Span4Mux_v
    port map (
            O => \N__43784\,
            I => \N__43772\
        );

    \I__9781\ : LocalMux
    port map (
            O => \N__43781\,
            I => \N__43769\
        );

    \I__9780\ : LocalMux
    port map (
            O => \N__43778\,
            I => \N__43766\
        );

    \I__9779\ : Span4Mux_h
    port map (
            O => \N__43775\,
            I => \N__43763\
        );

    \I__9778\ : Span4Mux_h
    port map (
            O => \N__43772\,
            I => \N__43758\
        );

    \I__9777\ : Span4Mux_h
    port map (
            O => \N__43769\,
            I => \N__43758\
        );

    \I__9776\ : Span4Mux_h
    port map (
            O => \N__43766\,
            I => \N__43755\
        );

    \I__9775\ : Odrv4
    port map (
            O => \N__43763\,
            I => \delay_measurement_inst.delay_hc_timer.N_198_i\
        );

    \I__9774\ : Odrv4
    port map (
            O => \N__43758\,
            I => \delay_measurement_inst.delay_hc_timer.N_198_i\
        );

    \I__9773\ : Odrv4
    port map (
            O => \N__43755\,
            I => \delay_measurement_inst.delay_hc_timer.N_198_i\
        );

    \I__9772\ : InMux
    port map (
            O => \N__43748\,
            I => \N__43745\
        );

    \I__9771\ : LocalMux
    port map (
            O => \N__43745\,
            I => \N__43741\
        );

    \I__9770\ : InMux
    port map (
            O => \N__43744\,
            I => \N__43737\
        );

    \I__9769\ : Span12Mux_h
    port map (
            O => \N__43741\,
            I => \N__43734\
        );

    \I__9768\ : InMux
    port map (
            O => \N__43740\,
            I => \N__43731\
        );

    \I__9767\ : LocalMux
    port map (
            O => \N__43737\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__9766\ : Odrv12
    port map (
            O => \N__43734\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__9765\ : LocalMux
    port map (
            O => \N__43731\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__9764\ : InMux
    port map (
            O => \N__43724\,
            I => \N__43721\
        );

    \I__9763\ : LocalMux
    port map (
            O => \N__43721\,
            I => \N__43717\
        );

    \I__9762\ : InMux
    port map (
            O => \N__43720\,
            I => \N__43713\
        );

    \I__9761\ : Span4Mux_v
    port map (
            O => \N__43717\,
            I => \N__43710\
        );

    \I__9760\ : InMux
    port map (
            O => \N__43716\,
            I => \N__43707\
        );

    \I__9759\ : LocalMux
    port map (
            O => \N__43713\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3\
        );

    \I__9758\ : Odrv4
    port map (
            O => \N__43710\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3\
        );

    \I__9757\ : LocalMux
    port map (
            O => \N__43707\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3\
        );

    \I__9756\ : InMux
    port map (
            O => \N__43700\,
            I => \N__43697\
        );

    \I__9755\ : LocalMux
    port map (
            O => \N__43697\,
            I => \N__43693\
        );

    \I__9754\ : InMux
    port map (
            O => \N__43696\,
            I => \N__43689\
        );

    \I__9753\ : Span4Mux_v
    port map (
            O => \N__43693\,
            I => \N__43686\
        );

    \I__9752\ : InMux
    port map (
            O => \N__43692\,
            I => \N__43683\
        );

    \I__9751\ : LocalMux
    port map (
            O => \N__43689\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4\
        );

    \I__9750\ : Odrv4
    port map (
            O => \N__43686\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4\
        );

    \I__9749\ : LocalMux
    port map (
            O => \N__43683\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4\
        );

    \I__9748\ : CascadeMux
    port map (
            O => \N__43676\,
            I => \N__43673\
        );

    \I__9747\ : InMux
    port map (
            O => \N__43673\,
            I => \N__43670\
        );

    \I__9746\ : LocalMux
    port map (
            O => \N__43670\,
            I => \N__43667\
        );

    \I__9745\ : Span4Mux_v
    port map (
            O => \N__43667\,
            I => \N__43664\
        );

    \I__9744\ : Odrv4
    port map (
            O => \N__43664\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt18\
        );

    \I__9743\ : InMux
    port map (
            O => \N__43661\,
            I => \N__43658\
        );

    \I__9742\ : LocalMux
    port map (
            O => \N__43658\,
            I => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\
        );

    \I__9741\ : CascadeMux
    port map (
            O => \N__43655\,
            I => \N__43652\
        );

    \I__9740\ : InMux
    port map (
            O => \N__43652\,
            I => \N__43649\
        );

    \I__9739\ : LocalMux
    port map (
            O => \N__43649\,
            I => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\
        );

    \I__9738\ : InMux
    port map (
            O => \N__43646\,
            I => \N__43643\
        );

    \I__9737\ : LocalMux
    port map (
            O => \N__43643\,
            I => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\
        );

    \I__9736\ : CascadeMux
    port map (
            O => \N__43640\,
            I => \N__43637\
        );

    \I__9735\ : InMux
    port map (
            O => \N__43637\,
            I => \N__43634\
        );

    \I__9734\ : LocalMux
    port map (
            O => \N__43634\,
            I => \N__43631\
        );

    \I__9733\ : Span4Mux_h
    port map (
            O => \N__43631\,
            I => \N__43628\
        );

    \I__9732\ : Span4Mux_v
    port map (
            O => \N__43628\,
            I => \N__43625\
        );

    \I__9731\ : Odrv4
    port map (
            O => \N__43625\,
            I => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\
        );

    \I__9730\ : InMux
    port map (
            O => \N__43622\,
            I => \N__43619\
        );

    \I__9729\ : LocalMux
    port map (
            O => \N__43619\,
            I => \N__43616\
        );

    \I__9728\ : Span4Mux_v
    port map (
            O => \N__43616\,
            I => \N__43613\
        );

    \I__9727\ : Odrv4
    port map (
            O => \N__43613\,
            I => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\
        );

    \I__9726\ : CascadeMux
    port map (
            O => \N__43610\,
            I => \N__43607\
        );

    \I__9725\ : InMux
    port map (
            O => \N__43607\,
            I => \N__43604\
        );

    \I__9724\ : LocalMux
    port map (
            O => \N__43604\,
            I => \N__43601\
        );

    \I__9723\ : Span12Mux_s11_v
    port map (
            O => \N__43601\,
            I => \N__43598\
        );

    \I__9722\ : Odrv12
    port map (
            O => \N__43598\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\
        );

    \I__9721\ : InMux
    port map (
            O => \N__43595\,
            I => \current_shift_inst.un10_control_input_cry_30\
        );

    \I__9720\ : InMux
    port map (
            O => \N__43592\,
            I => \N__43586\
        );

    \I__9719\ : InMux
    port map (
            O => \N__43591\,
            I => \N__43583\
        );

    \I__9718\ : CascadeMux
    port map (
            O => \N__43590\,
            I => \N__43568\
        );

    \I__9717\ : CascadeMux
    port map (
            O => \N__43589\,
            I => \N__43563\
        );

    \I__9716\ : LocalMux
    port map (
            O => \N__43586\,
            I => \N__43546\
        );

    \I__9715\ : LocalMux
    port map (
            O => \N__43583\,
            I => \N__43546\
        );

    \I__9714\ : InMux
    port map (
            O => \N__43582\,
            I => \N__43543\
        );

    \I__9713\ : InMux
    port map (
            O => \N__43581\,
            I => \N__43532\
        );

    \I__9712\ : InMux
    port map (
            O => \N__43580\,
            I => \N__43532\
        );

    \I__9711\ : InMux
    port map (
            O => \N__43579\,
            I => \N__43532\
        );

    \I__9710\ : InMux
    port map (
            O => \N__43578\,
            I => \N__43532\
        );

    \I__9709\ : InMux
    port map (
            O => \N__43577\,
            I => \N__43532\
        );

    \I__9708\ : InMux
    port map (
            O => \N__43576\,
            I => \N__43529\
        );

    \I__9707\ : InMux
    port map (
            O => \N__43575\,
            I => \N__43520\
        );

    \I__9706\ : InMux
    port map (
            O => \N__43574\,
            I => \N__43520\
        );

    \I__9705\ : InMux
    port map (
            O => \N__43573\,
            I => \N__43520\
        );

    \I__9704\ : InMux
    port map (
            O => \N__43572\,
            I => \N__43520\
        );

    \I__9703\ : InMux
    port map (
            O => \N__43571\,
            I => \N__43517\
        );

    \I__9702\ : InMux
    port map (
            O => \N__43568\,
            I => \N__43512\
        );

    \I__9701\ : InMux
    port map (
            O => \N__43567\,
            I => \N__43501\
        );

    \I__9700\ : InMux
    port map (
            O => \N__43566\,
            I => \N__43501\
        );

    \I__9699\ : InMux
    port map (
            O => \N__43563\,
            I => \N__43501\
        );

    \I__9698\ : InMux
    port map (
            O => \N__43562\,
            I => \N__43501\
        );

    \I__9697\ : InMux
    port map (
            O => \N__43561\,
            I => \N__43501\
        );

    \I__9696\ : InMux
    port map (
            O => \N__43560\,
            I => \N__43496\
        );

    \I__9695\ : InMux
    port map (
            O => \N__43559\,
            I => \N__43496\
        );

    \I__9694\ : InMux
    port map (
            O => \N__43558\,
            I => \N__43491\
        );

    \I__9693\ : InMux
    port map (
            O => \N__43557\,
            I => \N__43491\
        );

    \I__9692\ : InMux
    port map (
            O => \N__43556\,
            I => \N__43488\
        );

    \I__9691\ : InMux
    port map (
            O => \N__43555\,
            I => \N__43477\
        );

    \I__9690\ : InMux
    port map (
            O => \N__43554\,
            I => \N__43477\
        );

    \I__9689\ : InMux
    port map (
            O => \N__43553\,
            I => \N__43477\
        );

    \I__9688\ : InMux
    port map (
            O => \N__43552\,
            I => \N__43477\
        );

    \I__9687\ : InMux
    port map (
            O => \N__43551\,
            I => \N__43477\
        );

    \I__9686\ : Span4Mux_v
    port map (
            O => \N__43546\,
            I => \N__43466\
        );

    \I__9685\ : LocalMux
    port map (
            O => \N__43543\,
            I => \N__43466\
        );

    \I__9684\ : LocalMux
    port map (
            O => \N__43532\,
            I => \N__43466\
        );

    \I__9683\ : LocalMux
    port map (
            O => \N__43529\,
            I => \N__43466\
        );

    \I__9682\ : LocalMux
    port map (
            O => \N__43520\,
            I => \N__43466\
        );

    \I__9681\ : LocalMux
    port map (
            O => \N__43517\,
            I => \N__43463\
        );

    \I__9680\ : InMux
    port map (
            O => \N__43516\,
            I => \N__43458\
        );

    \I__9679\ : InMux
    port map (
            O => \N__43515\,
            I => \N__43458\
        );

    \I__9678\ : LocalMux
    port map (
            O => \N__43512\,
            I => \N__43451\
        );

    \I__9677\ : LocalMux
    port map (
            O => \N__43501\,
            I => \N__43451\
        );

    \I__9676\ : LocalMux
    port map (
            O => \N__43496\,
            I => \N__43451\
        );

    \I__9675\ : LocalMux
    port map (
            O => \N__43491\,
            I => \N__43442\
        );

    \I__9674\ : LocalMux
    port map (
            O => \N__43488\,
            I => \N__43442\
        );

    \I__9673\ : LocalMux
    port map (
            O => \N__43477\,
            I => \N__43442\
        );

    \I__9672\ : Span4Mux_h
    port map (
            O => \N__43466\,
            I => \N__43442\
        );

    \I__9671\ : Span4Mux_h
    port map (
            O => \N__43463\,
            I => \N__43439\
        );

    \I__9670\ : LocalMux
    port map (
            O => \N__43458\,
            I => \N__43436\
        );

    \I__9669\ : Span4Mux_h
    port map (
            O => \N__43451\,
            I => \N__43433\
        );

    \I__9668\ : Span4Mux_v
    port map (
            O => \N__43442\,
            I => \N__43430\
        );

    \I__9667\ : Span4Mux_h
    port map (
            O => \N__43439\,
            I => \N__43427\
        );

    \I__9666\ : Span12Mux_h
    port map (
            O => \N__43436\,
            I => \N__43424\
        );

    \I__9665\ : Span4Mux_v
    port map (
            O => \N__43433\,
            I => \N__43419\
        );

    \I__9664\ : Span4Mux_v
    port map (
            O => \N__43430\,
            I => \N__43419\
        );

    \I__9663\ : Odrv4
    port map (
            O => \N__43427\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__9662\ : Odrv12
    port map (
            O => \N__43424\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__9661\ : Odrv4
    port map (
            O => \N__43419\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__9660\ : CascadeMux
    port map (
            O => \N__43412\,
            I => \N__43409\
        );

    \I__9659\ : InMux
    port map (
            O => \N__43409\,
            I => \N__43406\
        );

    \I__9658\ : LocalMux
    port map (
            O => \N__43406\,
            I => \N__43403\
        );

    \I__9657\ : Span4Mux_v
    port map (
            O => \N__43403\,
            I => \N__43400\
        );

    \I__9656\ : Odrv4
    port map (
            O => \N__43400\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt20\
        );

    \I__9655\ : InMux
    port map (
            O => \N__43397\,
            I => \N__43394\
        );

    \I__9654\ : LocalMux
    port map (
            O => \N__43394\,
            I => \N__43391\
        );

    \I__9653\ : Odrv12
    port map (
            O => \N__43391\,
            I => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\
        );

    \I__9652\ : CascadeMux
    port map (
            O => \N__43388\,
            I => \N__43385\
        );

    \I__9651\ : InMux
    port map (
            O => \N__43385\,
            I => \N__43382\
        );

    \I__9650\ : LocalMux
    port map (
            O => \N__43382\,
            I => \N__43379\
        );

    \I__9649\ : Span4Mux_v
    port map (
            O => \N__43379\,
            I => \N__43376\
        );

    \I__9648\ : Odrv4
    port map (
            O => \N__43376\,
            I => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\
        );

    \I__9647\ : InMux
    port map (
            O => \N__43373\,
            I => \N__43370\
        );

    \I__9646\ : LocalMux
    port map (
            O => \N__43370\,
            I => \N__43367\
        );

    \I__9645\ : Span4Mux_v
    port map (
            O => \N__43367\,
            I => \N__43364\
        );

    \I__9644\ : Odrv4
    port map (
            O => \N__43364\,
            I => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\
        );

    \I__9643\ : CascadeMux
    port map (
            O => \N__43361\,
            I => \N__43358\
        );

    \I__9642\ : InMux
    port map (
            O => \N__43358\,
            I => \N__43355\
        );

    \I__9641\ : LocalMux
    port map (
            O => \N__43355\,
            I => \N__43352\
        );

    \I__9640\ : Span4Mux_v
    port map (
            O => \N__43352\,
            I => \N__43349\
        );

    \I__9639\ : Odrv4
    port map (
            O => \N__43349\,
            I => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\
        );

    \I__9638\ : InMux
    port map (
            O => \N__43346\,
            I => \N__43343\
        );

    \I__9637\ : LocalMux
    port map (
            O => \N__43343\,
            I => \N__43340\
        );

    \I__9636\ : Odrv12
    port map (
            O => \N__43340\,
            I => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\
        );

    \I__9635\ : CascadeMux
    port map (
            O => \N__43337\,
            I => \N__43334\
        );

    \I__9634\ : InMux
    port map (
            O => \N__43334\,
            I => \N__43331\
        );

    \I__9633\ : LocalMux
    port map (
            O => \N__43331\,
            I => \N__43328\
        );

    \I__9632\ : Odrv4
    port map (
            O => \N__43328\,
            I => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\
        );

    \I__9631\ : InMux
    port map (
            O => \N__43325\,
            I => \N__43322\
        );

    \I__9630\ : LocalMux
    port map (
            O => \N__43322\,
            I => \N__43319\
        );

    \I__9629\ : Odrv12
    port map (
            O => \N__43319\,
            I => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\
        );

    \I__9628\ : CascadeMux
    port map (
            O => \N__43316\,
            I => \N__43313\
        );

    \I__9627\ : InMux
    port map (
            O => \N__43313\,
            I => \N__43310\
        );

    \I__9626\ : LocalMux
    port map (
            O => \N__43310\,
            I => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\
        );

    \I__9625\ : CascadeMux
    port map (
            O => \N__43307\,
            I => \N__43304\
        );

    \I__9624\ : InMux
    port map (
            O => \N__43304\,
            I => \N__43301\
        );

    \I__9623\ : LocalMux
    port map (
            O => \N__43301\,
            I => \N__43298\
        );

    \I__9622\ : Span4Mux_v
    port map (
            O => \N__43298\,
            I => \N__43295\
        );

    \I__9621\ : Odrv4
    port map (
            O => \N__43295\,
            I => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\
        );

    \I__9620\ : InMux
    port map (
            O => \N__43292\,
            I => \N__43289\
        );

    \I__9619\ : LocalMux
    port map (
            O => \N__43289\,
            I => \N__43286\
        );

    \I__9618\ : Odrv12
    port map (
            O => \N__43286\,
            I => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\
        );

    \I__9617\ : CascadeMux
    port map (
            O => \N__43283\,
            I => \N__43280\
        );

    \I__9616\ : InMux
    port map (
            O => \N__43280\,
            I => \N__43277\
        );

    \I__9615\ : LocalMux
    port map (
            O => \N__43277\,
            I => \N__43274\
        );

    \I__9614\ : Span4Mux_v
    port map (
            O => \N__43274\,
            I => \N__43271\
        );

    \I__9613\ : Odrv4
    port map (
            O => \N__43271\,
            I => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\
        );

    \I__9612\ : CascadeMux
    port map (
            O => \N__43268\,
            I => \N__43265\
        );

    \I__9611\ : InMux
    port map (
            O => \N__43265\,
            I => \N__43262\
        );

    \I__9610\ : LocalMux
    port map (
            O => \N__43262\,
            I => \N__43259\
        );

    \I__9609\ : Span4Mux_v
    port map (
            O => \N__43259\,
            I => \N__43256\
        );

    \I__9608\ : Odrv4
    port map (
            O => \N__43256\,
            I => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\
        );

    \I__9607\ : InMux
    port map (
            O => \N__43253\,
            I => \N__43250\
        );

    \I__9606\ : LocalMux
    port map (
            O => \N__43250\,
            I => \N__43247\
        );

    \I__9605\ : Odrv12
    port map (
            O => \N__43247\,
            I => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\
        );

    \I__9604\ : CascadeMux
    port map (
            O => \N__43244\,
            I => \N__43241\
        );

    \I__9603\ : InMux
    port map (
            O => \N__43241\,
            I => \N__43238\
        );

    \I__9602\ : LocalMux
    port map (
            O => \N__43238\,
            I => \N__43235\
        );

    \I__9601\ : Odrv12
    port map (
            O => \N__43235\,
            I => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\
        );

    \I__9600\ : InMux
    port map (
            O => \N__43232\,
            I => \N__43229\
        );

    \I__9599\ : LocalMux
    port map (
            O => \N__43229\,
            I => \N__43226\
        );

    \I__9598\ : Odrv12
    port map (
            O => \N__43226\,
            I => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\
        );

    \I__9597\ : CascadeMux
    port map (
            O => \N__43223\,
            I => \N__43220\
        );

    \I__9596\ : InMux
    port map (
            O => \N__43220\,
            I => \N__43217\
        );

    \I__9595\ : LocalMux
    port map (
            O => \N__43217\,
            I => \N__43214\
        );

    \I__9594\ : Odrv12
    port map (
            O => \N__43214\,
            I => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\
        );

    \I__9593\ : CascadeMux
    port map (
            O => \N__43211\,
            I => \N__43208\
        );

    \I__9592\ : InMux
    port map (
            O => \N__43208\,
            I => \N__43205\
        );

    \I__9591\ : LocalMux
    port map (
            O => \N__43205\,
            I => \N__43202\
        );

    \I__9590\ : Span4Mux_v
    port map (
            O => \N__43202\,
            I => \N__43199\
        );

    \I__9589\ : Odrv4
    port map (
            O => \N__43199\,
            I => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\
        );

    \I__9588\ : InMux
    port map (
            O => \N__43196\,
            I => \N__43193\
        );

    \I__9587\ : LocalMux
    port map (
            O => \N__43193\,
            I => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\
        );

    \I__9586\ : CascadeMux
    port map (
            O => \N__43190\,
            I => \N__43187\
        );

    \I__9585\ : InMux
    port map (
            O => \N__43187\,
            I => \N__43184\
        );

    \I__9584\ : LocalMux
    port map (
            O => \N__43184\,
            I => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\
        );

    \I__9583\ : InMux
    port map (
            O => \N__43181\,
            I => \N__43178\
        );

    \I__9582\ : LocalMux
    port map (
            O => \N__43178\,
            I => \N__43175\
        );

    \I__9581\ : Span4Mux_v
    port map (
            O => \N__43175\,
            I => \N__43172\
        );

    \I__9580\ : Odrv4
    port map (
            O => \N__43172\,
            I => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\
        );

    \I__9579\ : CascadeMux
    port map (
            O => \N__43169\,
            I => \N__43166\
        );

    \I__9578\ : InMux
    port map (
            O => \N__43166\,
            I => \N__43163\
        );

    \I__9577\ : LocalMux
    port map (
            O => \N__43163\,
            I => \N__43160\
        );

    \I__9576\ : Odrv12
    port map (
            O => \N__43160\,
            I => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\
        );

    \I__9575\ : InMux
    port map (
            O => \N__43157\,
            I => \N__43154\
        );

    \I__9574\ : LocalMux
    port map (
            O => \N__43154\,
            I => \N__43151\
        );

    \I__9573\ : Odrv12
    port map (
            O => \N__43151\,
            I => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\
        );

    \I__9572\ : CascadeMux
    port map (
            O => \N__43148\,
            I => \N__43145\
        );

    \I__9571\ : InMux
    port map (
            O => \N__43145\,
            I => \N__43142\
        );

    \I__9570\ : LocalMux
    port map (
            O => \N__43142\,
            I => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\
        );

    \I__9569\ : CascadeMux
    port map (
            O => \N__43139\,
            I => \N__43133\
        );

    \I__9568\ : InMux
    port map (
            O => \N__43138\,
            I => \N__43130\
        );

    \I__9567\ : InMux
    port map (
            O => \N__43137\,
            I => \N__43125\
        );

    \I__9566\ : InMux
    port map (
            O => \N__43136\,
            I => \N__43125\
        );

    \I__9565\ : InMux
    port map (
            O => \N__43133\,
            I => \N__43122\
        );

    \I__9564\ : LocalMux
    port map (
            O => \N__43130\,
            I => \N__43119\
        );

    \I__9563\ : LocalMux
    port map (
            O => \N__43125\,
            I => \N__43116\
        );

    \I__9562\ : LocalMux
    port map (
            O => \N__43122\,
            I => \N__43113\
        );

    \I__9561\ : Span4Mux_v
    port map (
            O => \N__43119\,
            I => \N__43108\
        );

    \I__9560\ : Span4Mux_v
    port map (
            O => \N__43116\,
            I => \N__43108\
        );

    \I__9559\ : Span4Mux_h
    port map (
            O => \N__43113\,
            I => \N__43105\
        );

    \I__9558\ : Span4Mux_h
    port map (
            O => \N__43108\,
            I => \N__43102\
        );

    \I__9557\ : Odrv4
    port map (
            O => \N__43105\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__9556\ : Odrv4
    port map (
            O => \N__43102\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__9555\ : InMux
    port map (
            O => \N__43097\,
            I => \N__43094\
        );

    \I__9554\ : LocalMux
    port map (
            O => \N__43094\,
            I => \N__43091\
        );

    \I__9553\ : Span4Mux_h
    port map (
            O => \N__43091\,
            I => \N__43086\
        );

    \I__9552\ : InMux
    port map (
            O => \N__43090\,
            I => \N__43083\
        );

    \I__9551\ : InMux
    port map (
            O => \N__43089\,
            I => \N__43080\
        );

    \I__9550\ : Odrv4
    port map (
            O => \N__43086\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__9549\ : LocalMux
    port map (
            O => \N__43083\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__9548\ : LocalMux
    port map (
            O => \N__43080\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__9547\ : InMux
    port map (
            O => \N__43073\,
            I => \N__43070\
        );

    \I__9546\ : LocalMux
    port map (
            O => \N__43070\,
            I => \N__43065\
        );

    \I__9545\ : InMux
    port map (
            O => \N__43069\,
            I => \N__43062\
        );

    \I__9544\ : InMux
    port map (
            O => \N__43068\,
            I => \N__43059\
        );

    \I__9543\ : Span4Mux_h
    port map (
            O => \N__43065\,
            I => \N__43056\
        );

    \I__9542\ : LocalMux
    port map (
            O => \N__43062\,
            I => \N__43050\
        );

    \I__9541\ : LocalMux
    port map (
            O => \N__43059\,
            I => \N__43050\
        );

    \I__9540\ : Span4Mux_h
    port map (
            O => \N__43056\,
            I => \N__43047\
        );

    \I__9539\ : InMux
    port map (
            O => \N__43055\,
            I => \N__43044\
        );

    \I__9538\ : Span4Mux_v
    port map (
            O => \N__43050\,
            I => \N__43041\
        );

    \I__9537\ : Odrv4
    port map (
            O => \N__43047\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__9536\ : LocalMux
    port map (
            O => \N__43044\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__9535\ : Odrv4
    port map (
            O => \N__43041\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__9534\ : CascadeMux
    port map (
            O => \N__43034\,
            I => \N__43030\
        );

    \I__9533\ : InMux
    port map (
            O => \N__43033\,
            I => \N__43026\
        );

    \I__9532\ : InMux
    port map (
            O => \N__43030\,
            I => \N__43023\
        );

    \I__9531\ : CascadeMux
    port map (
            O => \N__43029\,
            I => \N__43020\
        );

    \I__9530\ : LocalMux
    port map (
            O => \N__43026\,
            I => \N__43017\
        );

    \I__9529\ : LocalMux
    port map (
            O => \N__43023\,
            I => \N__43014\
        );

    \I__9528\ : InMux
    port map (
            O => \N__43020\,
            I => \N__43011\
        );

    \I__9527\ : Span4Mux_v
    port map (
            O => \N__43017\,
            I => \N__43008\
        );

    \I__9526\ : Odrv4
    port map (
            O => \N__43014\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__9525\ : LocalMux
    port map (
            O => \N__43011\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__9524\ : Odrv4
    port map (
            O => \N__43008\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__9523\ : CascadeMux
    port map (
            O => \N__43001\,
            I => \N__42997\
        );

    \I__9522\ : InMux
    port map (
            O => \N__43000\,
            I => \N__42993\
        );

    \I__9521\ : InMux
    port map (
            O => \N__42997\,
            I => \N__42990\
        );

    \I__9520\ : CascadeMux
    port map (
            O => \N__42996\,
            I => \N__42987\
        );

    \I__9519\ : LocalMux
    port map (
            O => \N__42993\,
            I => \N__42984\
        );

    \I__9518\ : LocalMux
    port map (
            O => \N__42990\,
            I => \N__42981\
        );

    \I__9517\ : InMux
    port map (
            O => \N__42987\,
            I => \N__42978\
        );

    \I__9516\ : Span4Mux_h
    port map (
            O => \N__42984\,
            I => \N__42975\
        );

    \I__9515\ : Odrv4
    port map (
            O => \N__42981\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__9514\ : LocalMux
    port map (
            O => \N__42978\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__9513\ : Odrv4
    port map (
            O => \N__42975\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__9512\ : CascadeMux
    port map (
            O => \N__42968\,
            I => \N__42965\
        );

    \I__9511\ : InMux
    port map (
            O => \N__42965\,
            I => \N__42962\
        );

    \I__9510\ : LocalMux
    port map (
            O => \N__42962\,
            I => \N__42959\
        );

    \I__9509\ : Span4Mux_v
    port map (
            O => \N__42959\,
            I => \N__42956\
        );

    \I__9508\ : Odrv4
    port map (
            O => \N__42956\,
            I => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\
        );

    \I__9507\ : CascadeMux
    port map (
            O => \N__42953\,
            I => \N__42949\
        );

    \I__9506\ : InMux
    port map (
            O => \N__42952\,
            I => \N__42945\
        );

    \I__9505\ : InMux
    port map (
            O => \N__42949\,
            I => \N__42940\
        );

    \I__9504\ : InMux
    port map (
            O => \N__42948\,
            I => \N__42940\
        );

    \I__9503\ : LocalMux
    port map (
            O => \N__42945\,
            I => \N__42935\
        );

    \I__9502\ : LocalMux
    port map (
            O => \N__42940\,
            I => \N__42935\
        );

    \I__9501\ : Span4Mux_v
    port map (
            O => \N__42935\,
            I => \N__42931\
        );

    \I__9500\ : InMux
    port map (
            O => \N__42934\,
            I => \N__42928\
        );

    \I__9499\ : Odrv4
    port map (
            O => \N__42931\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__9498\ : LocalMux
    port map (
            O => \N__42928\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__9497\ : CascadeMux
    port map (
            O => \N__42923\,
            I => \N__42920\
        );

    \I__9496\ : InMux
    port map (
            O => \N__42920\,
            I => \N__42917\
        );

    \I__9495\ : LocalMux
    port map (
            O => \N__42917\,
            I => \N__42914\
        );

    \I__9494\ : Odrv4
    port map (
            O => \N__42914\,
            I => \current_shift_inst.un4_control_input_1_axb_9\
        );

    \I__9493\ : CascadeMux
    port map (
            O => \N__42911\,
            I => \N__42903\
        );

    \I__9492\ : CascadeMux
    port map (
            O => \N__42910\,
            I => \N__42899\
        );

    \I__9491\ : CascadeMux
    port map (
            O => \N__42909\,
            I => \N__42884\
        );

    \I__9490\ : InMux
    port map (
            O => \N__42908\,
            I => \N__42871\
        );

    \I__9489\ : InMux
    port map (
            O => \N__42907\,
            I => \N__42871\
        );

    \I__9488\ : InMux
    port map (
            O => \N__42906\,
            I => \N__42866\
        );

    \I__9487\ : InMux
    port map (
            O => \N__42903\,
            I => \N__42866\
        );

    \I__9486\ : CascadeMux
    port map (
            O => \N__42902\,
            I => \N__42851\
        );

    \I__9485\ : InMux
    port map (
            O => \N__42899\,
            I => \N__42848\
        );

    \I__9484\ : CascadeMux
    port map (
            O => \N__42898\,
            I => \N__42843\
        );

    \I__9483\ : CascadeMux
    port map (
            O => \N__42897\,
            I => \N__42834\
        );

    \I__9482\ : CascadeMux
    port map (
            O => \N__42896\,
            I => \N__42828\
        );

    \I__9481\ : CascadeMux
    port map (
            O => \N__42895\,
            I => \N__42820\
        );

    \I__9480\ : CascadeMux
    port map (
            O => \N__42894\,
            I => \N__42816\
        );

    \I__9479\ : CascadeMux
    port map (
            O => \N__42893\,
            I => \N__42812\
        );

    \I__9478\ : CascadeMux
    port map (
            O => \N__42892\,
            I => \N__42809\
        );

    \I__9477\ : CascadeMux
    port map (
            O => \N__42891\,
            I => \N__42805\
        );

    \I__9476\ : CascadeMux
    port map (
            O => \N__42890\,
            I => \N__42801\
        );

    \I__9475\ : CascadeMux
    port map (
            O => \N__42889\,
            I => \N__42797\
        );

    \I__9474\ : InMux
    port map (
            O => \N__42888\,
            I => \N__42789\
        );

    \I__9473\ : InMux
    port map (
            O => \N__42887\,
            I => \N__42773\
        );

    \I__9472\ : InMux
    port map (
            O => \N__42884\,
            I => \N__42773\
        );

    \I__9471\ : CascadeMux
    port map (
            O => \N__42883\,
            I => \N__42768\
        );

    \I__9470\ : CascadeMux
    port map (
            O => \N__42882\,
            I => \N__42765\
        );

    \I__9469\ : InMux
    port map (
            O => \N__42881\,
            I => \N__42762\
        );

    \I__9468\ : InMux
    port map (
            O => \N__42880\,
            I => \N__42757\
        );

    \I__9467\ : InMux
    port map (
            O => \N__42879\,
            I => \N__42757\
        );

    \I__9466\ : CascadeMux
    port map (
            O => \N__42878\,
            I => \N__42754\
        );

    \I__9465\ : CascadeMux
    port map (
            O => \N__42877\,
            I => \N__42750\
        );

    \I__9464\ : CascadeMux
    port map (
            O => \N__42876\,
            I => \N__42746\
        );

    \I__9463\ : LocalMux
    port map (
            O => \N__42871\,
            I => \N__42740\
        );

    \I__9462\ : LocalMux
    port map (
            O => \N__42866\,
            I => \N__42740\
        );

    \I__9461\ : CascadeMux
    port map (
            O => \N__42865\,
            I => \N__42737\
        );

    \I__9460\ : CascadeMux
    port map (
            O => \N__42864\,
            I => \N__42734\
        );

    \I__9459\ : CascadeMux
    port map (
            O => \N__42863\,
            I => \N__42731\
        );

    \I__9458\ : CascadeMux
    port map (
            O => \N__42862\,
            I => \N__42727\
        );

    \I__9457\ : CascadeMux
    port map (
            O => \N__42861\,
            I => \N__42724\
        );

    \I__9456\ : InMux
    port map (
            O => \N__42860\,
            I => \N__42713\
        );

    \I__9455\ : InMux
    port map (
            O => \N__42859\,
            I => \N__42710\
        );

    \I__9454\ : InMux
    port map (
            O => \N__42858\,
            I => \N__42697\
        );

    \I__9453\ : InMux
    port map (
            O => \N__42857\,
            I => \N__42697\
        );

    \I__9452\ : InMux
    port map (
            O => \N__42856\,
            I => \N__42697\
        );

    \I__9451\ : InMux
    port map (
            O => \N__42855\,
            I => \N__42697\
        );

    \I__9450\ : InMux
    port map (
            O => \N__42854\,
            I => \N__42697\
        );

    \I__9449\ : InMux
    port map (
            O => \N__42851\,
            I => \N__42697\
        );

    \I__9448\ : LocalMux
    port map (
            O => \N__42848\,
            I => \N__42694\
        );

    \I__9447\ : InMux
    port map (
            O => \N__42847\,
            I => \N__42689\
        );

    \I__9446\ : InMux
    port map (
            O => \N__42846\,
            I => \N__42689\
        );

    \I__9445\ : InMux
    port map (
            O => \N__42843\,
            I => \N__42674\
        );

    \I__9444\ : InMux
    port map (
            O => \N__42842\,
            I => \N__42674\
        );

    \I__9443\ : InMux
    port map (
            O => \N__42841\,
            I => \N__42674\
        );

    \I__9442\ : InMux
    port map (
            O => \N__42840\,
            I => \N__42674\
        );

    \I__9441\ : InMux
    port map (
            O => \N__42839\,
            I => \N__42674\
        );

    \I__9440\ : InMux
    port map (
            O => \N__42838\,
            I => \N__42674\
        );

    \I__9439\ : InMux
    port map (
            O => \N__42837\,
            I => \N__42674\
        );

    \I__9438\ : InMux
    port map (
            O => \N__42834\,
            I => \N__42659\
        );

    \I__9437\ : InMux
    port map (
            O => \N__42833\,
            I => \N__42659\
        );

    \I__9436\ : InMux
    port map (
            O => \N__42832\,
            I => \N__42659\
        );

    \I__9435\ : InMux
    port map (
            O => \N__42831\,
            I => \N__42659\
        );

    \I__9434\ : InMux
    port map (
            O => \N__42828\,
            I => \N__42659\
        );

    \I__9433\ : InMux
    port map (
            O => \N__42827\,
            I => \N__42659\
        );

    \I__9432\ : InMux
    port map (
            O => \N__42826\,
            I => \N__42659\
        );

    \I__9431\ : InMux
    port map (
            O => \N__42825\,
            I => \N__42656\
        );

    \I__9430\ : InMux
    port map (
            O => \N__42824\,
            I => \N__42641\
        );

    \I__9429\ : InMux
    port map (
            O => \N__42823\,
            I => \N__42641\
        );

    \I__9428\ : InMux
    port map (
            O => \N__42820\,
            I => \N__42641\
        );

    \I__9427\ : InMux
    port map (
            O => \N__42819\,
            I => \N__42641\
        );

    \I__9426\ : InMux
    port map (
            O => \N__42816\,
            I => \N__42641\
        );

    \I__9425\ : InMux
    port map (
            O => \N__42815\,
            I => \N__42641\
        );

    \I__9424\ : InMux
    port map (
            O => \N__42812\,
            I => \N__42641\
        );

    \I__9423\ : InMux
    port map (
            O => \N__42809\,
            I => \N__42624\
        );

    \I__9422\ : InMux
    port map (
            O => \N__42808\,
            I => \N__42624\
        );

    \I__9421\ : InMux
    port map (
            O => \N__42805\,
            I => \N__42624\
        );

    \I__9420\ : InMux
    port map (
            O => \N__42804\,
            I => \N__42624\
        );

    \I__9419\ : InMux
    port map (
            O => \N__42801\,
            I => \N__42624\
        );

    \I__9418\ : InMux
    port map (
            O => \N__42800\,
            I => \N__42624\
        );

    \I__9417\ : InMux
    port map (
            O => \N__42797\,
            I => \N__42624\
        );

    \I__9416\ : InMux
    port map (
            O => \N__42796\,
            I => \N__42624\
        );

    \I__9415\ : CascadeMux
    port map (
            O => \N__42795\,
            I => \N__42621\
        );

    \I__9414\ : CascadeMux
    port map (
            O => \N__42794\,
            I => \N__42617\
        );

    \I__9413\ : CascadeMux
    port map (
            O => \N__42793\,
            I => \N__42613\
        );

    \I__9412\ : CascadeMux
    port map (
            O => \N__42792\,
            I => \N__42609\
        );

    \I__9411\ : LocalMux
    port map (
            O => \N__42789\,
            I => \N__42602\
        );

    \I__9410\ : InMux
    port map (
            O => \N__42788\,
            I => \N__42595\
        );

    \I__9409\ : InMux
    port map (
            O => \N__42787\,
            I => \N__42595\
        );

    \I__9408\ : InMux
    port map (
            O => \N__42786\,
            I => \N__42595\
        );

    \I__9407\ : CascadeMux
    port map (
            O => \N__42785\,
            I => \N__42592\
        );

    \I__9406\ : CascadeMux
    port map (
            O => \N__42784\,
            I => \N__42588\
        );

    \I__9405\ : CascadeMux
    port map (
            O => \N__42783\,
            I => \N__42584\
        );

    \I__9404\ : CascadeMux
    port map (
            O => \N__42782\,
            I => \N__42580\
        );

    \I__9403\ : CascadeMux
    port map (
            O => \N__42781\,
            I => \N__42576\
        );

    \I__9402\ : CascadeMux
    port map (
            O => \N__42780\,
            I => \N__42572\
        );

    \I__9401\ : CascadeMux
    port map (
            O => \N__42779\,
            I => \N__42568\
        );

    \I__9400\ : CascadeMux
    port map (
            O => \N__42778\,
            I => \N__42564\
        );

    \I__9399\ : LocalMux
    port map (
            O => \N__42773\,
            I => \N__42560\
        );

    \I__9398\ : InMux
    port map (
            O => \N__42772\,
            I => \N__42553\
        );

    \I__9397\ : InMux
    port map (
            O => \N__42771\,
            I => \N__42553\
        );

    \I__9396\ : InMux
    port map (
            O => \N__42768\,
            I => \N__42553\
        );

    \I__9395\ : InMux
    port map (
            O => \N__42765\,
            I => \N__42550\
        );

    \I__9394\ : LocalMux
    port map (
            O => \N__42762\,
            I => \N__42545\
        );

    \I__9393\ : LocalMux
    port map (
            O => \N__42757\,
            I => \N__42545\
        );

    \I__9392\ : InMux
    port map (
            O => \N__42754\,
            I => \N__42532\
        );

    \I__9391\ : InMux
    port map (
            O => \N__42753\,
            I => \N__42532\
        );

    \I__9390\ : InMux
    port map (
            O => \N__42750\,
            I => \N__42532\
        );

    \I__9389\ : InMux
    port map (
            O => \N__42749\,
            I => \N__42532\
        );

    \I__9388\ : InMux
    port map (
            O => \N__42746\,
            I => \N__42532\
        );

    \I__9387\ : InMux
    port map (
            O => \N__42745\,
            I => \N__42532\
        );

    \I__9386\ : Span4Mux_v
    port map (
            O => \N__42740\,
            I => \N__42529\
        );

    \I__9385\ : InMux
    port map (
            O => \N__42737\,
            I => \N__42524\
        );

    \I__9384\ : InMux
    port map (
            O => \N__42734\,
            I => \N__42524\
        );

    \I__9383\ : InMux
    port map (
            O => \N__42731\,
            I => \N__42513\
        );

    \I__9382\ : InMux
    port map (
            O => \N__42730\,
            I => \N__42513\
        );

    \I__9381\ : InMux
    port map (
            O => \N__42727\,
            I => \N__42513\
        );

    \I__9380\ : InMux
    port map (
            O => \N__42724\,
            I => \N__42513\
        );

    \I__9379\ : InMux
    port map (
            O => \N__42723\,
            I => \N__42513\
        );

    \I__9378\ : CascadeMux
    port map (
            O => \N__42722\,
            I => \N__42508\
        );

    \I__9377\ : CascadeMux
    port map (
            O => \N__42721\,
            I => \N__42505\
        );

    \I__9376\ : CascadeMux
    port map (
            O => \N__42720\,
            I => \N__42499\
        );

    \I__9375\ : CascadeMux
    port map (
            O => \N__42719\,
            I => \N__42495\
        );

    \I__9374\ : CascadeMux
    port map (
            O => \N__42718\,
            I => \N__42491\
        );

    \I__9373\ : CascadeMux
    port map (
            O => \N__42717\,
            I => \N__42487\
        );

    \I__9372\ : CascadeMux
    port map (
            O => \N__42716\,
            I => \N__42483\
        );

    \I__9371\ : LocalMux
    port map (
            O => \N__42713\,
            I => \N__42475\
        );

    \I__9370\ : LocalMux
    port map (
            O => \N__42710\,
            I => \N__42475\
        );

    \I__9369\ : LocalMux
    port map (
            O => \N__42697\,
            I => \N__42475\
        );

    \I__9368\ : Span4Mux_v
    port map (
            O => \N__42694\,
            I => \N__42460\
        );

    \I__9367\ : LocalMux
    port map (
            O => \N__42689\,
            I => \N__42460\
        );

    \I__9366\ : LocalMux
    port map (
            O => \N__42674\,
            I => \N__42460\
        );

    \I__9365\ : LocalMux
    port map (
            O => \N__42659\,
            I => \N__42460\
        );

    \I__9364\ : LocalMux
    port map (
            O => \N__42656\,
            I => \N__42460\
        );

    \I__9363\ : LocalMux
    port map (
            O => \N__42641\,
            I => \N__42460\
        );

    \I__9362\ : LocalMux
    port map (
            O => \N__42624\,
            I => \N__42460\
        );

    \I__9361\ : InMux
    port map (
            O => \N__42621\,
            I => \N__42443\
        );

    \I__9360\ : InMux
    port map (
            O => \N__42620\,
            I => \N__42443\
        );

    \I__9359\ : InMux
    port map (
            O => \N__42617\,
            I => \N__42443\
        );

    \I__9358\ : InMux
    port map (
            O => \N__42616\,
            I => \N__42443\
        );

    \I__9357\ : InMux
    port map (
            O => \N__42613\,
            I => \N__42443\
        );

    \I__9356\ : InMux
    port map (
            O => \N__42612\,
            I => \N__42443\
        );

    \I__9355\ : InMux
    port map (
            O => \N__42609\,
            I => \N__42443\
        );

    \I__9354\ : InMux
    port map (
            O => \N__42608\,
            I => \N__42443\
        );

    \I__9353\ : CascadeMux
    port map (
            O => \N__42607\,
            I => \N__42440\
        );

    \I__9352\ : CascadeMux
    port map (
            O => \N__42606\,
            I => \N__42436\
        );

    \I__9351\ : CascadeMux
    port map (
            O => \N__42605\,
            I => \N__42432\
        );

    \I__9350\ : Span4Mux_v
    port map (
            O => \N__42602\,
            I => \N__42426\
        );

    \I__9349\ : LocalMux
    port map (
            O => \N__42595\,
            I => \N__42426\
        );

    \I__9348\ : InMux
    port map (
            O => \N__42592\,
            I => \N__42423\
        );

    \I__9347\ : InMux
    port map (
            O => \N__42591\,
            I => \N__42408\
        );

    \I__9346\ : InMux
    port map (
            O => \N__42588\,
            I => \N__42408\
        );

    \I__9345\ : InMux
    port map (
            O => \N__42587\,
            I => \N__42408\
        );

    \I__9344\ : InMux
    port map (
            O => \N__42584\,
            I => \N__42408\
        );

    \I__9343\ : InMux
    port map (
            O => \N__42583\,
            I => \N__42408\
        );

    \I__9342\ : InMux
    port map (
            O => \N__42580\,
            I => \N__42408\
        );

    \I__9341\ : InMux
    port map (
            O => \N__42579\,
            I => \N__42408\
        );

    \I__9340\ : InMux
    port map (
            O => \N__42576\,
            I => \N__42391\
        );

    \I__9339\ : InMux
    port map (
            O => \N__42575\,
            I => \N__42391\
        );

    \I__9338\ : InMux
    port map (
            O => \N__42572\,
            I => \N__42391\
        );

    \I__9337\ : InMux
    port map (
            O => \N__42571\,
            I => \N__42391\
        );

    \I__9336\ : InMux
    port map (
            O => \N__42568\,
            I => \N__42391\
        );

    \I__9335\ : InMux
    port map (
            O => \N__42567\,
            I => \N__42391\
        );

    \I__9334\ : InMux
    port map (
            O => \N__42564\,
            I => \N__42391\
        );

    \I__9333\ : InMux
    port map (
            O => \N__42563\,
            I => \N__42391\
        );

    \I__9332\ : Span4Mux_v
    port map (
            O => \N__42560\,
            I => \N__42380\
        );

    \I__9331\ : LocalMux
    port map (
            O => \N__42553\,
            I => \N__42380\
        );

    \I__9330\ : LocalMux
    port map (
            O => \N__42550\,
            I => \N__42380\
        );

    \I__9329\ : Span4Mux_h
    port map (
            O => \N__42545\,
            I => \N__42380\
        );

    \I__9328\ : LocalMux
    port map (
            O => \N__42532\,
            I => \N__42380\
        );

    \I__9327\ : Span4Mux_h
    port map (
            O => \N__42529\,
            I => \N__42377\
        );

    \I__9326\ : LocalMux
    port map (
            O => \N__42524\,
            I => \N__42372\
        );

    \I__9325\ : LocalMux
    port map (
            O => \N__42513\,
            I => \N__42372\
        );

    \I__9324\ : InMux
    port map (
            O => \N__42512\,
            I => \N__42359\
        );

    \I__9323\ : InMux
    port map (
            O => \N__42511\,
            I => \N__42359\
        );

    \I__9322\ : InMux
    port map (
            O => \N__42508\,
            I => \N__42359\
        );

    \I__9321\ : InMux
    port map (
            O => \N__42505\,
            I => \N__42359\
        );

    \I__9320\ : InMux
    port map (
            O => \N__42504\,
            I => \N__42359\
        );

    \I__9319\ : InMux
    port map (
            O => \N__42503\,
            I => \N__42359\
        );

    \I__9318\ : InMux
    port map (
            O => \N__42502\,
            I => \N__42352\
        );

    \I__9317\ : InMux
    port map (
            O => \N__42499\,
            I => \N__42352\
        );

    \I__9316\ : InMux
    port map (
            O => \N__42498\,
            I => \N__42352\
        );

    \I__9315\ : InMux
    port map (
            O => \N__42495\,
            I => \N__42335\
        );

    \I__9314\ : InMux
    port map (
            O => \N__42494\,
            I => \N__42335\
        );

    \I__9313\ : InMux
    port map (
            O => \N__42491\,
            I => \N__42335\
        );

    \I__9312\ : InMux
    port map (
            O => \N__42490\,
            I => \N__42335\
        );

    \I__9311\ : InMux
    port map (
            O => \N__42487\,
            I => \N__42335\
        );

    \I__9310\ : InMux
    port map (
            O => \N__42486\,
            I => \N__42335\
        );

    \I__9309\ : InMux
    port map (
            O => \N__42483\,
            I => \N__42335\
        );

    \I__9308\ : InMux
    port map (
            O => \N__42482\,
            I => \N__42335\
        );

    \I__9307\ : Span4Mux_h
    port map (
            O => \N__42475\,
            I => \N__42328\
        );

    \I__9306\ : Span4Mux_v
    port map (
            O => \N__42460\,
            I => \N__42328\
        );

    \I__9305\ : LocalMux
    port map (
            O => \N__42443\,
            I => \N__42328\
        );

    \I__9304\ : InMux
    port map (
            O => \N__42440\,
            I => \N__42315\
        );

    \I__9303\ : InMux
    port map (
            O => \N__42439\,
            I => \N__42315\
        );

    \I__9302\ : InMux
    port map (
            O => \N__42436\,
            I => \N__42315\
        );

    \I__9301\ : InMux
    port map (
            O => \N__42435\,
            I => \N__42315\
        );

    \I__9300\ : InMux
    port map (
            O => \N__42432\,
            I => \N__42315\
        );

    \I__9299\ : InMux
    port map (
            O => \N__42431\,
            I => \N__42315\
        );

    \I__9298\ : Span4Mux_h
    port map (
            O => \N__42426\,
            I => \N__42304\
        );

    \I__9297\ : LocalMux
    port map (
            O => \N__42423\,
            I => \N__42304\
        );

    \I__9296\ : LocalMux
    port map (
            O => \N__42408\,
            I => \N__42304\
        );

    \I__9295\ : LocalMux
    port map (
            O => \N__42391\,
            I => \N__42304\
        );

    \I__9294\ : Span4Mux_h
    port map (
            O => \N__42380\,
            I => \N__42304\
        );

    \I__9293\ : Odrv4
    port map (
            O => \N__42377\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__9292\ : Odrv4
    port map (
            O => \N__42372\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__9291\ : LocalMux
    port map (
            O => \N__42359\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__9290\ : LocalMux
    port map (
            O => \N__42352\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__9289\ : LocalMux
    port map (
            O => \N__42335\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__9288\ : Odrv4
    port map (
            O => \N__42328\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__9287\ : LocalMux
    port map (
            O => \N__42315\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__9286\ : Odrv4
    port map (
            O => \N__42304\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__9285\ : CascadeMux
    port map (
            O => \N__42287\,
            I => \N__42282\
        );

    \I__9284\ : InMux
    port map (
            O => \N__42286\,
            I => \N__42279\
        );

    \I__9283\ : InMux
    port map (
            O => \N__42285\,
            I => \N__42276\
        );

    \I__9282\ : InMux
    port map (
            O => \N__42282\,
            I => \N__42273\
        );

    \I__9281\ : LocalMux
    port map (
            O => \N__42279\,
            I => \N__42270\
        );

    \I__9280\ : LocalMux
    port map (
            O => \N__42276\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__9279\ : LocalMux
    port map (
            O => \N__42273\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__9278\ : Odrv12
    port map (
            O => \N__42270\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__9277\ : CascadeMux
    port map (
            O => \N__42263\,
            I => \N__42260\
        );

    \I__9276\ : InMux
    port map (
            O => \N__42260\,
            I => \N__42257\
        );

    \I__9275\ : LocalMux
    port map (
            O => \N__42257\,
            I => \N__42252\
        );

    \I__9274\ : InMux
    port map (
            O => \N__42256\,
            I => \N__42249\
        );

    \I__9273\ : InMux
    port map (
            O => \N__42255\,
            I => \N__42246\
        );

    \I__9272\ : Span4Mux_h
    port map (
            O => \N__42252\,
            I => \N__42242\
        );

    \I__9271\ : LocalMux
    port map (
            O => \N__42249\,
            I => \N__42239\
        );

    \I__9270\ : LocalMux
    port map (
            O => \N__42246\,
            I => \N__42236\
        );

    \I__9269\ : InMux
    port map (
            O => \N__42245\,
            I => \N__42233\
        );

    \I__9268\ : Odrv4
    port map (
            O => \N__42242\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__9267\ : Odrv4
    port map (
            O => \N__42239\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__9266\ : Odrv4
    port map (
            O => \N__42236\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__9265\ : LocalMux
    port map (
            O => \N__42233\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__9264\ : InMux
    port map (
            O => \N__42224\,
            I => \N__42221\
        );

    \I__9263\ : LocalMux
    port map (
            O => \N__42221\,
            I => \N__42218\
        );

    \I__9262\ : Span4Mux_h
    port map (
            O => \N__42218\,
            I => \N__42215\
        );

    \I__9261\ : Span4Mux_h
    port map (
            O => \N__42215\,
            I => \N__42212\
        );

    \I__9260\ : Odrv4
    port map (
            O => \N__42212\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\
        );

    \I__9259\ : CascadeMux
    port map (
            O => \N__42209\,
            I => \N__42205\
        );

    \I__9258\ : InMux
    port map (
            O => \N__42208\,
            I => \N__42202\
        );

    \I__9257\ : InMux
    port map (
            O => \N__42205\,
            I => \N__42199\
        );

    \I__9256\ : LocalMux
    port map (
            O => \N__42202\,
            I => \N__42195\
        );

    \I__9255\ : LocalMux
    port map (
            O => \N__42199\,
            I => \N__42192\
        );

    \I__9254\ : InMux
    port map (
            O => \N__42198\,
            I => \N__42189\
        );

    \I__9253\ : Span4Mux_v
    port map (
            O => \N__42195\,
            I => \N__42185\
        );

    \I__9252\ : Span4Mux_h
    port map (
            O => \N__42192\,
            I => \N__42180\
        );

    \I__9251\ : LocalMux
    port map (
            O => \N__42189\,
            I => \N__42180\
        );

    \I__9250\ : InMux
    port map (
            O => \N__42188\,
            I => \N__42177\
        );

    \I__9249\ : Odrv4
    port map (
            O => \N__42185\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__9248\ : Odrv4
    port map (
            O => \N__42180\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__9247\ : LocalMux
    port map (
            O => \N__42177\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__9246\ : InMux
    port map (
            O => \N__42170\,
            I => \N__42166\
        );

    \I__9245\ : CascadeMux
    port map (
            O => \N__42169\,
            I => \N__42163\
        );

    \I__9244\ : LocalMux
    port map (
            O => \N__42166\,
            I => \N__42159\
        );

    \I__9243\ : InMux
    port map (
            O => \N__42163\,
            I => \N__42156\
        );

    \I__9242\ : InMux
    port map (
            O => \N__42162\,
            I => \N__42153\
        );

    \I__9241\ : Odrv4
    port map (
            O => \N__42159\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__9240\ : LocalMux
    port map (
            O => \N__42156\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__9239\ : LocalMux
    port map (
            O => \N__42153\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__9238\ : CascadeMux
    port map (
            O => \N__42146\,
            I => \N__42142\
        );

    \I__9237\ : InMux
    port map (
            O => \N__42145\,
            I => \N__42139\
        );

    \I__9236\ : InMux
    port map (
            O => \N__42142\,
            I => \N__42136\
        );

    \I__9235\ : LocalMux
    port map (
            O => \N__42139\,
            I => \N__42133\
        );

    \I__9234\ : LocalMux
    port map (
            O => \N__42136\,
            I => \N__42126\
        );

    \I__9233\ : Span4Mux_v
    port map (
            O => \N__42133\,
            I => \N__42126\
        );

    \I__9232\ : InMux
    port map (
            O => \N__42132\,
            I => \N__42123\
        );

    \I__9231\ : InMux
    port map (
            O => \N__42131\,
            I => \N__42120\
        );

    \I__9230\ : Odrv4
    port map (
            O => \N__42126\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__9229\ : LocalMux
    port map (
            O => \N__42123\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__9228\ : LocalMux
    port map (
            O => \N__42120\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__9227\ : InMux
    port map (
            O => \N__42113\,
            I => \N__42110\
        );

    \I__9226\ : LocalMux
    port map (
            O => \N__42110\,
            I => \N__42105\
        );

    \I__9225\ : InMux
    port map (
            O => \N__42109\,
            I => \N__42102\
        );

    \I__9224\ : InMux
    port map (
            O => \N__42108\,
            I => \N__42099\
        );

    \I__9223\ : Span4Mux_v
    port map (
            O => \N__42105\,
            I => \N__42094\
        );

    \I__9222\ : LocalMux
    port map (
            O => \N__42102\,
            I => \N__42094\
        );

    \I__9221\ : LocalMux
    port map (
            O => \N__42099\,
            I => \N__42091\
        );

    \I__9220\ : Span4Mux_v
    port map (
            O => \N__42094\,
            I => \N__42086\
        );

    \I__9219\ : Span4Mux_v
    port map (
            O => \N__42091\,
            I => \N__42086\
        );

    \I__9218\ : Odrv4
    port map (
            O => \N__42086\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__9217\ : CascadeMux
    port map (
            O => \N__42083\,
            I => \N__42080\
        );

    \I__9216\ : InMux
    port map (
            O => \N__42080\,
            I => \N__42077\
        );

    \I__9215\ : LocalMux
    port map (
            O => \N__42077\,
            I => \N__42072\
        );

    \I__9214\ : InMux
    port map (
            O => \N__42076\,
            I => \N__42069\
        );

    \I__9213\ : InMux
    port map (
            O => \N__42075\,
            I => \N__42066\
        );

    \I__9212\ : Span4Mux_h
    port map (
            O => \N__42072\,
            I => \N__42060\
        );

    \I__9211\ : LocalMux
    port map (
            O => \N__42069\,
            I => \N__42060\
        );

    \I__9210\ : LocalMux
    port map (
            O => \N__42066\,
            I => \N__42057\
        );

    \I__9209\ : InMux
    port map (
            O => \N__42065\,
            I => \N__42054\
        );

    \I__9208\ : Odrv4
    port map (
            O => \N__42060\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__9207\ : Odrv4
    port map (
            O => \N__42057\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__9206\ : LocalMux
    port map (
            O => \N__42054\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__9205\ : InMux
    port map (
            O => \N__42047\,
            I => \N__42044\
        );

    \I__9204\ : LocalMux
    port map (
            O => \N__42044\,
            I => \N__42041\
        );

    \I__9203\ : Span4Mux_h
    port map (
            O => \N__42041\,
            I => \N__42038\
        );

    \I__9202\ : Odrv4
    port map (
            O => \N__42038\,
            I => \current_shift_inst.un4_control_input_1_axb_13\
        );

    \I__9201\ : CascadeMux
    port map (
            O => \N__42035\,
            I => \N__42031\
        );

    \I__9200\ : CascadeMux
    port map (
            O => \N__42034\,
            I => \N__42028\
        );

    \I__9199\ : InMux
    port map (
            O => \N__42031\,
            I => \N__42023\
        );

    \I__9198\ : InMux
    port map (
            O => \N__42028\,
            I => \N__42023\
        );

    \I__9197\ : LocalMux
    port map (
            O => \N__42023\,
            I => \N__42018\
        );

    \I__9196\ : InMux
    port map (
            O => \N__42022\,
            I => \N__42015\
        );

    \I__9195\ : InMux
    port map (
            O => \N__42021\,
            I => \N__42012\
        );

    \I__9194\ : Span4Mux_h
    port map (
            O => \N__42018\,
            I => \N__42007\
        );

    \I__9193\ : LocalMux
    port map (
            O => \N__42015\,
            I => \N__42007\
        );

    \I__9192\ : LocalMux
    port map (
            O => \N__42012\,
            I => \N__42004\
        );

    \I__9191\ : Odrv4
    port map (
            O => \N__42007\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__9190\ : Odrv12
    port map (
            O => \N__42004\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__9189\ : InMux
    port map (
            O => \N__41999\,
            I => \N__41993\
        );

    \I__9188\ : InMux
    port map (
            O => \N__41998\,
            I => \N__41993\
        );

    \I__9187\ : LocalMux
    port map (
            O => \N__41993\,
            I => \N__41989\
        );

    \I__9186\ : InMux
    port map (
            O => \N__41992\,
            I => \N__41986\
        );

    \I__9185\ : Span4Mux_h
    port map (
            O => \N__41989\,
            I => \N__41981\
        );

    \I__9184\ : LocalMux
    port map (
            O => \N__41986\,
            I => \N__41981\
        );

    \I__9183\ : Span4Mux_v
    port map (
            O => \N__41981\,
            I => \N__41978\
        );

    \I__9182\ : Odrv4
    port map (
            O => \N__41978\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__9181\ : CascadeMux
    port map (
            O => \N__41975\,
            I => \N__41971\
        );

    \I__9180\ : CascadeMux
    port map (
            O => \N__41974\,
            I => \N__41968\
        );

    \I__9179\ : InMux
    port map (
            O => \N__41971\,
            I => \N__41965\
        );

    \I__9178\ : InMux
    port map (
            O => \N__41968\,
            I => \N__41962\
        );

    \I__9177\ : LocalMux
    port map (
            O => \N__41965\,
            I => \N__41959\
        );

    \I__9176\ : LocalMux
    port map (
            O => \N__41962\,
            I => \N__41955\
        );

    \I__9175\ : Sp12to4
    port map (
            O => \N__41959\,
            I => \N__41952\
        );

    \I__9174\ : InMux
    port map (
            O => \N__41958\,
            I => \N__41949\
        );

    \I__9173\ : Span4Mux_v
    port map (
            O => \N__41955\,
            I => \N__41945\
        );

    \I__9172\ : Span12Mux_v
    port map (
            O => \N__41952\,
            I => \N__41942\
        );

    \I__9171\ : LocalMux
    port map (
            O => \N__41949\,
            I => \N__41939\
        );

    \I__9170\ : InMux
    port map (
            O => \N__41948\,
            I => \N__41936\
        );

    \I__9169\ : Odrv4
    port map (
            O => \N__41945\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__9168\ : Odrv12
    port map (
            O => \N__41942\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__9167\ : Odrv4
    port map (
            O => \N__41939\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__9166\ : LocalMux
    port map (
            O => \N__41936\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__9165\ : InMux
    port map (
            O => \N__41927\,
            I => \N__41923\
        );

    \I__9164\ : InMux
    port map (
            O => \N__41926\,
            I => \N__41920\
        );

    \I__9163\ : LocalMux
    port map (
            O => \N__41923\,
            I => \N__41917\
        );

    \I__9162\ : LocalMux
    port map (
            O => \N__41920\,
            I => \N__41911\
        );

    \I__9161\ : Span4Mux_v
    port map (
            O => \N__41917\,
            I => \N__41911\
        );

    \I__9160\ : InMux
    port map (
            O => \N__41916\,
            I => \N__41908\
        );

    \I__9159\ : Odrv4
    port map (
            O => \N__41911\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__9158\ : LocalMux
    port map (
            O => \N__41908\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__9157\ : InMux
    port map (
            O => \N__41903\,
            I => \N__41900\
        );

    \I__9156\ : LocalMux
    port map (
            O => \N__41900\,
            I => \current_shift_inst.un4_control_input_1_axb_23\
        );

    \I__9155\ : InMux
    port map (
            O => \N__41897\,
            I => \N__41892\
        );

    \I__9154\ : InMux
    port map (
            O => \N__41896\,
            I => \N__41889\
        );

    \I__9153\ : InMux
    port map (
            O => \N__41895\,
            I => \N__41886\
        );

    \I__9152\ : LocalMux
    port map (
            O => \N__41892\,
            I => \N__41880\
        );

    \I__9151\ : LocalMux
    port map (
            O => \N__41889\,
            I => \N__41880\
        );

    \I__9150\ : LocalMux
    port map (
            O => \N__41886\,
            I => \N__41877\
        );

    \I__9149\ : InMux
    port map (
            O => \N__41885\,
            I => \N__41874\
        );

    \I__9148\ : Span4Mux_h
    port map (
            O => \N__41880\,
            I => \N__41867\
        );

    \I__9147\ : Span4Mux_v
    port map (
            O => \N__41877\,
            I => \N__41867\
        );

    \I__9146\ : LocalMux
    port map (
            O => \N__41874\,
            I => \N__41867\
        );

    \I__9145\ : Odrv4
    port map (
            O => \N__41867\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__9144\ : InMux
    port map (
            O => \N__41864\,
            I => \N__41861\
        );

    \I__9143\ : LocalMux
    port map (
            O => \N__41861\,
            I => \current_shift_inst.un4_control_input_1_axb_17\
        );

    \I__9142\ : CascadeMux
    port map (
            O => \N__41858\,
            I => \N__41853\
        );

    \I__9141\ : InMux
    port map (
            O => \N__41857\,
            I => \N__41850\
        );

    \I__9140\ : InMux
    port map (
            O => \N__41856\,
            I => \N__41847\
        );

    \I__9139\ : InMux
    port map (
            O => \N__41853\,
            I => \N__41844\
        );

    \I__9138\ : LocalMux
    port map (
            O => \N__41850\,
            I => \N__41840\
        );

    \I__9137\ : LocalMux
    port map (
            O => \N__41847\,
            I => \N__41837\
        );

    \I__9136\ : LocalMux
    port map (
            O => \N__41844\,
            I => \N__41834\
        );

    \I__9135\ : InMux
    port map (
            O => \N__41843\,
            I => \N__41831\
        );

    \I__9134\ : Span4Mux_h
    port map (
            O => \N__41840\,
            I => \N__41828\
        );

    \I__9133\ : Span4Mux_h
    port map (
            O => \N__41837\,
            I => \N__41825\
        );

    \I__9132\ : Span4Mux_v
    port map (
            O => \N__41834\,
            I => \N__41820\
        );

    \I__9131\ : LocalMux
    port map (
            O => \N__41831\,
            I => \N__41820\
        );

    \I__9130\ : Odrv4
    port map (
            O => \N__41828\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__9129\ : Odrv4
    port map (
            O => \N__41825\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__9128\ : Odrv4
    port map (
            O => \N__41820\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__9127\ : InMux
    port map (
            O => \N__41813\,
            I => \N__41810\
        );

    \I__9126\ : LocalMux
    port map (
            O => \N__41810\,
            I => \N__41805\
        );

    \I__9125\ : InMux
    port map (
            O => \N__41809\,
            I => \N__41802\
        );

    \I__9124\ : InMux
    port map (
            O => \N__41808\,
            I => \N__41799\
        );

    \I__9123\ : Odrv4
    port map (
            O => \N__41805\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__9122\ : LocalMux
    port map (
            O => \N__41802\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__9121\ : LocalMux
    port map (
            O => \N__41799\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__9120\ : CascadeMux
    port map (
            O => \N__41792\,
            I => \N__41788\
        );

    \I__9119\ : InMux
    port map (
            O => \N__41791\,
            I => \N__41785\
        );

    \I__9118\ : InMux
    port map (
            O => \N__41788\,
            I => \N__41782\
        );

    \I__9117\ : LocalMux
    port map (
            O => \N__41785\,
            I => \N__41778\
        );

    \I__9116\ : LocalMux
    port map (
            O => \N__41782\,
            I => \N__41775\
        );

    \I__9115\ : InMux
    port map (
            O => \N__41781\,
            I => \N__41772\
        );

    \I__9114\ : Span4Mux_v
    port map (
            O => \N__41778\,
            I => \N__41766\
        );

    \I__9113\ : Span4Mux_h
    port map (
            O => \N__41775\,
            I => \N__41766\
        );

    \I__9112\ : LocalMux
    port map (
            O => \N__41772\,
            I => \N__41763\
        );

    \I__9111\ : InMux
    port map (
            O => \N__41771\,
            I => \N__41760\
        );

    \I__9110\ : Odrv4
    port map (
            O => \N__41766\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__9109\ : Odrv4
    port map (
            O => \N__41763\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__9108\ : LocalMux
    port map (
            O => \N__41760\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__9107\ : InMux
    port map (
            O => \N__41753\,
            I => \N__41749\
        );

    \I__9106\ : CascadeMux
    port map (
            O => \N__41752\,
            I => \N__41746\
        );

    \I__9105\ : LocalMux
    port map (
            O => \N__41749\,
            I => \N__41743\
        );

    \I__9104\ : InMux
    port map (
            O => \N__41746\,
            I => \N__41739\
        );

    \I__9103\ : Span4Mux_h
    port map (
            O => \N__41743\,
            I => \N__41736\
        );

    \I__9102\ : InMux
    port map (
            O => \N__41742\,
            I => \N__41733\
        );

    \I__9101\ : LocalMux
    port map (
            O => \N__41739\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__9100\ : Odrv4
    port map (
            O => \N__41736\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__9099\ : LocalMux
    port map (
            O => \N__41733\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__9098\ : CascadeMux
    port map (
            O => \N__41726\,
            I => \N__41722\
        );

    \I__9097\ : InMux
    port map (
            O => \N__41725\,
            I => \N__41716\
        );

    \I__9096\ : InMux
    port map (
            O => \N__41722\,
            I => \N__41716\
        );

    \I__9095\ : InMux
    port map (
            O => \N__41721\,
            I => \N__41713\
        );

    \I__9094\ : LocalMux
    port map (
            O => \N__41716\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__9093\ : LocalMux
    port map (
            O => \N__41713\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__9092\ : InMux
    port map (
            O => \N__41708\,
            I => \N__41700\
        );

    \I__9091\ : InMux
    port map (
            O => \N__41707\,
            I => \N__41700\
        );

    \I__9090\ : InMux
    port map (
            O => \N__41706\,
            I => \N__41695\
        );

    \I__9089\ : InMux
    port map (
            O => \N__41705\,
            I => \N__41695\
        );

    \I__9088\ : LocalMux
    port map (
            O => \N__41700\,
            I => \N__41692\
        );

    \I__9087\ : LocalMux
    port map (
            O => \N__41695\,
            I => \N__41689\
        );

    \I__9086\ : Odrv4
    port map (
            O => \N__41692\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__9085\ : Odrv4
    port map (
            O => \N__41689\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__9084\ : CascadeMux
    port map (
            O => \N__41684\,
            I => \N__41681\
        );

    \I__9083\ : InMux
    port map (
            O => \N__41681\,
            I => \N__41678\
        );

    \I__9082\ : LocalMux
    port map (
            O => \N__41678\,
            I => \current_shift_inst.un4_control_input_1_axb_20\
        );

    \I__9081\ : InMux
    port map (
            O => \N__41675\,
            I => \N__41672\
        );

    \I__9080\ : LocalMux
    port map (
            O => \N__41672\,
            I => \N__41667\
        );

    \I__9079\ : InMux
    port map (
            O => \N__41671\,
            I => \N__41664\
        );

    \I__9078\ : InMux
    port map (
            O => \N__41670\,
            I => \N__41661\
        );

    \I__9077\ : Span4Mux_v
    port map (
            O => \N__41667\,
            I => \N__41657\
        );

    \I__9076\ : LocalMux
    port map (
            O => \N__41664\,
            I => \N__41654\
        );

    \I__9075\ : LocalMux
    port map (
            O => \N__41661\,
            I => \N__41651\
        );

    \I__9074\ : InMux
    port map (
            O => \N__41660\,
            I => \N__41648\
        );

    \I__9073\ : Odrv4
    port map (
            O => \N__41657\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__9072\ : Odrv4
    port map (
            O => \N__41654\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__9071\ : Odrv4
    port map (
            O => \N__41651\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__9070\ : LocalMux
    port map (
            O => \N__41648\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__9069\ : CascadeMux
    port map (
            O => \N__41639\,
            I => \N__41635\
        );

    \I__9068\ : InMux
    port map (
            O => \N__41638\,
            I => \N__41632\
        );

    \I__9067\ : InMux
    port map (
            O => \N__41635\,
            I => \N__41628\
        );

    \I__9066\ : LocalMux
    port map (
            O => \N__41632\,
            I => \N__41625\
        );

    \I__9065\ : InMux
    port map (
            O => \N__41631\,
            I => \N__41622\
        );

    \I__9064\ : LocalMux
    port map (
            O => \N__41628\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__9063\ : Odrv4
    port map (
            O => \N__41625\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__9062\ : LocalMux
    port map (
            O => \N__41622\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__9061\ : CascadeMux
    port map (
            O => \N__41615\,
            I => \N__41611\
        );

    \I__9060\ : CascadeMux
    port map (
            O => \N__41614\,
            I => \N__41608\
        );

    \I__9059\ : InMux
    port map (
            O => \N__41611\,
            I => \N__41604\
        );

    \I__9058\ : InMux
    port map (
            O => \N__41608\,
            I => \N__41599\
        );

    \I__9057\ : InMux
    port map (
            O => \N__41607\,
            I => \N__41599\
        );

    \I__9056\ : LocalMux
    port map (
            O => \N__41604\,
            I => \N__41595\
        );

    \I__9055\ : LocalMux
    port map (
            O => \N__41599\,
            I => \N__41592\
        );

    \I__9054\ : InMux
    port map (
            O => \N__41598\,
            I => \N__41589\
        );

    \I__9053\ : Span4Mux_v
    port map (
            O => \N__41595\,
            I => \N__41586\
        );

    \I__9052\ : Span4Mux_h
    port map (
            O => \N__41592\,
            I => \N__41583\
        );

    \I__9051\ : LocalMux
    port map (
            O => \N__41589\,
            I => \N__41580\
        );

    \I__9050\ : Odrv4
    port map (
            O => \N__41586\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__9049\ : Odrv4
    port map (
            O => \N__41583\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__9048\ : Odrv12
    port map (
            O => \N__41580\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__9047\ : InMux
    port map (
            O => \N__41573\,
            I => \N__41570\
        );

    \I__9046\ : LocalMux
    port map (
            O => \N__41570\,
            I => \N__41567\
        );

    \I__9045\ : Span4Mux_h
    port map (
            O => \N__41567\,
            I => \N__41562\
        );

    \I__9044\ : InMux
    port map (
            O => \N__41566\,
            I => \N__41557\
        );

    \I__9043\ : InMux
    port map (
            O => \N__41565\,
            I => \N__41557\
        );

    \I__9042\ : Odrv4
    port map (
            O => \N__41562\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__9041\ : LocalMux
    port map (
            O => \N__41557\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__9040\ : CascadeMux
    port map (
            O => \N__41552\,
            I => \N__41549\
        );

    \I__9039\ : InMux
    port map (
            O => \N__41549\,
            I => \N__41546\
        );

    \I__9038\ : LocalMux
    port map (
            O => \N__41546\,
            I => \N__41543\
        );

    \I__9037\ : Span4Mux_h
    port map (
            O => \N__41543\,
            I => \N__41540\
        );

    \I__9036\ : Odrv4
    port map (
            O => \N__41540\,
            I => \current_shift_inst.un38_control_input_cry_0_s0_sf\
        );

    \I__9035\ : InMux
    port map (
            O => \N__41537\,
            I => \N__41532\
        );

    \I__9034\ : InMux
    port map (
            O => \N__41536\,
            I => \N__41529\
        );

    \I__9033\ : InMux
    port map (
            O => \N__41535\,
            I => \N__41526\
        );

    \I__9032\ : LocalMux
    port map (
            O => \N__41532\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__9031\ : LocalMux
    port map (
            O => \N__41529\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__9030\ : LocalMux
    port map (
            O => \N__41526\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__9029\ : InMux
    port map (
            O => \N__41519\,
            I => \N__41514\
        );

    \I__9028\ : InMux
    port map (
            O => \N__41518\,
            I => \N__41508\
        );

    \I__9027\ : InMux
    port map (
            O => \N__41517\,
            I => \N__41508\
        );

    \I__9026\ : LocalMux
    port map (
            O => \N__41514\,
            I => \N__41505\
        );

    \I__9025\ : InMux
    port map (
            O => \N__41513\,
            I => \N__41502\
        );

    \I__9024\ : LocalMux
    port map (
            O => \N__41508\,
            I => \N__41499\
        );

    \I__9023\ : Span4Mux_h
    port map (
            O => \N__41505\,
            I => \N__41496\
        );

    \I__9022\ : LocalMux
    port map (
            O => \N__41502\,
            I => \N__41493\
        );

    \I__9021\ : Span4Mux_v
    port map (
            O => \N__41499\,
            I => \N__41490\
        );

    \I__9020\ : Odrv4
    port map (
            O => \N__41496\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__9019\ : Odrv4
    port map (
            O => \N__41493\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__9018\ : Odrv4
    port map (
            O => \N__41490\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__9017\ : InMux
    port map (
            O => \N__41483\,
            I => \N__41480\
        );

    \I__9016\ : LocalMux
    port map (
            O => \N__41480\,
            I => \N__41476\
        );

    \I__9015\ : InMux
    port map (
            O => \N__41479\,
            I => \N__41473\
        );

    \I__9014\ : Span4Mux_h
    port map (
            O => \N__41476\,
            I => \N__41469\
        );

    \I__9013\ : LocalMux
    port map (
            O => \N__41473\,
            I => \N__41466\
        );

    \I__9012\ : InMux
    port map (
            O => \N__41472\,
            I => \N__41463\
        );

    \I__9011\ : Odrv4
    port map (
            O => \N__41469\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__9010\ : Odrv4
    port map (
            O => \N__41466\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__9009\ : LocalMux
    port map (
            O => \N__41463\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__9008\ : CascadeMux
    port map (
            O => \N__41456\,
            I => \N__41453\
        );

    \I__9007\ : InMux
    port map (
            O => \N__41453\,
            I => \N__41450\
        );

    \I__9006\ : LocalMux
    port map (
            O => \N__41450\,
            I => \N__41447\
        );

    \I__9005\ : Span4Mux_h
    port map (
            O => \N__41447\,
            I => \N__41444\
        );

    \I__9004\ : Odrv4
    port map (
            O => \N__41444\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI34N61_5\
        );

    \I__9003\ : CascadeMux
    port map (
            O => \N__41441\,
            I => \N__41437\
        );

    \I__9002\ : CascadeMux
    port map (
            O => \N__41440\,
            I => \N__41434\
        );

    \I__9001\ : InMux
    port map (
            O => \N__41437\,
            I => \N__41431\
        );

    \I__9000\ : InMux
    port map (
            O => \N__41434\,
            I => \N__41428\
        );

    \I__8999\ : LocalMux
    port map (
            O => \N__41431\,
            I => \N__41422\
        );

    \I__8998\ : LocalMux
    port map (
            O => \N__41428\,
            I => \N__41422\
        );

    \I__8997\ : InMux
    port map (
            O => \N__41427\,
            I => \N__41419\
        );

    \I__8996\ : Span4Mux_h
    port map (
            O => \N__41422\,
            I => \N__41413\
        );

    \I__8995\ : LocalMux
    port map (
            O => \N__41419\,
            I => \N__41413\
        );

    \I__8994\ : InMux
    port map (
            O => \N__41418\,
            I => \N__41410\
        );

    \I__8993\ : Odrv4
    port map (
            O => \N__41413\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__8992\ : LocalMux
    port map (
            O => \N__41410\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__8991\ : InMux
    port map (
            O => \N__41405\,
            I => \N__41402\
        );

    \I__8990\ : LocalMux
    port map (
            O => \N__41402\,
            I => \N__41398\
        );

    \I__8989\ : InMux
    port map (
            O => \N__41401\,
            I => \N__41394\
        );

    \I__8988\ : Span4Mux_h
    port map (
            O => \N__41398\,
            I => \N__41391\
        );

    \I__8987\ : InMux
    port map (
            O => \N__41397\,
            I => \N__41388\
        );

    \I__8986\ : LocalMux
    port map (
            O => \N__41394\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__8985\ : Odrv4
    port map (
            O => \N__41391\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__8984\ : LocalMux
    port map (
            O => \N__41388\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__8983\ : CascadeMux
    port map (
            O => \N__41381\,
            I => \N__41378\
        );

    \I__8982\ : InMux
    port map (
            O => \N__41378\,
            I => \N__41373\
        );

    \I__8981\ : InMux
    port map (
            O => \N__41377\,
            I => \N__41370\
        );

    \I__8980\ : InMux
    port map (
            O => \N__41376\,
            I => \N__41366\
        );

    \I__8979\ : LocalMux
    port map (
            O => \N__41373\,
            I => \N__41361\
        );

    \I__8978\ : LocalMux
    port map (
            O => \N__41370\,
            I => \N__41361\
        );

    \I__8977\ : InMux
    port map (
            O => \N__41369\,
            I => \N__41358\
        );

    \I__8976\ : LocalMux
    port map (
            O => \N__41366\,
            I => \N__41355\
        );

    \I__8975\ : Span4Mux_h
    port map (
            O => \N__41361\,
            I => \N__41350\
        );

    \I__8974\ : LocalMux
    port map (
            O => \N__41358\,
            I => \N__41350\
        );

    \I__8973\ : Odrv4
    port map (
            O => \N__41355\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__8972\ : Odrv4
    port map (
            O => \N__41350\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__8971\ : InMux
    port map (
            O => \N__41345\,
            I => \N__41341\
        );

    \I__8970\ : InMux
    port map (
            O => \N__41344\,
            I => \N__41338\
        );

    \I__8969\ : LocalMux
    port map (
            O => \N__41341\,
            I => \N__41334\
        );

    \I__8968\ : LocalMux
    port map (
            O => \N__41338\,
            I => \N__41331\
        );

    \I__8967\ : InMux
    port map (
            O => \N__41337\,
            I => \N__41328\
        );

    \I__8966\ : Odrv4
    port map (
            O => \N__41334\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__8965\ : Odrv12
    port map (
            O => \N__41331\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__8964\ : LocalMux
    port map (
            O => \N__41328\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__8963\ : CascadeMux
    port map (
            O => \N__41321\,
            I => \N__41318\
        );

    \I__8962\ : InMux
    port map (
            O => \N__41318\,
            I => \N__41315\
        );

    \I__8961\ : LocalMux
    port map (
            O => \N__41315\,
            I => \N__41312\
        );

    \I__8960\ : Span4Mux_h
    port map (
            O => \N__41312\,
            I => \N__41309\
        );

    \I__8959\ : Span4Mux_h
    port map (
            O => \N__41309\,
            I => \N__41306\
        );

    \I__8958\ : Odrv4
    port map (
            O => \N__41306\,
            I => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\
        );

    \I__8957\ : InMux
    port map (
            O => \N__41303\,
            I => \N__41298\
        );

    \I__8956\ : InMux
    port map (
            O => \N__41302\,
            I => \N__41295\
        );

    \I__8955\ : InMux
    port map (
            O => \N__41301\,
            I => \N__41292\
        );

    \I__8954\ : LocalMux
    port map (
            O => \N__41298\,
            I => \N__41289\
        );

    \I__8953\ : LocalMux
    port map (
            O => \N__41295\,
            I => \N__41286\
        );

    \I__8952\ : LocalMux
    port map (
            O => \N__41292\,
            I => \N__41283\
        );

    \I__8951\ : Span4Mux_v
    port map (
            O => \N__41289\,
            I => \N__41280\
        );

    \I__8950\ : Span4Mux_h
    port map (
            O => \N__41286\,
            I => \N__41275\
        );

    \I__8949\ : Span4Mux_v
    port map (
            O => \N__41283\,
            I => \N__41275\
        );

    \I__8948\ : Span4Mux_h
    port map (
            O => \N__41280\,
            I => \N__41269\
        );

    \I__8947\ : Span4Mux_v
    port map (
            O => \N__41275\,
            I => \N__41269\
        );

    \I__8946\ : InMux
    port map (
            O => \N__41274\,
            I => \N__41266\
        );

    \I__8945\ : Sp12to4
    port map (
            O => \N__41269\,
            I => \N__41263\
        );

    \I__8944\ : LocalMux
    port map (
            O => \N__41266\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__8943\ : Odrv12
    port map (
            O => \N__41263\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__8942\ : InMux
    port map (
            O => \N__41258\,
            I => \N__41255\
        );

    \I__8941\ : LocalMux
    port map (
            O => \N__41255\,
            I => \current_shift_inst.un4_control_input_1_axb_26\
        );

    \I__8940\ : InMux
    port map (
            O => \N__41252\,
            I => \N__41247\
        );

    \I__8939\ : CascadeMux
    port map (
            O => \N__41251\,
            I => \N__41244\
        );

    \I__8938\ : InMux
    port map (
            O => \N__41250\,
            I => \N__41241\
        );

    \I__8937\ : LocalMux
    port map (
            O => \N__41247\,
            I => \N__41238\
        );

    \I__8936\ : InMux
    port map (
            O => \N__41244\,
            I => \N__41235\
        );

    \I__8935\ : LocalMux
    port map (
            O => \N__41241\,
            I => \N__41232\
        );

    \I__8934\ : Span4Mux_v
    port map (
            O => \N__41238\,
            I => \N__41228\
        );

    \I__8933\ : LocalMux
    port map (
            O => \N__41235\,
            I => \N__41225\
        );

    \I__8932\ : Span4Mux_h
    port map (
            O => \N__41232\,
            I => \N__41222\
        );

    \I__8931\ : InMux
    port map (
            O => \N__41231\,
            I => \N__41219\
        );

    \I__8930\ : Odrv4
    port map (
            O => \N__41228\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__8929\ : Odrv4
    port map (
            O => \N__41225\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__8928\ : Odrv4
    port map (
            O => \N__41222\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__8927\ : LocalMux
    port map (
            O => \N__41219\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__8926\ : InMux
    port map (
            O => \N__41210\,
            I => \N__41206\
        );

    \I__8925\ : InMux
    port map (
            O => \N__41209\,
            I => \N__41203\
        );

    \I__8924\ : LocalMux
    port map (
            O => \N__41206\,
            I => \N__41200\
        );

    \I__8923\ : LocalMux
    port map (
            O => \N__41203\,
            I => \N__41196\
        );

    \I__8922\ : Span4Mux_h
    port map (
            O => \N__41200\,
            I => \N__41193\
        );

    \I__8921\ : InMux
    port map (
            O => \N__41199\,
            I => \N__41190\
        );

    \I__8920\ : Odrv12
    port map (
            O => \N__41196\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__8919\ : Odrv4
    port map (
            O => \N__41193\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__8918\ : LocalMux
    port map (
            O => \N__41190\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__8917\ : CascadeMux
    port map (
            O => \N__41183\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\
        );

    \I__8916\ : CascadeMux
    port map (
            O => \N__41180\,
            I => \N__41176\
        );

    \I__8915\ : InMux
    port map (
            O => \N__41179\,
            I => \N__41173\
        );

    \I__8914\ : InMux
    port map (
            O => \N__41176\,
            I => \N__41170\
        );

    \I__8913\ : LocalMux
    port map (
            O => \N__41173\,
            I => \N__41167\
        );

    \I__8912\ : LocalMux
    port map (
            O => \N__41170\,
            I => \N__41164\
        );

    \I__8911\ : Span4Mux_h
    port map (
            O => \N__41167\,
            I => \N__41159\
        );

    \I__8910\ : Span4Mux_v
    port map (
            O => \N__41164\,
            I => \N__41159\
        );

    \I__8909\ : Odrv4
    port map (
            O => \N__41159\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__8908\ : CascadeMux
    port map (
            O => \N__41156\,
            I => \N__41153\
        );

    \I__8907\ : InMux
    port map (
            O => \N__41153\,
            I => \N__41150\
        );

    \I__8906\ : LocalMux
    port map (
            O => \N__41150\,
            I => \N__41147\
        );

    \I__8905\ : Span4Mux_h
    port map (
            O => \N__41147\,
            I => \N__41144\
        );

    \I__8904\ : Odrv4
    port map (
            O => \N__41144\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\
        );

    \I__8903\ : InMux
    port map (
            O => \N__41141\,
            I => \N__41138\
        );

    \I__8902\ : LocalMux
    port map (
            O => \N__41138\,
            I => \N__41135\
        );

    \I__8901\ : Span4Mux_h
    port map (
            O => \N__41135\,
            I => \N__41129\
        );

    \I__8900\ : InMux
    port map (
            O => \N__41134\,
            I => \N__41126\
        );

    \I__8899\ : InMux
    port map (
            O => \N__41133\,
            I => \N__41121\
        );

    \I__8898\ : InMux
    port map (
            O => \N__41132\,
            I => \N__41121\
        );

    \I__8897\ : Span4Mux_h
    port map (
            O => \N__41129\,
            I => \N__41116\
        );

    \I__8896\ : LocalMux
    port map (
            O => \N__41126\,
            I => \N__41116\
        );

    \I__8895\ : LocalMux
    port map (
            O => \N__41121\,
            I => \N__41113\
        );

    \I__8894\ : Odrv4
    port map (
            O => \N__41116\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__8893\ : Odrv12
    port map (
            O => \N__41113\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__8892\ : InMux
    port map (
            O => \N__41108\,
            I => \N__41105\
        );

    \I__8891\ : LocalMux
    port map (
            O => \N__41105\,
            I => \N__41100\
        );

    \I__8890\ : InMux
    port map (
            O => \N__41104\,
            I => \N__41097\
        );

    \I__8889\ : InMux
    port map (
            O => \N__41103\,
            I => \N__41094\
        );

    \I__8888\ : Odrv4
    port map (
            O => \N__41100\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__8887\ : LocalMux
    port map (
            O => \N__41097\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__8886\ : LocalMux
    port map (
            O => \N__41094\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__8885\ : CascadeMux
    port map (
            O => \N__41087\,
            I => \N__41084\
        );

    \I__8884\ : InMux
    port map (
            O => \N__41084\,
            I => \N__41081\
        );

    \I__8883\ : LocalMux
    port map (
            O => \N__41081\,
            I => \N__41076\
        );

    \I__8882\ : InMux
    port map (
            O => \N__41080\,
            I => \N__41073\
        );

    \I__8881\ : InMux
    port map (
            O => \N__41079\,
            I => \N__41070\
        );

    \I__8880\ : Span4Mux_h
    port map (
            O => \N__41076\,
            I => \N__41065\
        );

    \I__8879\ : LocalMux
    port map (
            O => \N__41073\,
            I => \N__41065\
        );

    \I__8878\ : LocalMux
    port map (
            O => \N__41070\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__8877\ : Odrv4
    port map (
            O => \N__41065\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__8876\ : InMux
    port map (
            O => \N__41060\,
            I => \N__41056\
        );

    \I__8875\ : CascadeMux
    port map (
            O => \N__41059\,
            I => \N__41052\
        );

    \I__8874\ : LocalMux
    port map (
            O => \N__41056\,
            I => \N__41049\
        );

    \I__8873\ : InMux
    port map (
            O => \N__41055\,
            I => \N__41045\
        );

    \I__8872\ : InMux
    port map (
            O => \N__41052\,
            I => \N__41042\
        );

    \I__8871\ : Span4Mux_h
    port map (
            O => \N__41049\,
            I => \N__41039\
        );

    \I__8870\ : InMux
    port map (
            O => \N__41048\,
            I => \N__41036\
        );

    \I__8869\ : LocalMux
    port map (
            O => \N__41045\,
            I => \N__41033\
        );

    \I__8868\ : LocalMux
    port map (
            O => \N__41042\,
            I => \N__41030\
        );

    \I__8867\ : Span4Mux_v
    port map (
            O => \N__41039\,
            I => \N__41025\
        );

    \I__8866\ : LocalMux
    port map (
            O => \N__41036\,
            I => \N__41025\
        );

    \I__8865\ : Odrv12
    port map (
            O => \N__41033\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__8864\ : Odrv4
    port map (
            O => \N__41030\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__8863\ : Odrv4
    port map (
            O => \N__41025\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__8862\ : CascadeMux
    port map (
            O => \N__41018\,
            I => \N__41014\
        );

    \I__8861\ : InMux
    port map (
            O => \N__41017\,
            I => \N__41011\
        );

    \I__8860\ : InMux
    port map (
            O => \N__41014\,
            I => \N__41008\
        );

    \I__8859\ : LocalMux
    port map (
            O => \N__41011\,
            I => \N__41005\
        );

    \I__8858\ : LocalMux
    port map (
            O => \N__41008\,
            I => \N__41002\
        );

    \I__8857\ : Span4Mux_h
    port map (
            O => \N__41005\,
            I => \N__40999\
        );

    \I__8856\ : Span4Mux_h
    port map (
            O => \N__41002\,
            I => \N__40993\
        );

    \I__8855\ : Span4Mux_v
    port map (
            O => \N__40999\,
            I => \N__40993\
        );

    \I__8854\ : InMux
    port map (
            O => \N__40998\,
            I => \N__40990\
        );

    \I__8853\ : Odrv4
    port map (
            O => \N__40993\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__8852\ : LocalMux
    port map (
            O => \N__40990\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__8851\ : InMux
    port map (
            O => \N__40985\,
            I => \N__40980\
        );

    \I__8850\ : InMux
    port map (
            O => \N__40984\,
            I => \N__40977\
        );

    \I__8849\ : InMux
    port map (
            O => \N__40983\,
            I => \N__40974\
        );

    \I__8848\ : LocalMux
    port map (
            O => \N__40980\,
            I => \N__40971\
        );

    \I__8847\ : LocalMux
    port map (
            O => \N__40977\,
            I => \N__40968\
        );

    \I__8846\ : LocalMux
    port map (
            O => \N__40974\,
            I => \N__40965\
        );

    \I__8845\ : Span4Mux_v
    port map (
            O => \N__40971\,
            I => \N__40957\
        );

    \I__8844\ : Span4Mux_h
    port map (
            O => \N__40968\,
            I => \N__40957\
        );

    \I__8843\ : Span4Mux_h
    port map (
            O => \N__40965\,
            I => \N__40957\
        );

    \I__8842\ : InMux
    port map (
            O => \N__40964\,
            I => \N__40954\
        );

    \I__8841\ : Odrv4
    port map (
            O => \N__40957\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__8840\ : LocalMux
    port map (
            O => \N__40954\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__8839\ : CascadeMux
    port map (
            O => \N__40949\,
            I => \N__40945\
        );

    \I__8838\ : InMux
    port map (
            O => \N__40948\,
            I => \N__40942\
        );

    \I__8837\ : InMux
    port map (
            O => \N__40945\,
            I => \N__40939\
        );

    \I__8836\ : LocalMux
    port map (
            O => \N__40942\,
            I => \N__40936\
        );

    \I__8835\ : LocalMux
    port map (
            O => \N__40939\,
            I => \N__40933\
        );

    \I__8834\ : Span4Mux_h
    port map (
            O => \N__40936\,
            I => \N__40929\
        );

    \I__8833\ : Span4Mux_h
    port map (
            O => \N__40933\,
            I => \N__40926\
        );

    \I__8832\ : InMux
    port map (
            O => \N__40932\,
            I => \N__40923\
        );

    \I__8831\ : Odrv4
    port map (
            O => \N__40929\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__8830\ : Odrv4
    port map (
            O => \N__40926\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__8829\ : LocalMux
    port map (
            O => \N__40923\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__8828\ : InMux
    port map (
            O => \N__40916\,
            I => \N__40913\
        );

    \I__8827\ : LocalMux
    port map (
            O => \N__40913\,
            I => \current_shift_inst.un4_control_input_1_axb_1\
        );

    \I__8826\ : CascadeMux
    port map (
            O => \N__40910\,
            I => \N__40906\
        );

    \I__8825\ : CascadeMux
    port map (
            O => \N__40909\,
            I => \N__40903\
        );

    \I__8824\ : InMux
    port map (
            O => \N__40906\,
            I => \N__40900\
        );

    \I__8823\ : InMux
    port map (
            O => \N__40903\,
            I => \N__40896\
        );

    \I__8822\ : LocalMux
    port map (
            O => \N__40900\,
            I => \N__40893\
        );

    \I__8821\ : InMux
    port map (
            O => \N__40899\,
            I => \N__40890\
        );

    \I__8820\ : LocalMux
    port map (
            O => \N__40896\,
            I => \N__40887\
        );

    \I__8819\ : Span4Mux_v
    port map (
            O => \N__40893\,
            I => \N__40883\
        );

    \I__8818\ : LocalMux
    port map (
            O => \N__40890\,
            I => \N__40880\
        );

    \I__8817\ : Span4Mux_v
    port map (
            O => \N__40887\,
            I => \N__40877\
        );

    \I__8816\ : InMux
    port map (
            O => \N__40886\,
            I => \N__40874\
        );

    \I__8815\ : Span4Mux_h
    port map (
            O => \N__40883\,
            I => \N__40869\
        );

    \I__8814\ : Span4Mux_v
    port map (
            O => \N__40880\,
            I => \N__40869\
        );

    \I__8813\ : Odrv4
    port map (
            O => \N__40877\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__8812\ : LocalMux
    port map (
            O => \N__40874\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__8811\ : Odrv4
    port map (
            O => \N__40869\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__8810\ : CascadeMux
    port map (
            O => \N__40862\,
            I => \N__40859\
        );

    \I__8809\ : InMux
    port map (
            O => \N__40859\,
            I => \N__40856\
        );

    \I__8808\ : LocalMux
    port map (
            O => \N__40856\,
            I => \N__40853\
        );

    \I__8807\ : Span4Mux_v
    port map (
            O => \N__40853\,
            I => \N__40850\
        );

    \I__8806\ : Odrv4
    port map (
            O => \N__40850\,
            I => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\
        );

    \I__8805\ : InMux
    port map (
            O => \N__40847\,
            I => \N__40844\
        );

    \I__8804\ : LocalMux
    port map (
            O => \N__40844\,
            I => \N__40841\
        );

    \I__8803\ : Span4Mux_h
    port map (
            O => \N__40841\,
            I => \N__40838\
        );

    \I__8802\ : Span4Mux_v
    port map (
            O => \N__40838\,
            I => \N__40832\
        );

    \I__8801\ : InMux
    port map (
            O => \N__40837\,
            I => \N__40829\
        );

    \I__8800\ : InMux
    port map (
            O => \N__40836\,
            I => \N__40824\
        );

    \I__8799\ : InMux
    port map (
            O => \N__40835\,
            I => \N__40824\
        );

    \I__8798\ : Odrv4
    port map (
            O => \N__40832\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__8797\ : LocalMux
    port map (
            O => \N__40829\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__8796\ : LocalMux
    port map (
            O => \N__40824\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__8795\ : InMux
    port map (
            O => \N__40817\,
            I => \N__40814\
        );

    \I__8794\ : LocalMux
    port map (
            O => \N__40814\,
            I => \N__40811\
        );

    \I__8793\ : Span4Mux_v
    port map (
            O => \N__40811\,
            I => \N__40806\
        );

    \I__8792\ : InMux
    port map (
            O => \N__40810\,
            I => \N__40803\
        );

    \I__8791\ : InMux
    port map (
            O => \N__40809\,
            I => \N__40800\
        );

    \I__8790\ : Odrv4
    port map (
            O => \N__40806\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__8789\ : LocalMux
    port map (
            O => \N__40803\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__8788\ : LocalMux
    port map (
            O => \N__40800\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__8787\ : InMux
    port map (
            O => \N__40793\,
            I => \N__40790\
        );

    \I__8786\ : LocalMux
    port map (
            O => \N__40790\,
            I => \N__40787\
        );

    \I__8785\ : Span4Mux_h
    port map (
            O => \N__40787\,
            I => \N__40784\
        );

    \I__8784\ : Span4Mux_h
    port map (
            O => \N__40784\,
            I => \N__40781\
        );

    \I__8783\ : Odrv4
    port map (
            O => \N__40781\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\
        );

    \I__8782\ : InMux
    port map (
            O => \N__40778\,
            I => \N__40775\
        );

    \I__8781\ : LocalMux
    port map (
            O => \N__40775\,
            I => \N__40772\
        );

    \I__8780\ : Span4Mux_h
    port map (
            O => \N__40772\,
            I => \N__40769\
        );

    \I__8779\ : Odrv4
    port map (
            O => \N__40769\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\
        );

    \I__8778\ : InMux
    port map (
            O => \N__40766\,
            I => \N__40763\
        );

    \I__8777\ : LocalMux
    port map (
            O => \N__40763\,
            I => \N__40760\
        );

    \I__8776\ : Span4Mux_h
    port map (
            O => \N__40760\,
            I => \N__40757\
        );

    \I__8775\ : Span4Mux_v
    port map (
            O => \N__40757\,
            I => \N__40754\
        );

    \I__8774\ : Odrv4
    port map (
            O => \N__40754\,
            I => \current_shift_inst.un38_control_input_axb_31_s0\
        );

    \I__8773\ : CascadeMux
    port map (
            O => \N__40751\,
            I => \N__40747\
        );

    \I__8772\ : InMux
    port map (
            O => \N__40750\,
            I => \N__40739\
        );

    \I__8771\ : InMux
    port map (
            O => \N__40747\,
            I => \N__40739\
        );

    \I__8770\ : InMux
    port map (
            O => \N__40746\,
            I => \N__40739\
        );

    \I__8769\ : LocalMux
    port map (
            O => \N__40739\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__8768\ : InMux
    port map (
            O => \N__40736\,
            I => \N__40733\
        );

    \I__8767\ : LocalMux
    port map (
            O => \N__40733\,
            I => \N__40730\
        );

    \I__8766\ : Odrv4
    port map (
            O => \N__40730\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\
        );

    \I__8765\ : CascadeMux
    port map (
            O => \N__40727\,
            I => \N__40724\
        );

    \I__8764\ : InMux
    port map (
            O => \N__40724\,
            I => \N__40721\
        );

    \I__8763\ : LocalMux
    port map (
            O => \N__40721\,
            I => \N__40718\
        );

    \I__8762\ : Odrv12
    port map (
            O => \N__40718\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt30\
        );

    \I__8761\ : InMux
    port map (
            O => \N__40715\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30\
        );

    \I__8760\ : InMux
    port map (
            O => \N__40712\,
            I => \N__40709\
        );

    \I__8759\ : LocalMux
    port map (
            O => \N__40709\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt24\
        );

    \I__8758\ : CascadeMux
    port map (
            O => \N__40706\,
            I => \N__40703\
        );

    \I__8757\ : InMux
    port map (
            O => \N__40703\,
            I => \N__40700\
        );

    \I__8756\ : LocalMux
    port map (
            O => \N__40700\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24\
        );

    \I__8755\ : InMux
    port map (
            O => \N__40697\,
            I => \N__40694\
        );

    \I__8754\ : LocalMux
    port map (
            O => \N__40694\,
            I => \N__40691\
        );

    \I__8753\ : Span4Mux_h
    port map (
            O => \N__40691\,
            I => \N__40687\
        );

    \I__8752\ : InMux
    port map (
            O => \N__40690\,
            I => \N__40684\
        );

    \I__8751\ : Odrv4
    port map (
            O => \N__40687\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__8750\ : LocalMux
    port map (
            O => \N__40684\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__8749\ : CascadeMux
    port map (
            O => \N__40679\,
            I => \N__40675\
        );

    \I__8748\ : InMux
    port map (
            O => \N__40678\,
            I => \N__40672\
        );

    \I__8747\ : InMux
    port map (
            O => \N__40675\,
            I => \N__40667\
        );

    \I__8746\ : LocalMux
    port map (
            O => \N__40672\,
            I => \N__40664\
        );

    \I__8745\ : InMux
    port map (
            O => \N__40671\,
            I => \N__40659\
        );

    \I__8744\ : InMux
    port map (
            O => \N__40670\,
            I => \N__40659\
        );

    \I__8743\ : LocalMux
    port map (
            O => \N__40667\,
            I => \N__40656\
        );

    \I__8742\ : Span4Mux_h
    port map (
            O => \N__40664\,
            I => \N__40651\
        );

    \I__8741\ : LocalMux
    port map (
            O => \N__40659\,
            I => \N__40651\
        );

    \I__8740\ : Span4Mux_h
    port map (
            O => \N__40656\,
            I => \N__40648\
        );

    \I__8739\ : Odrv4
    port map (
            O => \N__40651\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__8738\ : Odrv4
    port map (
            O => \N__40648\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__8737\ : CascadeMux
    port map (
            O => \N__40643\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25_cascade_\
        );

    \I__8736\ : CascadeMux
    port map (
            O => \N__40640\,
            I => \N__40636\
        );

    \I__8735\ : InMux
    port map (
            O => \N__40639\,
            I => \N__40631\
        );

    \I__8734\ : InMux
    port map (
            O => \N__40636\,
            I => \N__40631\
        );

    \I__8733\ : LocalMux
    port map (
            O => \N__40631\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\
        );

    \I__8732\ : InMux
    port map (
            O => \N__40628\,
            I => \N__40623\
        );

    \I__8731\ : CascadeMux
    port map (
            O => \N__40627\,
            I => \N__40619\
        );

    \I__8730\ : InMux
    port map (
            O => \N__40626\,
            I => \N__40616\
        );

    \I__8729\ : LocalMux
    port map (
            O => \N__40623\,
            I => \N__40613\
        );

    \I__8728\ : InMux
    port map (
            O => \N__40622\,
            I => \N__40610\
        );

    \I__8727\ : InMux
    port map (
            O => \N__40619\,
            I => \N__40607\
        );

    \I__8726\ : LocalMux
    port map (
            O => \N__40616\,
            I => \N__40604\
        );

    \I__8725\ : Span4Mux_h
    port map (
            O => \N__40613\,
            I => \N__40601\
        );

    \I__8724\ : LocalMux
    port map (
            O => \N__40610\,
            I => \N__40598\
        );

    \I__8723\ : LocalMux
    port map (
            O => \N__40607\,
            I => \N__40595\
        );

    \I__8722\ : Odrv4
    port map (
            O => \N__40604\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__8721\ : Odrv4
    port map (
            O => \N__40601\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__8720\ : Odrv4
    port map (
            O => \N__40598\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__8719\ : Odrv4
    port map (
            O => \N__40595\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__8718\ : InMux
    port map (
            O => \N__40586\,
            I => \N__40583\
        );

    \I__8717\ : LocalMux
    port map (
            O => \N__40583\,
            I => \N__40579\
        );

    \I__8716\ : InMux
    port map (
            O => \N__40582\,
            I => \N__40575\
        );

    \I__8715\ : Span4Mux_v
    port map (
            O => \N__40579\,
            I => \N__40572\
        );

    \I__8714\ : InMux
    port map (
            O => \N__40578\,
            I => \N__40569\
        );

    \I__8713\ : LocalMux
    port map (
            O => \N__40575\,
            I => \N__40566\
        );

    \I__8712\ : Span4Mux_h
    port map (
            O => \N__40572\,
            I => \N__40563\
        );

    \I__8711\ : LocalMux
    port map (
            O => \N__40569\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24\
        );

    \I__8710\ : Odrv12
    port map (
            O => \N__40566\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24\
        );

    \I__8709\ : Odrv4
    port map (
            O => \N__40563\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24\
        );

    \I__8708\ : InMux
    port map (
            O => \N__40556\,
            I => \N__40550\
        );

    \I__8707\ : InMux
    port map (
            O => \N__40555\,
            I => \N__40550\
        );

    \I__8706\ : LocalMux
    port map (
            O => \N__40550\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\
        );

    \I__8705\ : CascadeMux
    port map (
            O => \N__40547\,
            I => \N__40544\
        );

    \I__8704\ : InMux
    port map (
            O => \N__40544\,
            I => \N__40541\
        );

    \I__8703\ : LocalMux
    port map (
            O => \N__40541\,
            I => \N__40538\
        );

    \I__8702\ : Span4Mux_h
    port map (
            O => \N__40538\,
            I => \N__40535\
        );

    \I__8701\ : Odrv4
    port map (
            O => \N__40535\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\
        );

    \I__8700\ : InMux
    port map (
            O => \N__40532\,
            I => \N__40529\
        );

    \I__8699\ : LocalMux
    port map (
            O => \N__40529\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\
        );

    \I__8698\ : CascadeMux
    port map (
            O => \N__40526\,
            I => \N__40523\
        );

    \I__8697\ : InMux
    port map (
            O => \N__40523\,
            I => \N__40520\
        );

    \I__8696\ : LocalMux
    port map (
            O => \N__40520\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\
        );

    \I__8695\ : CascadeMux
    port map (
            O => \N__40517\,
            I => \N__40514\
        );

    \I__8694\ : InMux
    port map (
            O => \N__40514\,
            I => \N__40511\
        );

    \I__8693\ : LocalMux
    port map (
            O => \N__40511\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\
        );

    \I__8692\ : CascadeMux
    port map (
            O => \N__40508\,
            I => \N__40505\
        );

    \I__8691\ : InMux
    port map (
            O => \N__40505\,
            I => \N__40502\
        );

    \I__8690\ : LocalMux
    port map (
            O => \N__40502\,
            I => \N__40499\
        );

    \I__8689\ : Odrv4
    port map (
            O => \N__40499\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\
        );

    \I__8688\ : InMux
    port map (
            O => \N__40496\,
            I => \N__40493\
        );

    \I__8687\ : LocalMux
    port map (
            O => \N__40493\,
            I => \N__40490\
        );

    \I__8686\ : Span4Mux_v
    port map (
            O => \N__40490\,
            I => \N__40487\
        );

    \I__8685\ : Odrv4
    port map (
            O => \N__40487\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\
        );

    \I__8684\ : CascadeMux
    port map (
            O => \N__40484\,
            I => \N__40481\
        );

    \I__8683\ : InMux
    port map (
            O => \N__40481\,
            I => \N__40478\
        );

    \I__8682\ : LocalMux
    port map (
            O => \N__40478\,
            I => \N__40475\
        );

    \I__8681\ : Odrv4
    port map (
            O => \N__40475\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\
        );

    \I__8680\ : CascadeMux
    port map (
            O => \N__40472\,
            I => \N__40469\
        );

    \I__8679\ : InMux
    port map (
            O => \N__40469\,
            I => \N__40466\
        );

    \I__8678\ : LocalMux
    port map (
            O => \N__40466\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\
        );

    \I__8677\ : InMux
    port map (
            O => \N__40463\,
            I => \N__40460\
        );

    \I__8676\ : LocalMux
    port map (
            O => \N__40460\,
            I => \N__40457\
        );

    \I__8675\ : Span4Mux_h
    port map (
            O => \N__40457\,
            I => \N__40454\
        );

    \I__8674\ : Odrv4
    port map (
            O => \N__40454\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\
        );

    \I__8673\ : CascadeMux
    port map (
            O => \N__40451\,
            I => \N__40448\
        );

    \I__8672\ : InMux
    port map (
            O => \N__40448\,
            I => \N__40445\
        );

    \I__8671\ : LocalMux
    port map (
            O => \N__40445\,
            I => \N__40442\
        );

    \I__8670\ : Odrv12
    port map (
            O => \N__40442\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\
        );

    \I__8669\ : InMux
    port map (
            O => \N__40439\,
            I => \N__40436\
        );

    \I__8668\ : LocalMux
    port map (
            O => \N__40436\,
            I => \N__40433\
        );

    \I__8667\ : Span4Mux_h
    port map (
            O => \N__40433\,
            I => \N__40430\
        );

    \I__8666\ : Odrv4
    port map (
            O => \N__40430\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\
        );

    \I__8665\ : CascadeMux
    port map (
            O => \N__40427\,
            I => \N__40424\
        );

    \I__8664\ : InMux
    port map (
            O => \N__40424\,
            I => \N__40421\
        );

    \I__8663\ : LocalMux
    port map (
            O => \N__40421\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\
        );

    \I__8662\ : InMux
    port map (
            O => \N__40418\,
            I => \N__40415\
        );

    \I__8661\ : LocalMux
    port map (
            O => \N__40415\,
            I => \N__40412\
        );

    \I__8660\ : Span4Mux_v
    port map (
            O => \N__40412\,
            I => \N__40409\
        );

    \I__8659\ : Odrv4
    port map (
            O => \N__40409\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\
        );

    \I__8658\ : CascadeMux
    port map (
            O => \N__40406\,
            I => \N__40403\
        );

    \I__8657\ : InMux
    port map (
            O => \N__40403\,
            I => \N__40400\
        );

    \I__8656\ : LocalMux
    port map (
            O => \N__40400\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\
        );

    \I__8655\ : InMux
    port map (
            O => \N__40397\,
            I => \N__40394\
        );

    \I__8654\ : LocalMux
    port map (
            O => \N__40394\,
            I => \N__40391\
        );

    \I__8653\ : Span4Mux_h
    port map (
            O => \N__40391\,
            I => \N__40388\
        );

    \I__8652\ : Odrv4
    port map (
            O => \N__40388\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\
        );

    \I__8651\ : CascadeMux
    port map (
            O => \N__40385\,
            I => \N__40382\
        );

    \I__8650\ : InMux
    port map (
            O => \N__40382\,
            I => \N__40379\
        );

    \I__8649\ : LocalMux
    port map (
            O => \N__40379\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\
        );

    \I__8648\ : InMux
    port map (
            O => \N__40376\,
            I => \N__40373\
        );

    \I__8647\ : LocalMux
    port map (
            O => \N__40373\,
            I => \N__40370\
        );

    \I__8646\ : Odrv12
    port map (
            O => \N__40370\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\
        );

    \I__8645\ : CascadeMux
    port map (
            O => \N__40367\,
            I => \N__40364\
        );

    \I__8644\ : InMux
    port map (
            O => \N__40364\,
            I => \N__40361\
        );

    \I__8643\ : LocalMux
    port map (
            O => \N__40361\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\
        );

    \I__8642\ : InMux
    port map (
            O => \N__40358\,
            I => \N__40352\
        );

    \I__8641\ : InMux
    port map (
            O => \N__40357\,
            I => \N__40352\
        );

    \I__8640\ : LocalMux
    port map (
            O => \N__40352\,
            I => \N__40349\
        );

    \I__8639\ : Span4Mux_v
    port map (
            O => \N__40349\,
            I => \N__40346\
        );

    \I__8638\ : Odrv4
    port map (
            O => \N__40346\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_30\
        );

    \I__8637\ : InMux
    port map (
            O => \N__40343\,
            I => \N__40337\
        );

    \I__8636\ : InMux
    port map (
            O => \N__40342\,
            I => \N__40337\
        );

    \I__8635\ : LocalMux
    port map (
            O => \N__40337\,
            I => \N__40334\
        );

    \I__8634\ : Odrv12
    port map (
            O => \N__40334\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_31\
        );

    \I__8633\ : InMux
    port map (
            O => \N__40331\,
            I => \N__40328\
        );

    \I__8632\ : LocalMux
    port map (
            O => \N__40328\,
            I => \N__40325\
        );

    \I__8631\ : Span4Mux_h
    port map (
            O => \N__40325\,
            I => \N__40319\
        );

    \I__8630\ : InMux
    port map (
            O => \N__40324\,
            I => \N__40316\
        );

    \I__8629\ : InMux
    port map (
            O => \N__40323\,
            I => \N__40313\
        );

    \I__8628\ : InMux
    port map (
            O => \N__40322\,
            I => \N__40310\
        );

    \I__8627\ : Odrv4
    port map (
            O => \N__40319\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__8626\ : LocalMux
    port map (
            O => \N__40316\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__8625\ : LocalMux
    port map (
            O => \N__40313\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__8624\ : LocalMux
    port map (
            O => \N__40310\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__8623\ : InMux
    port map (
            O => \N__40301\,
            I => \N__40298\
        );

    \I__8622\ : LocalMux
    port map (
            O => \N__40298\,
            I => \N__40294\
        );

    \I__8621\ : InMux
    port map (
            O => \N__40297\,
            I => \N__40290\
        );

    \I__8620\ : Span4Mux_v
    port map (
            O => \N__40294\,
            I => \N__40287\
        );

    \I__8619\ : InMux
    port map (
            O => \N__40293\,
            I => \N__40284\
        );

    \I__8618\ : LocalMux
    port map (
            O => \N__40290\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5\
        );

    \I__8617\ : Odrv4
    port map (
            O => \N__40287\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5\
        );

    \I__8616\ : LocalMux
    port map (
            O => \N__40284\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5\
        );

    \I__8615\ : InMux
    port map (
            O => \N__40277\,
            I => \N__40272\
        );

    \I__8614\ : InMux
    port map (
            O => \N__40276\,
            I => \N__40269\
        );

    \I__8613\ : InMux
    port map (
            O => \N__40275\,
            I => \N__40266\
        );

    \I__8612\ : LocalMux
    port map (
            O => \N__40272\,
            I => \N__40262\
        );

    \I__8611\ : LocalMux
    port map (
            O => \N__40269\,
            I => \N__40259\
        );

    \I__8610\ : LocalMux
    port map (
            O => \N__40266\,
            I => \N__40256\
        );

    \I__8609\ : InMux
    port map (
            O => \N__40265\,
            I => \N__40253\
        );

    \I__8608\ : Span4Mux_v
    port map (
            O => \N__40262\,
            I => \N__40250\
        );

    \I__8607\ : Span4Mux_h
    port map (
            O => \N__40259\,
            I => \N__40247\
        );

    \I__8606\ : Span4Mux_v
    port map (
            O => \N__40256\,
            I => \N__40244\
        );

    \I__8605\ : LocalMux
    port map (
            O => \N__40253\,
            I => \N__40241\
        );

    \I__8604\ : Odrv4
    port map (
            O => \N__40250\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__8603\ : Odrv4
    port map (
            O => \N__40247\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__8602\ : Odrv4
    port map (
            O => \N__40244\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__8601\ : Odrv4
    port map (
            O => \N__40241\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__8600\ : InMux
    port map (
            O => \N__40232\,
            I => \N__40229\
        );

    \I__8599\ : LocalMux
    port map (
            O => \N__40229\,
            I => \N__40226\
        );

    \I__8598\ : Span4Mux_v
    port map (
            O => \N__40226\,
            I => \N__40223\
        );

    \I__8597\ : Odrv4
    port map (
            O => \N__40223\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\
        );

    \I__8596\ : CascadeMux
    port map (
            O => \N__40220\,
            I => \N__40217\
        );

    \I__8595\ : InMux
    port map (
            O => \N__40217\,
            I => \N__40214\
        );

    \I__8594\ : LocalMux
    port map (
            O => \N__40214\,
            I => \N__40211\
        );

    \I__8593\ : Odrv4
    port map (
            O => \N__40211\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\
        );

    \I__8592\ : CascadeMux
    port map (
            O => \N__40208\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\
        );

    \I__8591\ : CascadeMux
    port map (
            O => \N__40205\,
            I => \N__40202\
        );

    \I__8590\ : InMux
    port map (
            O => \N__40202\,
            I => \N__40199\
        );

    \I__8589\ : LocalMux
    port map (
            O => \N__40199\,
            I => \N__40196\
        );

    \I__8588\ : Odrv4
    port map (
            O => \N__40196\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\
        );

    \I__8587\ : InMux
    port map (
            O => \N__40193\,
            I => \N__40190\
        );

    \I__8586\ : LocalMux
    port map (
            O => \N__40190\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\
        );

    \I__8585\ : InMux
    port map (
            O => \N__40187\,
            I => \N__40184\
        );

    \I__8584\ : LocalMux
    port map (
            O => \N__40184\,
            I => \N__40181\
        );

    \I__8583\ : Odrv4
    port map (
            O => \N__40181\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\
        );

    \I__8582\ : CascadeMux
    port map (
            O => \N__40178\,
            I => \N__40175\
        );

    \I__8581\ : InMux
    port map (
            O => \N__40175\,
            I => \N__40172\
        );

    \I__8580\ : LocalMux
    port map (
            O => \N__40172\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\
        );

    \I__8579\ : InMux
    port map (
            O => \N__40169\,
            I => \N__40166\
        );

    \I__8578\ : LocalMux
    port map (
            O => \N__40166\,
            I => \N__40163\
        );

    \I__8577\ : Odrv4
    port map (
            O => \N__40163\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\
        );

    \I__8576\ : CascadeMux
    port map (
            O => \N__40160\,
            I => \N__40157\
        );

    \I__8575\ : InMux
    port map (
            O => \N__40157\,
            I => \N__40154\
        );

    \I__8574\ : LocalMux
    port map (
            O => \N__40154\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\
        );

    \I__8573\ : CascadeMux
    port map (
            O => \N__40151\,
            I => \N__40148\
        );

    \I__8572\ : InMux
    port map (
            O => \N__40148\,
            I => \N__40145\
        );

    \I__8571\ : LocalMux
    port map (
            O => \N__40145\,
            I => \N__40142\
        );

    \I__8570\ : Odrv4
    port map (
            O => \N__40142\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\
        );

    \I__8569\ : InMux
    port map (
            O => \N__40139\,
            I => \N__40136\
        );

    \I__8568\ : LocalMux
    port map (
            O => \N__40136\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\
        );

    \I__8567\ : InMux
    port map (
            O => \N__40133\,
            I => \N__40130\
        );

    \I__8566\ : LocalMux
    port map (
            O => \N__40130\,
            I => \N__40127\
        );

    \I__8565\ : Odrv4
    port map (
            O => \N__40127\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\
        );

    \I__8564\ : InMux
    port map (
            O => \N__40124\,
            I => \N__40121\
        );

    \I__8563\ : LocalMux
    port map (
            O => \N__40121\,
            I => \N__40115\
        );

    \I__8562\ : InMux
    port map (
            O => \N__40120\,
            I => \N__40112\
        );

    \I__8561\ : InMux
    port map (
            O => \N__40119\,
            I => \N__40109\
        );

    \I__8560\ : InMux
    port map (
            O => \N__40118\,
            I => \N__40106\
        );

    \I__8559\ : Odrv4
    port map (
            O => \N__40115\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__8558\ : LocalMux
    port map (
            O => \N__40112\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__8557\ : LocalMux
    port map (
            O => \N__40109\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__8556\ : LocalMux
    port map (
            O => \N__40106\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__8555\ : InMux
    port map (
            O => \N__40097\,
            I => \N__40094\
        );

    \I__8554\ : LocalMux
    port map (
            O => \N__40094\,
            I => \N__40090\
        );

    \I__8553\ : InMux
    port map (
            O => \N__40093\,
            I => \N__40086\
        );

    \I__8552\ : Span4Mux_h
    port map (
            O => \N__40090\,
            I => \N__40083\
        );

    \I__8551\ : InMux
    port map (
            O => \N__40089\,
            I => \N__40080\
        );

    \I__8550\ : LocalMux
    port map (
            O => \N__40086\,
            I => \elapsed_time_ns_1_RNIK63T9_0_8\
        );

    \I__8549\ : Odrv4
    port map (
            O => \N__40083\,
            I => \elapsed_time_ns_1_RNIK63T9_0_8\
        );

    \I__8548\ : LocalMux
    port map (
            O => \N__40080\,
            I => \elapsed_time_ns_1_RNIK63T9_0_8\
        );

    \I__8547\ : InMux
    port map (
            O => \N__40073\,
            I => \N__40069\
        );

    \I__8546\ : InMux
    port map (
            O => \N__40072\,
            I => \N__40066\
        );

    \I__8545\ : LocalMux
    port map (
            O => \N__40069\,
            I => \N__40061\
        );

    \I__8544\ : LocalMux
    port map (
            O => \N__40066\,
            I => \N__40058\
        );

    \I__8543\ : InMux
    port map (
            O => \N__40065\,
            I => \N__40055\
        );

    \I__8542\ : InMux
    port map (
            O => \N__40064\,
            I => \N__40052\
        );

    \I__8541\ : Odrv4
    port map (
            O => \N__40061\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__8540\ : Odrv4
    port map (
            O => \N__40058\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__8539\ : LocalMux
    port map (
            O => \N__40055\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__8538\ : LocalMux
    port map (
            O => \N__40052\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__8537\ : InMux
    port map (
            O => \N__40043\,
            I => \N__40040\
        );

    \I__8536\ : LocalMux
    port map (
            O => \N__40040\,
            I => \N__40036\
        );

    \I__8535\ : InMux
    port map (
            O => \N__40039\,
            I => \N__40032\
        );

    \I__8534\ : Span4Mux_h
    port map (
            O => \N__40036\,
            I => \N__40029\
        );

    \I__8533\ : InMux
    port map (
            O => \N__40035\,
            I => \N__40026\
        );

    \I__8532\ : LocalMux
    port map (
            O => \N__40032\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12\
        );

    \I__8531\ : Odrv4
    port map (
            O => \N__40029\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12\
        );

    \I__8530\ : LocalMux
    port map (
            O => \N__40026\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12\
        );

    \I__8529\ : InMux
    port map (
            O => \N__40019\,
            I => \N__40016\
        );

    \I__8528\ : LocalMux
    port map (
            O => \N__40016\,
            I => \N__40013\
        );

    \I__8527\ : Odrv12
    port map (
            O => \N__40013\,
            I => \current_shift_inst.un4_control_input_1_axb_19\
        );

    \I__8526\ : InMux
    port map (
            O => \N__40010\,
            I => \N__40003\
        );

    \I__8525\ : InMux
    port map (
            O => \N__40009\,
            I => \N__40003\
        );

    \I__8524\ : InMux
    port map (
            O => \N__40008\,
            I => \N__39999\
        );

    \I__8523\ : LocalMux
    port map (
            O => \N__40003\,
            I => \N__39996\
        );

    \I__8522\ : InMux
    port map (
            O => \N__40002\,
            I => \N__39993\
        );

    \I__8521\ : LocalMux
    port map (
            O => \N__39999\,
            I => \N__39990\
        );

    \I__8520\ : Span4Mux_h
    port map (
            O => \N__39996\,
            I => \N__39985\
        );

    \I__8519\ : LocalMux
    port map (
            O => \N__39993\,
            I => \N__39985\
        );

    \I__8518\ : Odrv4
    port map (
            O => \N__39990\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__8517\ : Odrv4
    port map (
            O => \N__39985\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__8516\ : CascadeMux
    port map (
            O => \N__39980\,
            I => \N__39975\
        );

    \I__8515\ : InMux
    port map (
            O => \N__39979\,
            I => \N__39972\
        );

    \I__8514\ : InMux
    port map (
            O => \N__39978\,
            I => \N__39967\
        );

    \I__8513\ : InMux
    port map (
            O => \N__39975\,
            I => \N__39967\
        );

    \I__8512\ : LocalMux
    port map (
            O => \N__39972\,
            I => \N__39964\
        );

    \I__8511\ : LocalMux
    port map (
            O => \N__39967\,
            I => \N__39961\
        );

    \I__8510\ : Span4Mux_v
    port map (
            O => \N__39964\,
            I => \N__39958\
        );

    \I__8509\ : Odrv4
    port map (
            O => \N__39961\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__8508\ : Odrv4
    port map (
            O => \N__39958\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__8507\ : CascadeMux
    port map (
            O => \N__39953\,
            I => \N__39950\
        );

    \I__8506\ : InMux
    port map (
            O => \N__39950\,
            I => \N__39946\
        );

    \I__8505\ : InMux
    port map (
            O => \N__39949\,
            I => \N__39943\
        );

    \I__8504\ : LocalMux
    port map (
            O => \N__39946\,
            I => \N__39940\
        );

    \I__8503\ : LocalMux
    port map (
            O => \N__39943\,
            I => \N__39935\
        );

    \I__8502\ : Span4Mux_h
    port map (
            O => \N__39940\,
            I => \N__39932\
        );

    \I__8501\ : InMux
    port map (
            O => \N__39939\,
            I => \N__39929\
        );

    \I__8500\ : InMux
    port map (
            O => \N__39938\,
            I => \N__39926\
        );

    \I__8499\ : Span4Mux_h
    port map (
            O => \N__39935\,
            I => \N__39923\
        );

    \I__8498\ : Span4Mux_v
    port map (
            O => \N__39932\,
            I => \N__39920\
        );

    \I__8497\ : LocalMux
    port map (
            O => \N__39929\,
            I => \N__39915\
        );

    \I__8496\ : LocalMux
    port map (
            O => \N__39926\,
            I => \N__39915\
        );

    \I__8495\ : Odrv4
    port map (
            O => \N__39923\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__8494\ : Odrv4
    port map (
            O => \N__39920\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__8493\ : Odrv12
    port map (
            O => \N__39915\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__8492\ : InMux
    port map (
            O => \N__39908\,
            I => \N__39905\
        );

    \I__8491\ : LocalMux
    port map (
            O => \N__39905\,
            I => \N__39900\
        );

    \I__8490\ : InMux
    port map (
            O => \N__39904\,
            I => \N__39897\
        );

    \I__8489\ : InMux
    port map (
            O => \N__39903\,
            I => \N__39894\
        );

    \I__8488\ : Span4Mux_v
    port map (
            O => \N__39900\,
            I => \N__39891\
        );

    \I__8487\ : LocalMux
    port map (
            O => \N__39897\,
            I => \N__39886\
        );

    \I__8486\ : LocalMux
    port map (
            O => \N__39894\,
            I => \N__39886\
        );

    \I__8485\ : Odrv4
    port map (
            O => \N__39891\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__8484\ : Odrv12
    port map (
            O => \N__39886\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__8483\ : CascadeMux
    port map (
            O => \N__39881\,
            I => \N__39878\
        );

    \I__8482\ : InMux
    port map (
            O => \N__39878\,
            I => \N__39875\
        );

    \I__8481\ : LocalMux
    port map (
            O => \N__39875\,
            I => \N__39872\
        );

    \I__8480\ : Span4Mux_h
    port map (
            O => \N__39872\,
            I => \N__39869\
        );

    \I__8479\ : Span4Mux_v
    port map (
            O => \N__39869\,
            I => \N__39866\
        );

    \I__8478\ : Odrv4
    port map (
            O => \N__39866\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISST11_17\
        );

    \I__8477\ : InMux
    port map (
            O => \N__39863\,
            I => \N__39860\
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__39860\,
            I => \N__39857\
        );

    \I__8475\ : Span4Mux_s1_v
    port map (
            O => \N__39857\,
            I => \N__39853\
        );

    \I__8474\ : InMux
    port map (
            O => \N__39856\,
            I => \N__39850\
        );

    \I__8473\ : Span4Mux_h
    port map (
            O => \N__39853\,
            I => \N__39847\
        );

    \I__8472\ : LocalMux
    port map (
            O => \N__39850\,
            I => \N__39840\
        );

    \I__8471\ : Sp12to4
    port map (
            O => \N__39847\,
            I => \N__39840\
        );

    \I__8470\ : InMux
    port map (
            O => \N__39846\,
            I => \N__39836\
        );

    \I__8469\ : InMux
    port map (
            O => \N__39845\,
            I => \N__39833\
        );

    \I__8468\ : Span12Mux_s10_v
    port map (
            O => \N__39840\,
            I => \N__39830\
        );

    \I__8467\ : InMux
    port map (
            O => \N__39839\,
            I => \N__39827\
        );

    \I__8466\ : LocalMux
    port map (
            O => \N__39836\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__8465\ : LocalMux
    port map (
            O => \N__39833\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__8464\ : Odrv12
    port map (
            O => \N__39830\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__8463\ : LocalMux
    port map (
            O => \N__39827\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__8462\ : IoInMux
    port map (
            O => \N__39818\,
            I => \N__39815\
        );

    \I__8461\ : LocalMux
    port map (
            O => \N__39815\,
            I => \N__39812\
        );

    \I__8460\ : Span4Mux_s0_v
    port map (
            O => \N__39812\,
            I => \N__39808\
        );

    \I__8459\ : InMux
    port map (
            O => \N__39811\,
            I => \N__39805\
        );

    \I__8458\ : Odrv4
    port map (
            O => \N__39808\,
            I => \T23_c\
        );

    \I__8457\ : LocalMux
    port map (
            O => \N__39805\,
            I => \T23_c\
        );

    \I__8456\ : InMux
    port map (
            O => \N__39800\,
            I => \N__39796\
        );

    \I__8455\ : InMux
    port map (
            O => \N__39799\,
            I => \N__39793\
        );

    \I__8454\ : LocalMux
    port map (
            O => \N__39796\,
            I => \N__39789\
        );

    \I__8453\ : LocalMux
    port map (
            O => \N__39793\,
            I => \N__39786\
        );

    \I__8452\ : InMux
    port map (
            O => \N__39792\,
            I => \N__39783\
        );

    \I__8451\ : Span4Mux_h
    port map (
            O => \N__39789\,
            I => \N__39780\
        );

    \I__8450\ : Span4Mux_v
    port map (
            O => \N__39786\,
            I => \N__39777\
        );

    \I__8449\ : LocalMux
    port map (
            O => \N__39783\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21\
        );

    \I__8448\ : Odrv4
    port map (
            O => \N__39780\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21\
        );

    \I__8447\ : Odrv4
    port map (
            O => \N__39777\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21\
        );

    \I__8446\ : InMux
    port map (
            O => \N__39770\,
            I => \N__39764\
        );

    \I__8445\ : InMux
    port map (
            O => \N__39769\,
            I => \N__39761\
        );

    \I__8444\ : InMux
    port map (
            O => \N__39768\,
            I => \N__39758\
        );

    \I__8443\ : InMux
    port map (
            O => \N__39767\,
            I => \N__39755\
        );

    \I__8442\ : LocalMux
    port map (
            O => \N__39764\,
            I => \N__39752\
        );

    \I__8441\ : LocalMux
    port map (
            O => \N__39761\,
            I => \N__39747\
        );

    \I__8440\ : LocalMux
    port map (
            O => \N__39758\,
            I => \N__39747\
        );

    \I__8439\ : LocalMux
    port map (
            O => \N__39755\,
            I => \N__39744\
        );

    \I__8438\ : Span4Mux_h
    port map (
            O => \N__39752\,
            I => \N__39739\
        );

    \I__8437\ : Span4Mux_v
    port map (
            O => \N__39747\,
            I => \N__39739\
        );

    \I__8436\ : Span4Mux_v
    port map (
            O => \N__39744\,
            I => \N__39736\
        );

    \I__8435\ : Odrv4
    port map (
            O => \N__39739\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__8434\ : Odrv4
    port map (
            O => \N__39736\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__8433\ : InMux
    port map (
            O => \N__39731\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\
        );

    \I__8432\ : InMux
    port map (
            O => \N__39728\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\
        );

    \I__8431\ : InMux
    port map (
            O => \N__39725\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\
        );

    \I__8430\ : InMux
    port map (
            O => \N__39722\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\
        );

    \I__8429\ : InMux
    port map (
            O => \N__39719\,
            I => \N__39716\
        );

    \I__8428\ : LocalMux
    port map (
            O => \N__39716\,
            I => \N__39713\
        );

    \I__8427\ : Odrv12
    port map (
            O => \N__39713\,
            I => \current_shift_inst.un4_control_input_1_axb_27\
        );

    \I__8426\ : CascadeMux
    port map (
            O => \N__39710\,
            I => \N__39707\
        );

    \I__8425\ : InMux
    port map (
            O => \N__39707\,
            I => \N__39704\
        );

    \I__8424\ : LocalMux
    port map (
            O => \N__39704\,
            I => \N__39701\
        );

    \I__8423\ : Span4Mux_h
    port map (
            O => \N__39701\,
            I => \N__39696\
        );

    \I__8422\ : InMux
    port map (
            O => \N__39700\,
            I => \N__39691\
        );

    \I__8421\ : InMux
    port map (
            O => \N__39699\,
            I => \N__39691\
        );

    \I__8420\ : Span4Mux_v
    port map (
            O => \N__39696\,
            I => \N__39687\
        );

    \I__8419\ : LocalMux
    port map (
            O => \N__39691\,
            I => \N__39684\
        );

    \I__8418\ : InMux
    port map (
            O => \N__39690\,
            I => \N__39681\
        );

    \I__8417\ : Odrv4
    port map (
            O => \N__39687\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__8416\ : Odrv4
    port map (
            O => \N__39684\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__8415\ : LocalMux
    port map (
            O => \N__39681\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__8414\ : InMux
    port map (
            O => \N__39674\,
            I => \N__39671\
        );

    \I__8413\ : LocalMux
    port map (
            O => \N__39671\,
            I => \N__39668\
        );

    \I__8412\ : Odrv12
    port map (
            O => \N__39668\,
            I => \current_shift_inst.un4_control_input_1_axb_28\
        );

    \I__8411\ : InMux
    port map (
            O => \N__39665\,
            I => \N__39662\
        );

    \I__8410\ : LocalMux
    port map (
            O => \N__39662\,
            I => \N__39659\
        );

    \I__8409\ : Odrv12
    port map (
            O => \N__39659\,
            I => \current_shift_inst.un4_control_input_1_axb_29\
        );

    \I__8408\ : InMux
    port map (
            O => \N__39656\,
            I => \N__39652\
        );

    \I__8407\ : CascadeMux
    port map (
            O => \N__39655\,
            I => \N__39649\
        );

    \I__8406\ : LocalMux
    port map (
            O => \N__39652\,
            I => \N__39646\
        );

    \I__8405\ : InMux
    port map (
            O => \N__39649\,
            I => \N__39643\
        );

    \I__8404\ : Span4Mux_h
    port map (
            O => \N__39646\,
            I => \N__39636\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__39643\,
            I => \N__39636\
        );

    \I__8402\ : InMux
    port map (
            O => \N__39642\,
            I => \N__39633\
        );

    \I__8401\ : InMux
    port map (
            O => \N__39641\,
            I => \N__39630\
        );

    \I__8400\ : Odrv4
    port map (
            O => \N__39636\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__8399\ : LocalMux
    port map (
            O => \N__39633\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__8398\ : LocalMux
    port map (
            O => \N__39630\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__8397\ : InMux
    port map (
            O => \N__39623\,
            I => \N__39620\
        );

    \I__8396\ : LocalMux
    port map (
            O => \N__39620\,
            I => \N__39615\
        );

    \I__8395\ : InMux
    port map (
            O => \N__39619\,
            I => \N__39612\
        );

    \I__8394\ : InMux
    port map (
            O => \N__39618\,
            I => \N__39609\
        );

    \I__8393\ : Span4Mux_v
    port map (
            O => \N__39615\,
            I => \N__39606\
        );

    \I__8392\ : LocalMux
    port map (
            O => \N__39612\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__8391\ : LocalMux
    port map (
            O => \N__39609\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__8390\ : Odrv4
    port map (
            O => \N__39606\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__8389\ : InMux
    port map (
            O => \N__39599\,
            I => \N__39594\
        );

    \I__8388\ : InMux
    port map (
            O => \N__39598\,
            I => \N__39591\
        );

    \I__8387\ : InMux
    port map (
            O => \N__39597\,
            I => \N__39588\
        );

    \I__8386\ : LocalMux
    port map (
            O => \N__39594\,
            I => \N__39585\
        );

    \I__8385\ : LocalMux
    port map (
            O => \N__39591\,
            I => \N__39582\
        );

    \I__8384\ : LocalMux
    port map (
            O => \N__39588\,
            I => \N__39579\
        );

    \I__8383\ : Span4Mux_h
    port map (
            O => \N__39585\,
            I => \N__39576\
        );

    \I__8382\ : Span4Mux_v
    port map (
            O => \N__39582\,
            I => \N__39573\
        );

    \I__8381\ : Odrv4
    port map (
            O => \N__39579\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__8380\ : Odrv4
    port map (
            O => \N__39576\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__8379\ : Odrv4
    port map (
            O => \N__39573\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__8378\ : InMux
    port map (
            O => \N__39566\,
            I => \bfn_16_21_0_\
        );

    \I__8377\ : InMux
    port map (
            O => \N__39563\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\
        );

    \I__8376\ : InMux
    port map (
            O => \N__39560\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\
        );

    \I__8375\ : InMux
    port map (
            O => \N__39557\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\
        );

    \I__8374\ : InMux
    port map (
            O => \N__39554\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\
        );

    \I__8373\ : InMux
    port map (
            O => \N__39551\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\
        );

    \I__8372\ : InMux
    port map (
            O => \N__39548\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\
        );

    \I__8371\ : InMux
    port map (
            O => \N__39545\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\
        );

    \I__8370\ : InMux
    port map (
            O => \N__39542\,
            I => \bfn_16_22_0_\
        );

    \I__8369\ : InMux
    port map (
            O => \N__39539\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\
        );

    \I__8368\ : InMux
    port map (
            O => \N__39536\,
            I => \bfn_16_20_0_\
        );

    \I__8367\ : InMux
    port map (
            O => \N__39533\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\
        );

    \I__8366\ : InMux
    port map (
            O => \N__39530\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\
        );

    \I__8365\ : InMux
    port map (
            O => \N__39527\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\
        );

    \I__8364\ : InMux
    port map (
            O => \N__39524\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\
        );

    \I__8363\ : InMux
    port map (
            O => \N__39521\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\
        );

    \I__8362\ : InMux
    port map (
            O => \N__39518\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\
        );

    \I__8361\ : InMux
    port map (
            O => \N__39515\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\
        );

    \I__8360\ : InMux
    port map (
            O => \N__39512\,
            I => \current_shift_inst.un4_control_input1_31\
        );

    \I__8359\ : InMux
    port map (
            O => \N__39509\,
            I => \N__39506\
        );

    \I__8358\ : LocalMux
    port map (
            O => \N__39506\,
            I => \N__39503\
        );

    \I__8357\ : Odrv12
    port map (
            O => \N__39503\,
            I => \current_shift_inst.un4_control_input_1_axb_2\
        );

    \I__8356\ : InMux
    port map (
            O => \N__39500\,
            I => \N__39497\
        );

    \I__8355\ : LocalMux
    port map (
            O => \N__39497\,
            I => \current_shift_inst.un4_control_input_1_axb_24\
        );

    \I__8354\ : InMux
    port map (
            O => \N__39494\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\
        );

    \I__8353\ : InMux
    port map (
            O => \N__39491\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\
        );

    \I__8352\ : InMux
    port map (
            O => \N__39488\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\
        );

    \I__8351\ : InMux
    port map (
            O => \N__39485\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\
        );

    \I__8350\ : InMux
    port map (
            O => \N__39482\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\
        );

    \I__8349\ : InMux
    port map (
            O => \N__39479\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\
        );

    \I__8348\ : InMux
    port map (
            O => \N__39476\,
            I => \N__39473\
        );

    \I__8347\ : LocalMux
    port map (
            O => \N__39473\,
            I => \current_shift_inst.un4_control_input_1_axb_22\
        );

    \I__8346\ : InMux
    port map (
            O => \N__39470\,
            I => \current_shift_inst.un4_control_input_1_cry_21\
        );

    \I__8345\ : InMux
    port map (
            O => \N__39467\,
            I => \current_shift_inst.un4_control_input_1_cry_22\
        );

    \I__8344\ : InMux
    port map (
            O => \N__39464\,
            I => \current_shift_inst.un4_control_input_1_cry_23\
        );

    \I__8343\ : InMux
    port map (
            O => \N__39461\,
            I => \N__39458\
        );

    \I__8342\ : LocalMux
    port map (
            O => \N__39458\,
            I => \N__39455\
        );

    \I__8341\ : Odrv4
    port map (
            O => \N__39455\,
            I => \current_shift_inst.un4_control_input_1_axb_25\
        );

    \I__8340\ : InMux
    port map (
            O => \N__39452\,
            I => \bfn_16_18_0_\
        );

    \I__8339\ : InMux
    port map (
            O => \N__39449\,
            I => \current_shift_inst.un4_control_input_1_cry_25\
        );

    \I__8338\ : InMux
    port map (
            O => \N__39446\,
            I => \current_shift_inst.un4_control_input_1_cry_26\
        );

    \I__8337\ : InMux
    port map (
            O => \N__39443\,
            I => \N__39439\
        );

    \I__8336\ : CascadeMux
    port map (
            O => \N__39442\,
            I => \N__39436\
        );

    \I__8335\ : LocalMux
    port map (
            O => \N__39439\,
            I => \N__39432\
        );

    \I__8334\ : InMux
    port map (
            O => \N__39436\,
            I => \N__39427\
        );

    \I__8333\ : InMux
    port map (
            O => \N__39435\,
            I => \N__39427\
        );

    \I__8332\ : Odrv12
    port map (
            O => \N__39432\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__8331\ : LocalMux
    port map (
            O => \N__39427\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__8330\ : InMux
    port map (
            O => \N__39422\,
            I => \current_shift_inst.un4_control_input_1_cry_27\
        );

    \I__8329\ : InMux
    port map (
            O => \N__39419\,
            I => \current_shift_inst.un4_control_input_1_cry_28\
        );

    \I__8328\ : InMux
    port map (
            O => \N__39416\,
            I => \current_shift_inst.un4_control_input_1_cry_12\
        );

    \I__8327\ : InMux
    port map (
            O => \N__39413\,
            I => \N__39410\
        );

    \I__8326\ : LocalMux
    port map (
            O => \N__39410\,
            I => \N__39407\
        );

    \I__8325\ : Odrv4
    port map (
            O => \N__39407\,
            I => \current_shift_inst.un4_control_input_1_axb_14\
        );

    \I__8324\ : InMux
    port map (
            O => \N__39404\,
            I => \current_shift_inst.un4_control_input_1_cry_13\
        );

    \I__8323\ : InMux
    port map (
            O => \N__39401\,
            I => \N__39398\
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__39398\,
            I => \N__39395\
        );

    \I__8321\ : Span4Mux_h
    port map (
            O => \N__39395\,
            I => \N__39392\
        );

    \I__8320\ : Odrv4
    port map (
            O => \N__39392\,
            I => \current_shift_inst.un4_control_input_1_axb_15\
        );

    \I__8319\ : InMux
    port map (
            O => \N__39389\,
            I => \current_shift_inst.un4_control_input_1_cry_14\
        );

    \I__8318\ : InMux
    port map (
            O => \N__39386\,
            I => \N__39383\
        );

    \I__8317\ : LocalMux
    port map (
            O => \N__39383\,
            I => \N__39380\
        );

    \I__8316\ : Span4Mux_h
    port map (
            O => \N__39380\,
            I => \N__39377\
        );

    \I__8315\ : Odrv4
    port map (
            O => \N__39377\,
            I => \current_shift_inst.un4_control_input_1_axb_16\
        );

    \I__8314\ : InMux
    port map (
            O => \N__39374\,
            I => \current_shift_inst.un4_control_input_1_cry_15\
        );

    \I__8313\ : InMux
    port map (
            O => \N__39371\,
            I => \bfn_16_17_0_\
        );

    \I__8312\ : InMux
    port map (
            O => \N__39368\,
            I => \N__39365\
        );

    \I__8311\ : LocalMux
    port map (
            O => \N__39365\,
            I => \N__39362\
        );

    \I__8310\ : Odrv4
    port map (
            O => \N__39362\,
            I => \current_shift_inst.un4_control_input_1_axb_18\
        );

    \I__8309\ : InMux
    port map (
            O => \N__39359\,
            I => \current_shift_inst.un4_control_input_1_cry_17\
        );

    \I__8308\ : InMux
    port map (
            O => \N__39356\,
            I => \current_shift_inst.un4_control_input_1_cry_18\
        );

    \I__8307\ : InMux
    port map (
            O => \N__39353\,
            I => \current_shift_inst.un4_control_input_1_cry_19\
        );

    \I__8306\ : InMux
    port map (
            O => \N__39350\,
            I => \N__39347\
        );

    \I__8305\ : LocalMux
    port map (
            O => \N__39347\,
            I => \N__39344\
        );

    \I__8304\ : Span4Mux_v
    port map (
            O => \N__39344\,
            I => \N__39341\
        );

    \I__8303\ : Odrv4
    port map (
            O => \N__39341\,
            I => \current_shift_inst.un4_control_input_1_axb_21\
        );

    \I__8302\ : InMux
    port map (
            O => \N__39338\,
            I => \current_shift_inst.un4_control_input_1_cry_20\
        );

    \I__8301\ : InMux
    port map (
            O => \N__39335\,
            I => \N__39332\
        );

    \I__8300\ : LocalMux
    port map (
            O => \N__39332\,
            I => \current_shift_inst.un4_control_input_1_axb_4\
        );

    \I__8299\ : InMux
    port map (
            O => \N__39329\,
            I => \current_shift_inst.un4_control_input_1_cry_3\
        );

    \I__8298\ : InMux
    port map (
            O => \N__39326\,
            I => \N__39323\
        );

    \I__8297\ : LocalMux
    port map (
            O => \N__39323\,
            I => \current_shift_inst.un4_control_input_1_axb_5\
        );

    \I__8296\ : InMux
    port map (
            O => \N__39320\,
            I => \current_shift_inst.un4_control_input_1_cry_4\
        );

    \I__8295\ : InMux
    port map (
            O => \N__39317\,
            I => \N__39314\
        );

    \I__8294\ : LocalMux
    port map (
            O => \N__39314\,
            I => \current_shift_inst.un4_control_input_1_axb_6\
        );

    \I__8293\ : InMux
    port map (
            O => \N__39311\,
            I => \current_shift_inst.un4_control_input_1_cry_5\
        );

    \I__8292\ : InMux
    port map (
            O => \N__39308\,
            I => \N__39305\
        );

    \I__8291\ : LocalMux
    port map (
            O => \N__39305\,
            I => \current_shift_inst.un4_control_input_1_axb_7\
        );

    \I__8290\ : InMux
    port map (
            O => \N__39302\,
            I => \current_shift_inst.un4_control_input_1_cry_6\
        );

    \I__8289\ : InMux
    port map (
            O => \N__39299\,
            I => \N__39296\
        );

    \I__8288\ : LocalMux
    port map (
            O => \N__39296\,
            I => \current_shift_inst.un4_control_input_1_axb_8\
        );

    \I__8287\ : InMux
    port map (
            O => \N__39293\,
            I => \current_shift_inst.un4_control_input_1_cry_7\
        );

    \I__8286\ : InMux
    port map (
            O => \N__39290\,
            I => \bfn_16_16_0_\
        );

    \I__8285\ : InMux
    port map (
            O => \N__39287\,
            I => \N__39284\
        );

    \I__8284\ : LocalMux
    port map (
            O => \N__39284\,
            I => \N__39281\
        );

    \I__8283\ : Span4Mux_h
    port map (
            O => \N__39281\,
            I => \N__39278\
        );

    \I__8282\ : Odrv4
    port map (
            O => \N__39278\,
            I => \current_shift_inst.un4_control_input_1_axb_10\
        );

    \I__8281\ : InMux
    port map (
            O => \N__39275\,
            I => \current_shift_inst.un4_control_input_1_cry_9\
        );

    \I__8280\ : InMux
    port map (
            O => \N__39272\,
            I => \current_shift_inst.un4_control_input_1_cry_10\
        );

    \I__8279\ : InMux
    port map (
            O => \N__39269\,
            I => \N__39266\
        );

    \I__8278\ : LocalMux
    port map (
            O => \N__39266\,
            I => \current_shift_inst.un4_control_input_1_axb_12\
        );

    \I__8277\ : InMux
    port map (
            O => \N__39263\,
            I => \current_shift_inst.un4_control_input_1_cry_11\
        );

    \I__8276\ : InMux
    port map (
            O => \N__39260\,
            I => \N__39257\
        );

    \I__8275\ : LocalMux
    port map (
            O => \N__39257\,
            I => \N__39254\
        );

    \I__8274\ : Span4Mux_h
    port map (
            O => \N__39254\,
            I => \N__39251\
        );

    \I__8273\ : Span4Mux_v
    port map (
            O => \N__39251\,
            I => \N__39248\
        );

    \I__8272\ : Odrv4
    port map (
            O => \N__39248\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\
        );

    \I__8271\ : InMux
    port map (
            O => \N__39245\,
            I => \N__39242\
        );

    \I__8270\ : LocalMux
    port map (
            O => \N__39242\,
            I => \N__39239\
        );

    \I__8269\ : Span4Mux_h
    port map (
            O => \N__39239\,
            I => \N__39236\
        );

    \I__8268\ : Odrv4
    port map (
            O => \N__39236\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI68O61_6\
        );

    \I__8267\ : InMux
    port map (
            O => \N__39233\,
            I => \current_shift_inst.un4_control_input_1_cry_1\
        );

    \I__8266\ : InMux
    port map (
            O => \N__39230\,
            I => \N__39227\
        );

    \I__8265\ : LocalMux
    port map (
            O => \N__39227\,
            I => \current_shift_inst.un4_control_input_1_axb_3\
        );

    \I__8264\ : InMux
    port map (
            O => \N__39224\,
            I => \current_shift_inst.un4_control_input_1_cry_2\
        );

    \I__8263\ : InMux
    port map (
            O => \N__39221\,
            I => \N__39218\
        );

    \I__8262\ : LocalMux
    port map (
            O => \N__39218\,
            I => \N__39214\
        );

    \I__8261\ : InMux
    port map (
            O => \N__39217\,
            I => \N__39211\
        );

    \I__8260\ : Span4Mux_v
    port map (
            O => \N__39214\,
            I => \N__39208\
        );

    \I__8259\ : LocalMux
    port map (
            O => \N__39211\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__8258\ : Odrv4
    port map (
            O => \N__39208\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__8257\ : CascadeMux
    port map (
            O => \N__39203\,
            I => \N__39200\
        );

    \I__8256\ : InMux
    port map (
            O => \N__39200\,
            I => \N__39195\
        );

    \I__8255\ : InMux
    port map (
            O => \N__39199\,
            I => \N__39192\
        );

    \I__8254\ : InMux
    port map (
            O => \N__39198\,
            I => \N__39189\
        );

    \I__8253\ : LocalMux
    port map (
            O => \N__39195\,
            I => \N__39184\
        );

    \I__8252\ : LocalMux
    port map (
            O => \N__39192\,
            I => \N__39184\
        );

    \I__8251\ : LocalMux
    port map (
            O => \N__39189\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__8250\ : Odrv12
    port map (
            O => \N__39184\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__8249\ : InMux
    port map (
            O => \N__39179\,
            I => \N__39176\
        );

    \I__8248\ : LocalMux
    port map (
            O => \N__39176\,
            I => \N__39170\
        );

    \I__8247\ : InMux
    port map (
            O => \N__39175\,
            I => \N__39167\
        );

    \I__8246\ : InMux
    port map (
            O => \N__39174\,
            I => \N__39162\
        );

    \I__8245\ : InMux
    port map (
            O => \N__39173\,
            I => \N__39162\
        );

    \I__8244\ : Span4Mux_h
    port map (
            O => \N__39170\,
            I => \N__39159\
        );

    \I__8243\ : LocalMux
    port map (
            O => \N__39167\,
            I => \N__39156\
        );

    \I__8242\ : LocalMux
    port map (
            O => \N__39162\,
            I => \N__39153\
        );

    \I__8241\ : Span4Mux_v
    port map (
            O => \N__39159\,
            I => \N__39150\
        );

    \I__8240\ : Span4Mux_v
    port map (
            O => \N__39156\,
            I => \N__39147\
        );

    \I__8239\ : Span4Mux_h
    port map (
            O => \N__39153\,
            I => \N__39144\
        );

    \I__8238\ : Odrv4
    port map (
            O => \N__39150\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__8237\ : Odrv4
    port map (
            O => \N__39147\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__8236\ : Odrv4
    port map (
            O => \N__39144\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__8235\ : InMux
    port map (
            O => \N__39137\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__8234\ : InMux
    port map (
            O => \N__39134\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__8233\ : InMux
    port map (
            O => \N__39131\,
            I => \N__39128\
        );

    \I__8232\ : LocalMux
    port map (
            O => \N__39128\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt16\
        );

    \I__8231\ : CascadeMux
    port map (
            O => \N__39125\,
            I => \N__39121\
        );

    \I__8230\ : InMux
    port map (
            O => \N__39124\,
            I => \N__39116\
        );

    \I__8229\ : InMux
    port map (
            O => \N__39121\,
            I => \N__39116\
        );

    \I__8228\ : LocalMux
    port map (
            O => \N__39116\,
            I => \N__39112\
        );

    \I__8227\ : InMux
    port map (
            O => \N__39115\,
            I => \N__39109\
        );

    \I__8226\ : Span4Mux_h
    port map (
            O => \N__39112\,
            I => \N__39106\
        );

    \I__8225\ : LocalMux
    port map (
            O => \N__39109\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__8224\ : Odrv4
    port map (
            O => \N__39106\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__8223\ : CascadeMux
    port map (
            O => \N__39101\,
            I => \N__39096\
        );

    \I__8222\ : InMux
    port map (
            O => \N__39100\,
            I => \N__39093\
        );

    \I__8221\ : InMux
    port map (
            O => \N__39099\,
            I => \N__39088\
        );

    \I__8220\ : InMux
    port map (
            O => \N__39096\,
            I => \N__39088\
        );

    \I__8219\ : LocalMux
    port map (
            O => \N__39093\,
            I => \N__39083\
        );

    \I__8218\ : LocalMux
    port map (
            O => \N__39088\,
            I => \N__39083\
        );

    \I__8217\ : Odrv4
    port map (
            O => \N__39083\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__8216\ : CascadeMux
    port map (
            O => \N__39080\,
            I => \N__39077\
        );

    \I__8215\ : InMux
    port map (
            O => \N__39077\,
            I => \N__39074\
        );

    \I__8214\ : LocalMux
    port map (
            O => \N__39074\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\
        );

    \I__8213\ : InMux
    port map (
            O => \N__39071\,
            I => \N__39065\
        );

    \I__8212\ : InMux
    port map (
            O => \N__39070\,
            I => \N__39065\
        );

    \I__8211\ : LocalMux
    port map (
            O => \N__39065\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\
        );

    \I__8210\ : InMux
    port map (
            O => \N__39062\,
            I => \N__39059\
        );

    \I__8209\ : LocalMux
    port map (
            O => \N__39059\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\
        );

    \I__8208\ : InMux
    port map (
            O => \N__39056\,
            I => \N__39053\
        );

    \I__8207\ : LocalMux
    port map (
            O => \N__39053\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\
        );

    \I__8206\ : InMux
    port map (
            O => \N__39050\,
            I => \N__39043\
        );

    \I__8205\ : InMux
    port map (
            O => \N__39049\,
            I => \N__39043\
        );

    \I__8204\ : InMux
    port map (
            O => \N__39048\,
            I => \N__39040\
        );

    \I__8203\ : LocalMux
    port map (
            O => \N__39043\,
            I => \N__39037\
        );

    \I__8202\ : LocalMux
    port map (
            O => \N__39040\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__8201\ : Odrv12
    port map (
            O => \N__39037\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__8200\ : InMux
    port map (
            O => \N__39032\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__8199\ : CascadeMux
    port map (
            O => \N__39029\,
            I => \N__39026\
        );

    \I__8198\ : InMux
    port map (
            O => \N__39026\,
            I => \N__39021\
        );

    \I__8197\ : InMux
    port map (
            O => \N__39025\,
            I => \N__39018\
        );

    \I__8196\ : InMux
    port map (
            O => \N__39024\,
            I => \N__39015\
        );

    \I__8195\ : LocalMux
    port map (
            O => \N__39021\,
            I => \N__39010\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__39018\,
            I => \N__39010\
        );

    \I__8193\ : LocalMux
    port map (
            O => \N__39015\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__8192\ : Odrv12
    port map (
            O => \N__39010\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__8191\ : InMux
    port map (
            O => \N__39005\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__8190\ : CascadeMux
    port map (
            O => \N__39002\,
            I => \N__38998\
        );

    \I__8189\ : InMux
    port map (
            O => \N__39001\,
            I => \N__38995\
        );

    \I__8188\ : InMux
    port map (
            O => \N__38998\,
            I => \N__38992\
        );

    \I__8187\ : LocalMux
    port map (
            O => \N__38995\,
            I => \N__38988\
        );

    \I__8186\ : LocalMux
    port map (
            O => \N__38992\,
            I => \N__38985\
        );

    \I__8185\ : InMux
    port map (
            O => \N__38991\,
            I => \N__38982\
        );

    \I__8184\ : Span4Mux_v
    port map (
            O => \N__38988\,
            I => \N__38977\
        );

    \I__8183\ : Span4Mux_v
    port map (
            O => \N__38985\,
            I => \N__38977\
        );

    \I__8182\ : LocalMux
    port map (
            O => \N__38982\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__8181\ : Odrv4
    port map (
            O => \N__38977\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__8180\ : InMux
    port map (
            O => \N__38972\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__8179\ : InMux
    port map (
            O => \N__38969\,
            I => \N__38963\
        );

    \I__8178\ : InMux
    port map (
            O => \N__38968\,
            I => \N__38963\
        );

    \I__8177\ : LocalMux
    port map (
            O => \N__38963\,
            I => \N__38959\
        );

    \I__8176\ : InMux
    port map (
            O => \N__38962\,
            I => \N__38956\
        );

    \I__8175\ : Span4Mux_v
    port map (
            O => \N__38959\,
            I => \N__38953\
        );

    \I__8174\ : LocalMux
    port map (
            O => \N__38956\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__8173\ : Odrv4
    port map (
            O => \N__38953\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__8172\ : InMux
    port map (
            O => \N__38948\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__8171\ : CascadeMux
    port map (
            O => \N__38945\,
            I => \N__38941\
        );

    \I__8170\ : CascadeMux
    port map (
            O => \N__38944\,
            I => \N__38938\
        );

    \I__8169\ : InMux
    port map (
            O => \N__38941\,
            I => \N__38933\
        );

    \I__8168\ : InMux
    port map (
            O => \N__38938\,
            I => \N__38933\
        );

    \I__8167\ : LocalMux
    port map (
            O => \N__38933\,
            I => \N__38929\
        );

    \I__8166\ : InMux
    port map (
            O => \N__38932\,
            I => \N__38926\
        );

    \I__8165\ : Span4Mux_v
    port map (
            O => \N__38929\,
            I => \N__38923\
        );

    \I__8164\ : LocalMux
    port map (
            O => \N__38926\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__8163\ : Odrv4
    port map (
            O => \N__38923\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__8162\ : InMux
    port map (
            O => \N__38918\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__8161\ : CascadeMux
    port map (
            O => \N__38915\,
            I => \N__38911\
        );

    \I__8160\ : CascadeMux
    port map (
            O => \N__38914\,
            I => \N__38908\
        );

    \I__8159\ : InMux
    port map (
            O => \N__38911\,
            I => \N__38905\
        );

    \I__8158\ : InMux
    port map (
            O => \N__38908\,
            I => \N__38902\
        );

    \I__8157\ : LocalMux
    port map (
            O => \N__38905\,
            I => \N__38896\
        );

    \I__8156\ : LocalMux
    port map (
            O => \N__38902\,
            I => \N__38896\
        );

    \I__8155\ : InMux
    port map (
            O => \N__38901\,
            I => \N__38893\
        );

    \I__8154\ : Span4Mux_v
    port map (
            O => \N__38896\,
            I => \N__38890\
        );

    \I__8153\ : LocalMux
    port map (
            O => \N__38893\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__8152\ : Odrv4
    port map (
            O => \N__38890\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__8151\ : InMux
    port map (
            O => \N__38885\,
            I => \bfn_16_12_0_\
        );

    \I__8150\ : CascadeMux
    port map (
            O => \N__38882\,
            I => \N__38879\
        );

    \I__8149\ : InMux
    port map (
            O => \N__38879\,
            I => \N__38874\
        );

    \I__8148\ : InMux
    port map (
            O => \N__38878\,
            I => \N__38871\
        );

    \I__8147\ : InMux
    port map (
            O => \N__38877\,
            I => \N__38868\
        );

    \I__8146\ : LocalMux
    port map (
            O => \N__38874\,
            I => \N__38863\
        );

    \I__8145\ : LocalMux
    port map (
            O => \N__38871\,
            I => \N__38863\
        );

    \I__8144\ : LocalMux
    port map (
            O => \N__38868\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__8143\ : Odrv12
    port map (
            O => \N__38863\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__8142\ : InMux
    port map (
            O => \N__38858\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__8141\ : InMux
    port map (
            O => \N__38855\,
            I => \N__38848\
        );

    \I__8140\ : InMux
    port map (
            O => \N__38854\,
            I => \N__38848\
        );

    \I__8139\ : InMux
    port map (
            O => \N__38853\,
            I => \N__38845\
        );

    \I__8138\ : LocalMux
    port map (
            O => \N__38848\,
            I => \N__38842\
        );

    \I__8137\ : LocalMux
    port map (
            O => \N__38845\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__8136\ : Odrv12
    port map (
            O => \N__38842\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__8135\ : CascadeMux
    port map (
            O => \N__38837\,
            I => \N__38834\
        );

    \I__8134\ : InMux
    port map (
            O => \N__38834\,
            I => \N__38830\
        );

    \I__8133\ : InMux
    port map (
            O => \N__38833\,
            I => \N__38827\
        );

    \I__8132\ : LocalMux
    port map (
            O => \N__38830\,
            I => \N__38824\
        );

    \I__8131\ : LocalMux
    port map (
            O => \N__38827\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__8130\ : Odrv12
    port map (
            O => \N__38824\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__8129\ : InMux
    port map (
            O => \N__38819\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__8128\ : InMux
    port map (
            O => \N__38816\,
            I => \N__38811\
        );

    \I__8127\ : InMux
    port map (
            O => \N__38815\,
            I => \N__38808\
        );

    \I__8126\ : InMux
    port map (
            O => \N__38814\,
            I => \N__38805\
        );

    \I__8125\ : LocalMux
    port map (
            O => \N__38811\,
            I => \N__38802\
        );

    \I__8124\ : LocalMux
    port map (
            O => \N__38808\,
            I => \N__38797\
        );

    \I__8123\ : LocalMux
    port map (
            O => \N__38805\,
            I => \N__38797\
        );

    \I__8122\ : Span4Mux_v
    port map (
            O => \N__38802\,
            I => \N__38791\
        );

    \I__8121\ : Span4Mux_v
    port map (
            O => \N__38797\,
            I => \N__38791\
        );

    \I__8120\ : InMux
    port map (
            O => \N__38796\,
            I => \N__38788\
        );

    \I__8119\ : Odrv4
    port map (
            O => \N__38791\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__8118\ : LocalMux
    port map (
            O => \N__38788\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__8117\ : InMux
    port map (
            O => \N__38783\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__8116\ : InMux
    port map (
            O => \N__38780\,
            I => \N__38774\
        );

    \I__8115\ : InMux
    port map (
            O => \N__38779\,
            I => \N__38774\
        );

    \I__8114\ : LocalMux
    port map (
            O => \N__38774\,
            I => \N__38770\
        );

    \I__8113\ : InMux
    port map (
            O => \N__38773\,
            I => \N__38767\
        );

    \I__8112\ : Span4Mux_v
    port map (
            O => \N__38770\,
            I => \N__38764\
        );

    \I__8111\ : LocalMux
    port map (
            O => \N__38767\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__8110\ : Odrv4
    port map (
            O => \N__38764\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__8109\ : InMux
    port map (
            O => \N__38759\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__8108\ : CascadeMux
    port map (
            O => \N__38756\,
            I => \N__38752\
        );

    \I__8107\ : CascadeMux
    port map (
            O => \N__38755\,
            I => \N__38749\
        );

    \I__8106\ : InMux
    port map (
            O => \N__38752\,
            I => \N__38743\
        );

    \I__8105\ : InMux
    port map (
            O => \N__38749\,
            I => \N__38743\
        );

    \I__8104\ : InMux
    port map (
            O => \N__38748\,
            I => \N__38740\
        );

    \I__8103\ : LocalMux
    port map (
            O => \N__38743\,
            I => \N__38737\
        );

    \I__8102\ : LocalMux
    port map (
            O => \N__38740\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__8101\ : Odrv12
    port map (
            O => \N__38737\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__8100\ : InMux
    port map (
            O => \N__38732\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__8099\ : CascadeMux
    port map (
            O => \N__38729\,
            I => \N__38725\
        );

    \I__8098\ : CascadeMux
    port map (
            O => \N__38728\,
            I => \N__38722\
        );

    \I__8097\ : InMux
    port map (
            O => \N__38725\,
            I => \N__38716\
        );

    \I__8096\ : InMux
    port map (
            O => \N__38722\,
            I => \N__38716\
        );

    \I__8095\ : InMux
    port map (
            O => \N__38721\,
            I => \N__38713\
        );

    \I__8094\ : LocalMux
    port map (
            O => \N__38716\,
            I => \N__38710\
        );

    \I__8093\ : LocalMux
    port map (
            O => \N__38713\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__8092\ : Odrv12
    port map (
            O => \N__38710\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__8091\ : InMux
    port map (
            O => \N__38705\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__8090\ : InMux
    port map (
            O => \N__38702\,
            I => \N__38696\
        );

    \I__8089\ : InMux
    port map (
            O => \N__38701\,
            I => \N__38696\
        );

    \I__8088\ : LocalMux
    port map (
            O => \N__38696\,
            I => \N__38692\
        );

    \I__8087\ : InMux
    port map (
            O => \N__38695\,
            I => \N__38689\
        );

    \I__8086\ : Span4Mux_v
    port map (
            O => \N__38692\,
            I => \N__38686\
        );

    \I__8085\ : LocalMux
    port map (
            O => \N__38689\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__8084\ : Odrv4
    port map (
            O => \N__38686\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__8083\ : InMux
    port map (
            O => \N__38681\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__8082\ : CascadeMux
    port map (
            O => \N__38678\,
            I => \N__38675\
        );

    \I__8081\ : InMux
    port map (
            O => \N__38675\,
            I => \N__38670\
        );

    \I__8080\ : InMux
    port map (
            O => \N__38674\,
            I => \N__38667\
        );

    \I__8079\ : InMux
    port map (
            O => \N__38673\,
            I => \N__38664\
        );

    \I__8078\ : LocalMux
    port map (
            O => \N__38670\,
            I => \N__38659\
        );

    \I__8077\ : LocalMux
    port map (
            O => \N__38667\,
            I => \N__38659\
        );

    \I__8076\ : LocalMux
    port map (
            O => \N__38664\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__8075\ : Odrv12
    port map (
            O => \N__38659\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__8074\ : InMux
    port map (
            O => \N__38654\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__8073\ : CascadeMux
    port map (
            O => \N__38651\,
            I => \N__38647\
        );

    \I__8072\ : InMux
    port map (
            O => \N__38650\,
            I => \N__38644\
        );

    \I__8071\ : InMux
    port map (
            O => \N__38647\,
            I => \N__38641\
        );

    \I__8070\ : LocalMux
    port map (
            O => \N__38644\,
            I => \N__38635\
        );

    \I__8069\ : LocalMux
    port map (
            O => \N__38641\,
            I => \N__38635\
        );

    \I__8068\ : InMux
    port map (
            O => \N__38640\,
            I => \N__38632\
        );

    \I__8067\ : Span4Mux_v
    port map (
            O => \N__38635\,
            I => \N__38629\
        );

    \I__8066\ : LocalMux
    port map (
            O => \N__38632\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__8065\ : Odrv4
    port map (
            O => \N__38629\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__8064\ : InMux
    port map (
            O => \N__38624\,
            I => \bfn_16_11_0_\
        );

    \I__8063\ : CascadeMux
    port map (
            O => \N__38621\,
            I => \N__38618\
        );

    \I__8062\ : InMux
    port map (
            O => \N__38618\,
            I => \N__38613\
        );

    \I__8061\ : InMux
    port map (
            O => \N__38617\,
            I => \N__38610\
        );

    \I__8060\ : InMux
    port map (
            O => \N__38616\,
            I => \N__38607\
        );

    \I__8059\ : LocalMux
    port map (
            O => \N__38613\,
            I => \N__38602\
        );

    \I__8058\ : LocalMux
    port map (
            O => \N__38610\,
            I => \N__38602\
        );

    \I__8057\ : LocalMux
    port map (
            O => \N__38607\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__8056\ : Odrv12
    port map (
            O => \N__38602\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__8055\ : InMux
    port map (
            O => \N__38597\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__8054\ : CascadeMux
    port map (
            O => \N__38594\,
            I => \N__38590\
        );

    \I__8053\ : CascadeMux
    port map (
            O => \N__38593\,
            I => \N__38587\
        );

    \I__8052\ : InMux
    port map (
            O => \N__38590\,
            I => \N__38581\
        );

    \I__8051\ : InMux
    port map (
            O => \N__38587\,
            I => \N__38581\
        );

    \I__8050\ : InMux
    port map (
            O => \N__38586\,
            I => \N__38578\
        );

    \I__8049\ : LocalMux
    port map (
            O => \N__38581\,
            I => \N__38575\
        );

    \I__8048\ : LocalMux
    port map (
            O => \N__38578\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__8047\ : Odrv12
    port map (
            O => \N__38575\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__8046\ : InMux
    port map (
            O => \N__38570\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__8045\ : InMux
    port map (
            O => \N__38567\,
            I => \N__38563\
        );

    \I__8044\ : CascadeMux
    port map (
            O => \N__38566\,
            I => \N__38560\
        );

    \I__8043\ : LocalMux
    port map (
            O => \N__38563\,
            I => \N__38556\
        );

    \I__8042\ : InMux
    port map (
            O => \N__38560\,
            I => \N__38553\
        );

    \I__8041\ : InMux
    port map (
            O => \N__38559\,
            I => \N__38550\
        );

    \I__8040\ : Sp12to4
    port map (
            O => \N__38556\,
            I => \N__38545\
        );

    \I__8039\ : LocalMux
    port map (
            O => \N__38553\,
            I => \N__38545\
        );

    \I__8038\ : LocalMux
    port map (
            O => \N__38550\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__8037\ : Odrv12
    port map (
            O => \N__38545\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__8036\ : InMux
    port map (
            O => \N__38540\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__8035\ : InMux
    port map (
            O => \N__38537\,
            I => \N__38531\
        );

    \I__8034\ : InMux
    port map (
            O => \N__38536\,
            I => \N__38531\
        );

    \I__8033\ : LocalMux
    port map (
            O => \N__38531\,
            I => \N__38527\
        );

    \I__8032\ : InMux
    port map (
            O => \N__38530\,
            I => \N__38524\
        );

    \I__8031\ : Span4Mux_v
    port map (
            O => \N__38527\,
            I => \N__38521\
        );

    \I__8030\ : LocalMux
    port map (
            O => \N__38524\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__8029\ : Odrv4
    port map (
            O => \N__38521\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__8028\ : InMux
    port map (
            O => \N__38516\,
            I => \N__38513\
        );

    \I__8027\ : LocalMux
    port map (
            O => \N__38513\,
            I => \N__38509\
        );

    \I__8026\ : InMux
    port map (
            O => \N__38512\,
            I => \N__38506\
        );

    \I__8025\ : Span4Mux_v
    port map (
            O => \N__38509\,
            I => \N__38501\
        );

    \I__8024\ : LocalMux
    port map (
            O => \N__38506\,
            I => \N__38498\
        );

    \I__8023\ : InMux
    port map (
            O => \N__38505\,
            I => \N__38495\
        );

    \I__8022\ : InMux
    port map (
            O => \N__38504\,
            I => \N__38492\
        );

    \I__8021\ : Odrv4
    port map (
            O => \N__38501\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__8020\ : Odrv4
    port map (
            O => \N__38498\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__8019\ : LocalMux
    port map (
            O => \N__38495\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__8018\ : LocalMux
    port map (
            O => \N__38492\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__8017\ : InMux
    port map (
            O => \N__38483\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__8016\ : CascadeMux
    port map (
            O => \N__38480\,
            I => \N__38476\
        );

    \I__8015\ : CascadeMux
    port map (
            O => \N__38479\,
            I => \N__38473\
        );

    \I__8014\ : InMux
    port map (
            O => \N__38476\,
            I => \N__38467\
        );

    \I__8013\ : InMux
    port map (
            O => \N__38473\,
            I => \N__38467\
        );

    \I__8012\ : InMux
    port map (
            O => \N__38472\,
            I => \N__38464\
        );

    \I__8011\ : LocalMux
    port map (
            O => \N__38467\,
            I => \N__38461\
        );

    \I__8010\ : LocalMux
    port map (
            O => \N__38464\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__8009\ : Odrv12
    port map (
            O => \N__38461\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__8008\ : InMux
    port map (
            O => \N__38456\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__8007\ : CascadeMux
    port map (
            O => \N__38453\,
            I => \N__38449\
        );

    \I__8006\ : CascadeMux
    port map (
            O => \N__38452\,
            I => \N__38446\
        );

    \I__8005\ : InMux
    port map (
            O => \N__38449\,
            I => \N__38440\
        );

    \I__8004\ : InMux
    port map (
            O => \N__38446\,
            I => \N__38440\
        );

    \I__8003\ : InMux
    port map (
            O => \N__38445\,
            I => \N__38437\
        );

    \I__8002\ : LocalMux
    port map (
            O => \N__38440\,
            I => \N__38434\
        );

    \I__8001\ : LocalMux
    port map (
            O => \N__38437\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__8000\ : Odrv12
    port map (
            O => \N__38434\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__7999\ : InMux
    port map (
            O => \N__38429\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__7998\ : InMux
    port map (
            O => \N__38426\,
            I => \N__38420\
        );

    \I__7997\ : InMux
    port map (
            O => \N__38425\,
            I => \N__38420\
        );

    \I__7996\ : LocalMux
    port map (
            O => \N__38420\,
            I => \N__38416\
        );

    \I__7995\ : InMux
    port map (
            O => \N__38419\,
            I => \N__38413\
        );

    \I__7994\ : Span4Mux_v
    port map (
            O => \N__38416\,
            I => \N__38410\
        );

    \I__7993\ : LocalMux
    port map (
            O => \N__38413\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__7992\ : Odrv4
    port map (
            O => \N__38410\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__7991\ : InMux
    port map (
            O => \N__38405\,
            I => \N__38401\
        );

    \I__7990\ : InMux
    port map (
            O => \N__38404\,
            I => \N__38396\
        );

    \I__7989\ : LocalMux
    port map (
            O => \N__38401\,
            I => \N__38393\
        );

    \I__7988\ : CascadeMux
    port map (
            O => \N__38400\,
            I => \N__38390\
        );

    \I__7987\ : InMux
    port map (
            O => \N__38399\,
            I => \N__38387\
        );

    \I__7986\ : LocalMux
    port map (
            O => \N__38396\,
            I => \N__38384\
        );

    \I__7985\ : Span4Mux_v
    port map (
            O => \N__38393\,
            I => \N__38381\
        );

    \I__7984\ : InMux
    port map (
            O => \N__38390\,
            I => \N__38378\
        );

    \I__7983\ : LocalMux
    port map (
            O => \N__38387\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__7982\ : Odrv4
    port map (
            O => \N__38384\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__7981\ : Odrv4
    port map (
            O => \N__38381\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__7980\ : LocalMux
    port map (
            O => \N__38378\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__7979\ : InMux
    port map (
            O => \N__38369\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__7978\ : InMux
    port map (
            O => \N__38366\,
            I => \N__38360\
        );

    \I__7977\ : InMux
    port map (
            O => \N__38365\,
            I => \N__38360\
        );

    \I__7976\ : LocalMux
    port map (
            O => \N__38360\,
            I => \N__38356\
        );

    \I__7975\ : InMux
    port map (
            O => \N__38359\,
            I => \N__38353\
        );

    \I__7974\ : Span4Mux_v
    port map (
            O => \N__38356\,
            I => \N__38350\
        );

    \I__7973\ : LocalMux
    port map (
            O => \N__38353\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__7972\ : Odrv4
    port map (
            O => \N__38350\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__7971\ : InMux
    port map (
            O => \N__38345\,
            I => \N__38342\
        );

    \I__7970\ : LocalMux
    port map (
            O => \N__38342\,
            I => \N__38339\
        );

    \I__7969\ : Span4Mux_h
    port map (
            O => \N__38339\,
            I => \N__38333\
        );

    \I__7968\ : InMux
    port map (
            O => \N__38338\,
            I => \N__38328\
        );

    \I__7967\ : InMux
    port map (
            O => \N__38337\,
            I => \N__38328\
        );

    \I__7966\ : InMux
    port map (
            O => \N__38336\,
            I => \N__38325\
        );

    \I__7965\ : Odrv4
    port map (
            O => \N__38333\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__7964\ : LocalMux
    port map (
            O => \N__38328\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__7963\ : LocalMux
    port map (
            O => \N__38325\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__7962\ : InMux
    port map (
            O => \N__38318\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__7961\ : CascadeMux
    port map (
            O => \N__38315\,
            I => \N__38311\
        );

    \I__7960\ : CascadeMux
    port map (
            O => \N__38314\,
            I => \N__38308\
        );

    \I__7959\ : InMux
    port map (
            O => \N__38311\,
            I => \N__38305\
        );

    \I__7958\ : InMux
    port map (
            O => \N__38308\,
            I => \N__38302\
        );

    \I__7957\ : LocalMux
    port map (
            O => \N__38305\,
            I => \N__38296\
        );

    \I__7956\ : LocalMux
    port map (
            O => \N__38302\,
            I => \N__38296\
        );

    \I__7955\ : InMux
    port map (
            O => \N__38301\,
            I => \N__38293\
        );

    \I__7954\ : Span4Mux_v
    port map (
            O => \N__38296\,
            I => \N__38290\
        );

    \I__7953\ : LocalMux
    port map (
            O => \N__38293\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__7952\ : Odrv4
    port map (
            O => \N__38290\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__7951\ : InMux
    port map (
            O => \N__38285\,
            I => \N__38281\
        );

    \I__7950\ : InMux
    port map (
            O => \N__38284\,
            I => \N__38278\
        );

    \I__7949\ : LocalMux
    port map (
            O => \N__38281\,
            I => \N__38275\
        );

    \I__7948\ : LocalMux
    port map (
            O => \N__38278\,
            I => \N__38270\
        );

    \I__7947\ : Span4Mux_h
    port map (
            O => \N__38275\,
            I => \N__38267\
        );

    \I__7946\ : InMux
    port map (
            O => \N__38274\,
            I => \N__38262\
        );

    \I__7945\ : InMux
    port map (
            O => \N__38273\,
            I => \N__38262\
        );

    \I__7944\ : Odrv4
    port map (
            O => \N__38270\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__7943\ : Odrv4
    port map (
            O => \N__38267\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__7942\ : LocalMux
    port map (
            O => \N__38262\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__7941\ : InMux
    port map (
            O => \N__38255\,
            I => \bfn_16_10_0_\
        );

    \I__7940\ : CascadeMux
    port map (
            O => \N__38252\,
            I => \N__38248\
        );

    \I__7939\ : CascadeMux
    port map (
            O => \N__38251\,
            I => \N__38245\
        );

    \I__7938\ : InMux
    port map (
            O => \N__38248\,
            I => \N__38242\
        );

    \I__7937\ : InMux
    port map (
            O => \N__38245\,
            I => \N__38239\
        );

    \I__7936\ : LocalMux
    port map (
            O => \N__38242\,
            I => \N__38233\
        );

    \I__7935\ : LocalMux
    port map (
            O => \N__38239\,
            I => \N__38233\
        );

    \I__7934\ : InMux
    port map (
            O => \N__38238\,
            I => \N__38230\
        );

    \I__7933\ : Span4Mux_v
    port map (
            O => \N__38233\,
            I => \N__38227\
        );

    \I__7932\ : LocalMux
    port map (
            O => \N__38230\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__7931\ : Odrv4
    port map (
            O => \N__38227\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__7930\ : InMux
    port map (
            O => \N__38222\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__7929\ : InMux
    port map (
            O => \N__38219\,
            I => \N__38213\
        );

    \I__7928\ : InMux
    port map (
            O => \N__38218\,
            I => \N__38213\
        );

    \I__7927\ : LocalMux
    port map (
            O => \N__38213\,
            I => \N__38209\
        );

    \I__7926\ : InMux
    port map (
            O => \N__38212\,
            I => \N__38206\
        );

    \I__7925\ : Span4Mux_v
    port map (
            O => \N__38209\,
            I => \N__38203\
        );

    \I__7924\ : LocalMux
    port map (
            O => \N__38206\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__7923\ : Odrv4
    port map (
            O => \N__38203\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__7922\ : InMux
    port map (
            O => \N__38198\,
            I => \bfn_16_8_0_\
        );

    \I__7921\ : InMux
    port map (
            O => \N__38195\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_24\
        );

    \I__7920\ : InMux
    port map (
            O => \N__38192\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_25\
        );

    \I__7919\ : InMux
    port map (
            O => \N__38189\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_26\
        );

    \I__7918\ : InMux
    port map (
            O => \N__38186\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_27\
        );

    \I__7917\ : InMux
    port map (
            O => \N__38183\,
            I => \N__38149\
        );

    \I__7916\ : InMux
    port map (
            O => \N__38182\,
            I => \N__38149\
        );

    \I__7915\ : InMux
    port map (
            O => \N__38181\,
            I => \N__38140\
        );

    \I__7914\ : InMux
    port map (
            O => \N__38180\,
            I => \N__38140\
        );

    \I__7913\ : InMux
    port map (
            O => \N__38179\,
            I => \N__38140\
        );

    \I__7912\ : InMux
    port map (
            O => \N__38178\,
            I => \N__38140\
        );

    \I__7911\ : InMux
    port map (
            O => \N__38177\,
            I => \N__38131\
        );

    \I__7910\ : InMux
    port map (
            O => \N__38176\,
            I => \N__38131\
        );

    \I__7909\ : InMux
    port map (
            O => \N__38175\,
            I => \N__38131\
        );

    \I__7908\ : InMux
    port map (
            O => \N__38174\,
            I => \N__38131\
        );

    \I__7907\ : InMux
    port map (
            O => \N__38173\,
            I => \N__38122\
        );

    \I__7906\ : InMux
    port map (
            O => \N__38172\,
            I => \N__38122\
        );

    \I__7905\ : InMux
    port map (
            O => \N__38171\,
            I => \N__38122\
        );

    \I__7904\ : InMux
    port map (
            O => \N__38170\,
            I => \N__38122\
        );

    \I__7903\ : InMux
    port map (
            O => \N__38169\,
            I => \N__38113\
        );

    \I__7902\ : InMux
    port map (
            O => \N__38168\,
            I => \N__38113\
        );

    \I__7901\ : InMux
    port map (
            O => \N__38167\,
            I => \N__38113\
        );

    \I__7900\ : InMux
    port map (
            O => \N__38166\,
            I => \N__38113\
        );

    \I__7899\ : InMux
    port map (
            O => \N__38165\,
            I => \N__38104\
        );

    \I__7898\ : InMux
    port map (
            O => \N__38164\,
            I => \N__38104\
        );

    \I__7897\ : InMux
    port map (
            O => \N__38163\,
            I => \N__38104\
        );

    \I__7896\ : InMux
    port map (
            O => \N__38162\,
            I => \N__38104\
        );

    \I__7895\ : InMux
    port map (
            O => \N__38161\,
            I => \N__38095\
        );

    \I__7894\ : InMux
    port map (
            O => \N__38160\,
            I => \N__38095\
        );

    \I__7893\ : InMux
    port map (
            O => \N__38159\,
            I => \N__38095\
        );

    \I__7892\ : InMux
    port map (
            O => \N__38158\,
            I => \N__38095\
        );

    \I__7891\ : InMux
    port map (
            O => \N__38157\,
            I => \N__38086\
        );

    \I__7890\ : InMux
    port map (
            O => \N__38156\,
            I => \N__38086\
        );

    \I__7889\ : InMux
    port map (
            O => \N__38155\,
            I => \N__38086\
        );

    \I__7888\ : InMux
    port map (
            O => \N__38154\,
            I => \N__38086\
        );

    \I__7887\ : LocalMux
    port map (
            O => \N__38149\,
            I => \N__38081\
        );

    \I__7886\ : LocalMux
    port map (
            O => \N__38140\,
            I => \N__38081\
        );

    \I__7885\ : LocalMux
    port map (
            O => \N__38131\,
            I => \N__38068\
        );

    \I__7884\ : LocalMux
    port map (
            O => \N__38122\,
            I => \N__38068\
        );

    \I__7883\ : LocalMux
    port map (
            O => \N__38113\,
            I => \N__38068\
        );

    \I__7882\ : LocalMux
    port map (
            O => \N__38104\,
            I => \N__38068\
        );

    \I__7881\ : LocalMux
    port map (
            O => \N__38095\,
            I => \N__38068\
        );

    \I__7880\ : LocalMux
    port map (
            O => \N__38086\,
            I => \N__38068\
        );

    \I__7879\ : Span4Mux_v
    port map (
            O => \N__38081\,
            I => \N__38063\
        );

    \I__7878\ : Span4Mux_v
    port map (
            O => \N__38068\,
            I => \N__38063\
        );

    \I__7877\ : Odrv4
    port map (
            O => \N__38063\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__7876\ : InMux
    port map (
            O => \N__38060\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_28\
        );

    \I__7875\ : CEMux
    port map (
            O => \N__38057\,
            I => \N__38051\
        );

    \I__7874\ : CEMux
    port map (
            O => \N__38056\,
            I => \N__38048\
        );

    \I__7873\ : CEMux
    port map (
            O => \N__38055\,
            I => \N__38045\
        );

    \I__7872\ : CEMux
    port map (
            O => \N__38054\,
            I => \N__38042\
        );

    \I__7871\ : LocalMux
    port map (
            O => \N__38051\,
            I => \N__38039\
        );

    \I__7870\ : LocalMux
    port map (
            O => \N__38048\,
            I => \N__38036\
        );

    \I__7869\ : LocalMux
    port map (
            O => \N__38045\,
            I => \N__38033\
        );

    \I__7868\ : LocalMux
    port map (
            O => \N__38042\,
            I => \N__38030\
        );

    \I__7867\ : Span4Mux_h
    port map (
            O => \N__38039\,
            I => \N__38027\
        );

    \I__7866\ : Span4Mux_h
    port map (
            O => \N__38036\,
            I => \N__38024\
        );

    \I__7865\ : Span4Mux_h
    port map (
            O => \N__38033\,
            I => \N__38021\
        );

    \I__7864\ : Span4Mux_v
    port map (
            O => \N__38030\,
            I => \N__38018\
        );

    \I__7863\ : Odrv4
    port map (
            O => \N__38027\,
            I => \delay_measurement_inst.delay_hc_timer.N_199_i\
        );

    \I__7862\ : Odrv4
    port map (
            O => \N__38024\,
            I => \delay_measurement_inst.delay_hc_timer.N_199_i\
        );

    \I__7861\ : Odrv4
    port map (
            O => \N__38021\,
            I => \delay_measurement_inst.delay_hc_timer.N_199_i\
        );

    \I__7860\ : Odrv4
    port map (
            O => \N__38018\,
            I => \delay_measurement_inst.delay_hc_timer.N_199_i\
        );

    \I__7859\ : InMux
    port map (
            O => \N__38009\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__7858\ : InMux
    port map (
            O => \N__38006\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_13\
        );

    \I__7857\ : InMux
    port map (
            O => \N__38003\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_14\
        );

    \I__7856\ : InMux
    port map (
            O => \N__38000\,
            I => \bfn_16_7_0_\
        );

    \I__7855\ : InMux
    port map (
            O => \N__37997\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_16\
        );

    \I__7854\ : InMux
    port map (
            O => \N__37994\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_17\
        );

    \I__7853\ : InMux
    port map (
            O => \N__37991\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_18\
        );

    \I__7852\ : InMux
    port map (
            O => \N__37988\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_19\
        );

    \I__7851\ : InMux
    port map (
            O => \N__37985\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_20\
        );

    \I__7850\ : InMux
    port map (
            O => \N__37982\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_21\
        );

    \I__7849\ : InMux
    port map (
            O => \N__37979\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_22\
        );

    \I__7848\ : InMux
    port map (
            O => \N__37976\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_4\
        );

    \I__7847\ : InMux
    port map (
            O => \N__37973\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_5\
        );

    \I__7846\ : InMux
    port map (
            O => \N__37970\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_6\
        );

    \I__7845\ : InMux
    port map (
            O => \N__37967\,
            I => \bfn_16_6_0_\
        );

    \I__7844\ : InMux
    port map (
            O => \N__37964\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_8\
        );

    \I__7843\ : InMux
    port map (
            O => \N__37961\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_9\
        );

    \I__7842\ : InMux
    port map (
            O => \N__37958\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_10\
        );

    \I__7841\ : InMux
    port map (
            O => \N__37955\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_11\
        );

    \I__7840\ : InMux
    port map (
            O => \N__37952\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_12\
        );

    \I__7839\ : InMux
    port map (
            O => \N__37949\,
            I => \N__37944\
        );

    \I__7838\ : InMux
    port map (
            O => \N__37948\,
            I => \N__37940\
        );

    \I__7837\ : InMux
    port map (
            O => \N__37947\,
            I => \N__37937\
        );

    \I__7836\ : LocalMux
    port map (
            O => \N__37944\,
            I => \N__37934\
        );

    \I__7835\ : InMux
    port map (
            O => \N__37943\,
            I => \N__37931\
        );

    \I__7834\ : LocalMux
    port map (
            O => \N__37940\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__7833\ : LocalMux
    port map (
            O => \N__37937\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__7832\ : Odrv12
    port map (
            O => \N__37934\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__7831\ : LocalMux
    port map (
            O => \N__37931\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__7830\ : InMux
    port map (
            O => \N__37922\,
            I => \bfn_16_5_0_\
        );

    \I__7829\ : InMux
    port map (
            O => \N__37919\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_0\
        );

    \I__7828\ : InMux
    port map (
            O => \N__37916\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_1\
        );

    \I__7827\ : InMux
    port map (
            O => \N__37913\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_2\
        );

    \I__7826\ : InMux
    port map (
            O => \N__37910\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_3\
        );

    \I__7825\ : CascadeMux
    port map (
            O => \N__37907\,
            I => \N__37904\
        );

    \I__7824\ : InMux
    port map (
            O => \N__37904\,
            I => \N__37901\
        );

    \I__7823\ : LocalMux
    port map (
            O => \N__37901\,
            I => \N__37898\
        );

    \I__7822\ : Odrv4
    port map (
            O => \N__37898\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\
        );

    \I__7821\ : InMux
    port map (
            O => \N__37895\,
            I => \N__37892\
        );

    \I__7820\ : LocalMux
    port map (
            O => \N__37892\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\
        );

    \I__7819\ : CascadeMux
    port map (
            O => \N__37889\,
            I => \N__37886\
        );

    \I__7818\ : InMux
    port map (
            O => \N__37886\,
            I => \N__37883\
        );

    \I__7817\ : LocalMux
    port map (
            O => \N__37883\,
            I => \N__37880\
        );

    \I__7816\ : Odrv12
    port map (
            O => \N__37880\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\
        );

    \I__7815\ : CascadeMux
    port map (
            O => \N__37877\,
            I => \N__37874\
        );

    \I__7814\ : InMux
    port map (
            O => \N__37874\,
            I => \N__37871\
        );

    \I__7813\ : LocalMux
    port map (
            O => \N__37871\,
            I => \N__37868\
        );

    \I__7812\ : Span4Mux_v
    port map (
            O => \N__37868\,
            I => \N__37865\
        );

    \I__7811\ : Span4Mux_h
    port map (
            O => \N__37865\,
            I => \N__37862\
        );

    \I__7810\ : Odrv4
    port map (
            O => \N__37862\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\
        );

    \I__7809\ : InMux
    port map (
            O => \N__37859\,
            I => \N__37856\
        );

    \I__7808\ : LocalMux
    port map (
            O => \N__37856\,
            I => \N__37853\
        );

    \I__7807\ : Odrv12
    port map (
            O => \N__37853\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\
        );

    \I__7806\ : InMux
    port map (
            O => \N__37850\,
            I => \N__37847\
        );

    \I__7805\ : LocalMux
    port map (
            O => \N__37847\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\
        );

    \I__7804\ : CascadeMux
    port map (
            O => \N__37844\,
            I => \N__37841\
        );

    \I__7803\ : InMux
    port map (
            O => \N__37841\,
            I => \N__37838\
        );

    \I__7802\ : LocalMux
    port map (
            O => \N__37838\,
            I => \N__37835\
        );

    \I__7801\ : Odrv4
    port map (
            O => \N__37835\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\
        );

    \I__7800\ : InMux
    port map (
            O => \N__37832\,
            I => \N__37829\
        );

    \I__7799\ : LocalMux
    port map (
            O => \N__37829\,
            I => \N__37826\
        );

    \I__7798\ : Odrv12
    port map (
            O => \N__37826\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\
        );

    \I__7797\ : CascadeMux
    port map (
            O => \N__37823\,
            I => \N__37820\
        );

    \I__7796\ : InMux
    port map (
            O => \N__37820\,
            I => \N__37817\
        );

    \I__7795\ : LocalMux
    port map (
            O => \N__37817\,
            I => \N__37814\
        );

    \I__7794\ : Odrv4
    port map (
            O => \N__37814\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\
        );

    \I__7793\ : InMux
    port map (
            O => \N__37811\,
            I => \N__37808\
        );

    \I__7792\ : LocalMux
    port map (
            O => \N__37808\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\
        );

    \I__7791\ : CascadeMux
    port map (
            O => \N__37805\,
            I => \N__37802\
        );

    \I__7790\ : InMux
    port map (
            O => \N__37802\,
            I => \N__37799\
        );

    \I__7789\ : LocalMux
    port map (
            O => \N__37799\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\
        );

    \I__7788\ : CascadeMux
    port map (
            O => \N__37796\,
            I => \N__37793\
        );

    \I__7787\ : InMux
    port map (
            O => \N__37793\,
            I => \N__37790\
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__37790\,
            I => \N__37787\
        );

    \I__7785\ : Span4Mux_h
    port map (
            O => \N__37787\,
            I => \N__37784\
        );

    \I__7784\ : Odrv4
    port map (
            O => \N__37784\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\
        );

    \I__7783\ : InMux
    port map (
            O => \N__37781\,
            I => \N__37778\
        );

    \I__7782\ : LocalMux
    port map (
            O => \N__37778\,
            I => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\
        );

    \I__7781\ : CascadeMux
    port map (
            O => \N__37775\,
            I => \N__37772\
        );

    \I__7780\ : InMux
    port map (
            O => \N__37772\,
            I => \N__37769\
        );

    \I__7779\ : LocalMux
    port map (
            O => \N__37769\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\
        );

    \I__7778\ : InMux
    port map (
            O => \N__37766\,
            I => \N__37763\
        );

    \I__7777\ : LocalMux
    port map (
            O => \N__37763\,
            I => \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\
        );

    \I__7776\ : InMux
    port map (
            O => \N__37760\,
            I => \N__37757\
        );

    \I__7775\ : LocalMux
    port map (
            O => \N__37757\,
            I => \N__37754\
        );

    \I__7774\ : Odrv12
    port map (
            O => \N__37754\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\
        );

    \I__7773\ : InMux
    port map (
            O => \N__37751\,
            I => \N__37748\
        );

    \I__7772\ : LocalMux
    port map (
            O => \N__37748\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\
        );

    \I__7771\ : InMux
    port map (
            O => \N__37745\,
            I => \N__37742\
        );

    \I__7770\ : LocalMux
    port map (
            O => \N__37742\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\
        );

    \I__7769\ : CascadeMux
    port map (
            O => \N__37739\,
            I => \N__37736\
        );

    \I__7768\ : InMux
    port map (
            O => \N__37736\,
            I => \N__37733\
        );

    \I__7767\ : LocalMux
    port map (
            O => \N__37733\,
            I => \N__37730\
        );

    \I__7766\ : Span4Mux_h
    port map (
            O => \N__37730\,
            I => \N__37727\
        );

    \I__7765\ : Odrv4
    port map (
            O => \N__37727\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI25021_19\
        );

    \I__7764\ : InMux
    port map (
            O => \N__37724\,
            I => \N__37721\
        );

    \I__7763\ : LocalMux
    port map (
            O => \N__37721\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\
        );

    \I__7762\ : InMux
    port map (
            O => \N__37718\,
            I => \N__37715\
        );

    \I__7761\ : LocalMux
    port map (
            O => \N__37715\,
            I => \N__37712\
        );

    \I__7760\ : Span4Mux_h
    port map (
            O => \N__37712\,
            I => \N__37709\
        );

    \I__7759\ : Odrv4
    port map (
            O => \N__37709\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24\
        );

    \I__7758\ : CascadeMux
    port map (
            O => \N__37706\,
            I => \N__37703\
        );

    \I__7757\ : InMux
    port map (
            O => \N__37703\,
            I => \N__37700\
        );

    \I__7756\ : LocalMux
    port map (
            O => \N__37700\,
            I => \N__37697\
        );

    \I__7755\ : Span4Mux_v
    port map (
            O => \N__37697\,
            I => \N__37694\
        );

    \I__7754\ : Odrv4
    port map (
            O => \N__37694\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt24\
        );

    \I__7753\ : InMux
    port map (
            O => \N__37691\,
            I => \N__37688\
        );

    \I__7752\ : LocalMux
    port map (
            O => \N__37688\,
            I => \N__37685\
        );

    \I__7751\ : Span4Mux_v
    port map (
            O => \N__37685\,
            I => \N__37682\
        );

    \I__7750\ : Odrv4
    port map (
            O => \N__37682\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\
        );

    \I__7749\ : CascadeMux
    port map (
            O => \N__37679\,
            I => \N__37676\
        );

    \I__7748\ : InMux
    port map (
            O => \N__37676\,
            I => \N__37673\
        );

    \I__7747\ : LocalMux
    port map (
            O => \N__37673\,
            I => \N__37670\
        );

    \I__7746\ : Span4Mux_v
    port map (
            O => \N__37670\,
            I => \N__37667\
        );

    \I__7745\ : Odrv4
    port map (
            O => \N__37667\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt30\
        );

    \I__7744\ : InMux
    port map (
            O => \N__37664\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_30\
        );

    \I__7743\ : InMux
    port map (
            O => \N__37661\,
            I => \N__37658\
        );

    \I__7742\ : LocalMux
    port map (
            O => \N__37658\,
            I => \N__37653\
        );

    \I__7741\ : InMux
    port map (
            O => \N__37657\,
            I => \N__37648\
        );

    \I__7740\ : InMux
    port map (
            O => \N__37656\,
            I => \N__37648\
        );

    \I__7739\ : Span4Mux_v
    port map (
            O => \N__37653\,
            I => \N__37645\
        );

    \I__7738\ : LocalMux
    port map (
            O => \N__37648\,
            I => \N__37642\
        );

    \I__7737\ : Span4Mux_h
    port map (
            O => \N__37645\,
            I => \N__37637\
        );

    \I__7736\ : Span4Mux_v
    port map (
            O => \N__37642\,
            I => \N__37637\
        );

    \I__7735\ : Odrv4
    port map (
            O => \N__37637\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__7734\ : InMux
    port map (
            O => \N__37634\,
            I => \N__37631\
        );

    \I__7733\ : LocalMux
    port map (
            O => \N__37631\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\
        );

    \I__7732\ : CascadeMux
    port map (
            O => \N__37628\,
            I => \N__37625\
        );

    \I__7731\ : InMux
    port map (
            O => \N__37625\,
            I => \N__37622\
        );

    \I__7730\ : LocalMux
    port map (
            O => \N__37622\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\
        );

    \I__7729\ : CascadeMux
    port map (
            O => \N__37619\,
            I => \N__37616\
        );

    \I__7728\ : InMux
    port map (
            O => \N__37616\,
            I => \N__37613\
        );

    \I__7727\ : LocalMux
    port map (
            O => \N__37613\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\
        );

    \I__7726\ : InMux
    port map (
            O => \N__37610\,
            I => \N__37607\
        );

    \I__7725\ : LocalMux
    port map (
            O => \N__37607\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\
        );

    \I__7724\ : InMux
    port map (
            O => \N__37604\,
            I => \N__37601\
        );

    \I__7723\ : LocalMux
    port map (
            O => \N__37601\,
            I => \N__37598\
        );

    \I__7722\ : Odrv12
    port map (
            O => \N__37598\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\
        );

    \I__7721\ : InMux
    port map (
            O => \N__37595\,
            I => \N__37591\
        );

    \I__7720\ : InMux
    port map (
            O => \N__37594\,
            I => \N__37588\
        );

    \I__7719\ : LocalMux
    port map (
            O => \N__37591\,
            I => \N__37585\
        );

    \I__7718\ : LocalMux
    port map (
            O => \N__37588\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__7717\ : Odrv4
    port map (
            O => \N__37585\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__7716\ : CascadeMux
    port map (
            O => \N__37580\,
            I => \N__37577\
        );

    \I__7715\ : InMux
    port map (
            O => \N__37577\,
            I => \N__37574\
        );

    \I__7714\ : LocalMux
    port map (
            O => \N__37574\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\
        );

    \I__7713\ : InMux
    port map (
            O => \N__37571\,
            I => \N__37567\
        );

    \I__7712\ : InMux
    port map (
            O => \N__37570\,
            I => \N__37564\
        );

    \I__7711\ : LocalMux
    port map (
            O => \N__37567\,
            I => \N__37561\
        );

    \I__7710\ : LocalMux
    port map (
            O => \N__37564\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__7709\ : Odrv4
    port map (
            O => \N__37561\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__7708\ : InMux
    port map (
            O => \N__37556\,
            I => \N__37553\
        );

    \I__7707\ : LocalMux
    port map (
            O => \N__37553\,
            I => \N__37550\
        );

    \I__7706\ : Span4Mux_v
    port map (
            O => \N__37550\,
            I => \N__37547\
        );

    \I__7705\ : Odrv4
    port map (
            O => \N__37547\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\
        );

    \I__7704\ : CascadeMux
    port map (
            O => \N__37544\,
            I => \N__37541\
        );

    \I__7703\ : InMux
    port map (
            O => \N__37541\,
            I => \N__37538\
        );

    \I__7702\ : LocalMux
    port map (
            O => \N__37538\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\
        );

    \I__7701\ : InMux
    port map (
            O => \N__37535\,
            I => \N__37531\
        );

    \I__7700\ : InMux
    port map (
            O => \N__37534\,
            I => \N__37528\
        );

    \I__7699\ : LocalMux
    port map (
            O => \N__37531\,
            I => \N__37525\
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__37528\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__7697\ : Odrv4
    port map (
            O => \N__37525\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__7696\ : CascadeMux
    port map (
            O => \N__37520\,
            I => \N__37517\
        );

    \I__7695\ : InMux
    port map (
            O => \N__37517\,
            I => \N__37514\
        );

    \I__7694\ : LocalMux
    port map (
            O => \N__37514\,
            I => \N__37511\
        );

    \I__7693\ : Odrv4
    port map (
            O => \N__37511\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\
        );

    \I__7692\ : InMux
    port map (
            O => \N__37508\,
            I => \N__37505\
        );

    \I__7691\ : LocalMux
    port map (
            O => \N__37505\,
            I => \N__37502\
        );

    \I__7690\ : Span4Mux_v
    port map (
            O => \N__37502\,
            I => \N__37499\
        );

    \I__7689\ : Odrv4
    port map (
            O => \N__37499\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\
        );

    \I__7688\ : InMux
    port map (
            O => \N__37496\,
            I => \N__37492\
        );

    \I__7687\ : InMux
    port map (
            O => \N__37495\,
            I => \N__37489\
        );

    \I__7686\ : LocalMux
    port map (
            O => \N__37492\,
            I => \N__37486\
        );

    \I__7685\ : LocalMux
    port map (
            O => \N__37489\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__7684\ : Odrv4
    port map (
            O => \N__37486\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__7683\ : CascadeMux
    port map (
            O => \N__37481\,
            I => \N__37478\
        );

    \I__7682\ : InMux
    port map (
            O => \N__37478\,
            I => \N__37475\
        );

    \I__7681\ : LocalMux
    port map (
            O => \N__37475\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\
        );

    \I__7680\ : InMux
    port map (
            O => \N__37472\,
            I => \N__37469\
        );

    \I__7679\ : LocalMux
    port map (
            O => \N__37469\,
            I => \N__37466\
        );

    \I__7678\ : Odrv12
    port map (
            O => \N__37466\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt18\
        );

    \I__7677\ : CascadeMux
    port map (
            O => \N__37463\,
            I => \N__37460\
        );

    \I__7676\ : InMux
    port map (
            O => \N__37460\,
            I => \N__37457\
        );

    \I__7675\ : LocalMux
    port map (
            O => \N__37457\,
            I => \N__37454\
        );

    \I__7674\ : Odrv12
    port map (
            O => \N__37454\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\
        );

    \I__7673\ : InMux
    port map (
            O => \N__37451\,
            I => \N__37448\
        );

    \I__7672\ : LocalMux
    port map (
            O => \N__37448\,
            I => \N__37445\
        );

    \I__7671\ : Odrv12
    port map (
            O => \N__37445\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20\
        );

    \I__7670\ : CascadeMux
    port map (
            O => \N__37442\,
            I => \N__37439\
        );

    \I__7669\ : InMux
    port map (
            O => \N__37439\,
            I => \N__37436\
        );

    \I__7668\ : LocalMux
    port map (
            O => \N__37436\,
            I => \N__37433\
        );

    \I__7667\ : Span4Mux_v
    port map (
            O => \N__37433\,
            I => \N__37430\
        );

    \I__7666\ : Odrv4
    port map (
            O => \N__37430\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt20\
        );

    \I__7665\ : InMux
    port map (
            O => \N__37427\,
            I => \N__37424\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__37424\,
            I => \N__37421\
        );

    \I__7663\ : Span4Mux_v
    port map (
            O => \N__37421\,
            I => \N__37418\
        );

    \I__7662\ : Odrv4
    port map (
            O => \N__37418\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt22\
        );

    \I__7661\ : CascadeMux
    port map (
            O => \N__37415\,
            I => \N__37412\
        );

    \I__7660\ : InMux
    port map (
            O => \N__37412\,
            I => \N__37409\
        );

    \I__7659\ : LocalMux
    port map (
            O => \N__37409\,
            I => \N__37406\
        );

    \I__7658\ : Span4Mux_v
    port map (
            O => \N__37406\,
            I => \N__37403\
        );

    \I__7657\ : Odrv4
    port map (
            O => \N__37403\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22\
        );

    \I__7656\ : InMux
    port map (
            O => \N__37400\,
            I => \N__37396\
        );

    \I__7655\ : InMux
    port map (
            O => \N__37399\,
            I => \N__37393\
        );

    \I__7654\ : LocalMux
    port map (
            O => \N__37396\,
            I => \N__37390\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__37393\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__7652\ : Odrv4
    port map (
            O => \N__37390\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__7651\ : CascadeMux
    port map (
            O => \N__37385\,
            I => \N__37382\
        );

    \I__7650\ : InMux
    port map (
            O => \N__37382\,
            I => \N__37379\
        );

    \I__7649\ : LocalMux
    port map (
            O => \N__37379\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\
        );

    \I__7648\ : InMux
    port map (
            O => \N__37376\,
            I => \N__37373\
        );

    \I__7647\ : LocalMux
    port map (
            O => \N__37373\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\
        );

    \I__7646\ : InMux
    port map (
            O => \N__37370\,
            I => \N__37366\
        );

    \I__7645\ : InMux
    port map (
            O => \N__37369\,
            I => \N__37363\
        );

    \I__7644\ : LocalMux
    port map (
            O => \N__37366\,
            I => \N__37360\
        );

    \I__7643\ : LocalMux
    port map (
            O => \N__37363\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__7642\ : Odrv4
    port map (
            O => \N__37360\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__7641\ : InMux
    port map (
            O => \N__37355\,
            I => \N__37352\
        );

    \I__7640\ : LocalMux
    port map (
            O => \N__37352\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\
        );

    \I__7639\ : CascadeMux
    port map (
            O => \N__37349\,
            I => \N__37346\
        );

    \I__7638\ : InMux
    port map (
            O => \N__37346\,
            I => \N__37343\
        );

    \I__7637\ : LocalMux
    port map (
            O => \N__37343\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\
        );

    \I__7636\ : CascadeMux
    port map (
            O => \N__37340\,
            I => \N__37337\
        );

    \I__7635\ : InMux
    port map (
            O => \N__37337\,
            I => \N__37334\
        );

    \I__7634\ : LocalMux
    port map (
            O => \N__37334\,
            I => \N__37331\
        );

    \I__7633\ : Odrv4
    port map (
            O => \N__37331\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\
        );

    \I__7632\ : InMux
    port map (
            O => \N__37328\,
            I => \N__37324\
        );

    \I__7631\ : InMux
    port map (
            O => \N__37327\,
            I => \N__37321\
        );

    \I__7630\ : LocalMux
    port map (
            O => \N__37324\,
            I => \N__37318\
        );

    \I__7629\ : LocalMux
    port map (
            O => \N__37321\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__7628\ : Odrv4
    port map (
            O => \N__37318\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__7627\ : InMux
    port map (
            O => \N__37313\,
            I => \N__37310\
        );

    \I__7626\ : LocalMux
    port map (
            O => \N__37310\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\
        );

    \I__7625\ : InMux
    port map (
            O => \N__37307\,
            I => \N__37303\
        );

    \I__7624\ : InMux
    port map (
            O => \N__37306\,
            I => \N__37300\
        );

    \I__7623\ : LocalMux
    port map (
            O => \N__37303\,
            I => \N__37297\
        );

    \I__7622\ : LocalMux
    port map (
            O => \N__37300\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__7621\ : Odrv4
    port map (
            O => \N__37297\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__7620\ : InMux
    port map (
            O => \N__37292\,
            I => \N__37289\
        );

    \I__7619\ : LocalMux
    port map (
            O => \N__37289\,
            I => \N__37286\
        );

    \I__7618\ : Odrv4
    port map (
            O => \N__37286\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\
        );

    \I__7617\ : CascadeMux
    port map (
            O => \N__37283\,
            I => \N__37280\
        );

    \I__7616\ : InMux
    port map (
            O => \N__37280\,
            I => \N__37277\
        );

    \I__7615\ : LocalMux
    port map (
            O => \N__37277\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\
        );

    \I__7614\ : InMux
    port map (
            O => \N__37274\,
            I => \N__37271\
        );

    \I__7613\ : LocalMux
    port map (
            O => \N__37271\,
            I => \N__37268\
        );

    \I__7612\ : Span4Mux_h
    port map (
            O => \N__37268\,
            I => \N__37265\
        );

    \I__7611\ : Odrv4
    port map (
            O => \N__37265\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\
        );

    \I__7610\ : InMux
    port map (
            O => \N__37262\,
            I => \N__37259\
        );

    \I__7609\ : LocalMux
    port map (
            O => \N__37259\,
            I => \N__37255\
        );

    \I__7608\ : InMux
    port map (
            O => \N__37258\,
            I => \N__37252\
        );

    \I__7607\ : Span4Mux_v
    port map (
            O => \N__37255\,
            I => \N__37249\
        );

    \I__7606\ : LocalMux
    port map (
            O => \N__37252\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__7605\ : Odrv4
    port map (
            O => \N__37249\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__7604\ : CascadeMux
    port map (
            O => \N__37244\,
            I => \N__37241\
        );

    \I__7603\ : InMux
    port map (
            O => \N__37241\,
            I => \N__37238\
        );

    \I__7602\ : LocalMux
    port map (
            O => \N__37238\,
            I => \N__37235\
        );

    \I__7601\ : Odrv4
    port map (
            O => \N__37235\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\
        );

    \I__7600\ : InMux
    port map (
            O => \N__37232\,
            I => \N__37229\
        );

    \I__7599\ : LocalMux
    port map (
            O => \N__37229\,
            I => \N__37226\
        );

    \I__7598\ : Span4Mux_v
    port map (
            O => \N__37226\,
            I => \N__37223\
        );

    \I__7597\ : Odrv4
    port map (
            O => \N__37223\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\
        );

    \I__7596\ : InMux
    port map (
            O => \N__37220\,
            I => \N__37216\
        );

    \I__7595\ : InMux
    port map (
            O => \N__37219\,
            I => \N__37213\
        );

    \I__7594\ : LocalMux
    port map (
            O => \N__37216\,
            I => \N__37210\
        );

    \I__7593\ : LocalMux
    port map (
            O => \N__37213\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__7592\ : Odrv4
    port map (
            O => \N__37210\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__7591\ : CascadeMux
    port map (
            O => \N__37205\,
            I => \N__37202\
        );

    \I__7590\ : InMux
    port map (
            O => \N__37202\,
            I => \N__37199\
        );

    \I__7589\ : LocalMux
    port map (
            O => \N__37199\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\
        );

    \I__7588\ : InMux
    port map (
            O => \N__37196\,
            I => \N__37193\
        );

    \I__7587\ : LocalMux
    port map (
            O => \N__37193\,
            I => \N__37190\
        );

    \I__7586\ : Span4Mux_v
    port map (
            O => \N__37190\,
            I => \N__37187\
        );

    \I__7585\ : Odrv4
    port map (
            O => \N__37187\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\
        );

    \I__7584\ : InMux
    port map (
            O => \N__37184\,
            I => \N__37181\
        );

    \I__7583\ : LocalMux
    port map (
            O => \N__37181\,
            I => \N__37177\
        );

    \I__7582\ : InMux
    port map (
            O => \N__37180\,
            I => \N__37174\
        );

    \I__7581\ : Span4Mux_v
    port map (
            O => \N__37177\,
            I => \N__37171\
        );

    \I__7580\ : LocalMux
    port map (
            O => \N__37174\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__7579\ : Odrv4
    port map (
            O => \N__37171\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__7578\ : CascadeMux
    port map (
            O => \N__37166\,
            I => \N__37163\
        );

    \I__7577\ : InMux
    port map (
            O => \N__37163\,
            I => \N__37160\
        );

    \I__7576\ : LocalMux
    port map (
            O => \N__37160\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\
        );

    \I__7575\ : InMux
    port map (
            O => \N__37157\,
            I => \N__37153\
        );

    \I__7574\ : InMux
    port map (
            O => \N__37156\,
            I => \N__37149\
        );

    \I__7573\ : LocalMux
    port map (
            O => \N__37153\,
            I => \N__37146\
        );

    \I__7572\ : InMux
    port map (
            O => \N__37152\,
            I => \N__37143\
        );

    \I__7571\ : LocalMux
    port map (
            O => \N__37149\,
            I => \elapsed_time_ns_1_RNII43T9_0_6\
        );

    \I__7570\ : Odrv4
    port map (
            O => \N__37146\,
            I => \elapsed_time_ns_1_RNII43T9_0_6\
        );

    \I__7569\ : LocalMux
    port map (
            O => \N__37143\,
            I => \elapsed_time_ns_1_RNII43T9_0_6\
        );

    \I__7568\ : CascadeMux
    port map (
            O => \N__37136\,
            I => \N__37133\
        );

    \I__7567\ : InMux
    port map (
            O => \N__37133\,
            I => \N__37130\
        );

    \I__7566\ : LocalMux
    port map (
            O => \N__37130\,
            I => \N__37127\
        );

    \I__7565\ : Odrv12
    port map (
            O => \N__37127\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\
        );

    \I__7564\ : CascadeMux
    port map (
            O => \N__37124\,
            I => \N__37121\
        );

    \I__7563\ : InMux
    port map (
            O => \N__37121\,
            I => \N__37118\
        );

    \I__7562\ : LocalMux
    port map (
            O => \N__37118\,
            I => \N__37113\
        );

    \I__7561\ : InMux
    port map (
            O => \N__37117\,
            I => \N__37110\
        );

    \I__7560\ : InMux
    port map (
            O => \N__37116\,
            I => \N__37107\
        );

    \I__7559\ : Span4Mux_h
    port map (
            O => \N__37113\,
            I => \N__37104\
        );

    \I__7558\ : LocalMux
    port map (
            O => \N__37110\,
            I => \N__37101\
        );

    \I__7557\ : LocalMux
    port map (
            O => \N__37107\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__7556\ : Odrv4
    port map (
            O => \N__37104\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__7555\ : Odrv4
    port map (
            O => \N__37101\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__7554\ : InMux
    port map (
            O => \N__37094\,
            I => \N__37091\
        );

    \I__7553\ : LocalMux
    port map (
            O => \N__37091\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\
        );

    \I__7552\ : InMux
    port map (
            O => \N__37088\,
            I => \N__37084\
        );

    \I__7551\ : InMux
    port map (
            O => \N__37087\,
            I => \N__37081\
        );

    \I__7550\ : LocalMux
    port map (
            O => \N__37084\,
            I => \N__37078\
        );

    \I__7549\ : LocalMux
    port map (
            O => \N__37081\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__7548\ : Odrv4
    port map (
            O => \N__37078\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__7547\ : CascadeMux
    port map (
            O => \N__37073\,
            I => \N__37070\
        );

    \I__7546\ : InMux
    port map (
            O => \N__37070\,
            I => \N__37067\
        );

    \I__7545\ : LocalMux
    port map (
            O => \N__37067\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\
        );

    \I__7544\ : InMux
    port map (
            O => \N__37064\,
            I => \N__37061\
        );

    \I__7543\ : LocalMux
    port map (
            O => \N__37061\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\
        );

    \I__7542\ : InMux
    port map (
            O => \N__37058\,
            I => \N__37055\
        );

    \I__7541\ : LocalMux
    port map (
            O => \N__37055\,
            I => \N__37051\
        );

    \I__7540\ : InMux
    port map (
            O => \N__37054\,
            I => \N__37048\
        );

    \I__7539\ : Span4Mux_v
    port map (
            O => \N__37051\,
            I => \N__37045\
        );

    \I__7538\ : LocalMux
    port map (
            O => \N__37048\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__7537\ : Odrv4
    port map (
            O => \N__37045\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__7536\ : CascadeMux
    port map (
            O => \N__37040\,
            I => \N__37037\
        );

    \I__7535\ : InMux
    port map (
            O => \N__37037\,
            I => \N__37034\
        );

    \I__7534\ : LocalMux
    port map (
            O => \N__37034\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\
        );

    \I__7533\ : InMux
    port map (
            O => \N__37031\,
            I => \N__37028\
        );

    \I__7532\ : LocalMux
    port map (
            O => \N__37028\,
            I => \N__37024\
        );

    \I__7531\ : InMux
    port map (
            O => \N__37027\,
            I => \N__37021\
        );

    \I__7530\ : Span4Mux_v
    port map (
            O => \N__37024\,
            I => \N__37018\
        );

    \I__7529\ : LocalMux
    port map (
            O => \N__37021\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__7528\ : Odrv4
    port map (
            O => \N__37018\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__7527\ : InMux
    port map (
            O => \N__37013\,
            I => \N__37010\
        );

    \I__7526\ : LocalMux
    port map (
            O => \N__37010\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\
        );

    \I__7525\ : CascadeMux
    port map (
            O => \N__37007\,
            I => \N__37004\
        );

    \I__7524\ : InMux
    port map (
            O => \N__37004\,
            I => \N__37001\
        );

    \I__7523\ : LocalMux
    port map (
            O => \N__37001\,
            I => \N__36998\
        );

    \I__7522\ : Odrv4
    port map (
            O => \N__36998\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\
        );

    \I__7521\ : CascadeMux
    port map (
            O => \N__36995\,
            I => \N__36992\
        );

    \I__7520\ : InMux
    port map (
            O => \N__36992\,
            I => \N__36988\
        );

    \I__7519\ : InMux
    port map (
            O => \N__36991\,
            I => \N__36984\
        );

    \I__7518\ : LocalMux
    port map (
            O => \N__36988\,
            I => \N__36981\
        );

    \I__7517\ : InMux
    port map (
            O => \N__36987\,
            I => \N__36978\
        );

    \I__7516\ : LocalMux
    port map (
            O => \N__36984\,
            I => \N__36975\
        );

    \I__7515\ : Span4Mux_h
    port map (
            O => \N__36981\,
            I => \N__36972\
        );

    \I__7514\ : LocalMux
    port map (
            O => \N__36978\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11\
        );

    \I__7513\ : Odrv4
    port map (
            O => \N__36975\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11\
        );

    \I__7512\ : Odrv4
    port map (
            O => \N__36972\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11\
        );

    \I__7511\ : CascadeMux
    port map (
            O => \N__36965\,
            I => \N__36961\
        );

    \I__7510\ : InMux
    port map (
            O => \N__36964\,
            I => \N__36955\
        );

    \I__7509\ : InMux
    port map (
            O => \N__36961\,
            I => \N__36955\
        );

    \I__7508\ : InMux
    port map (
            O => \N__36960\,
            I => \N__36952\
        );

    \I__7507\ : LocalMux
    port map (
            O => \N__36955\,
            I => \N__36949\
        );

    \I__7506\ : LocalMux
    port map (
            O => \N__36952\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__7505\ : Odrv4
    port map (
            O => \N__36949\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__7504\ : CascadeMux
    port map (
            O => \N__36944\,
            I => \N__36941\
        );

    \I__7503\ : InMux
    port map (
            O => \N__36941\,
            I => \N__36937\
        );

    \I__7502\ : InMux
    port map (
            O => \N__36940\,
            I => \N__36934\
        );

    \I__7501\ : LocalMux
    port map (
            O => \N__36937\,
            I => \N__36928\
        );

    \I__7500\ : LocalMux
    port map (
            O => \N__36934\,
            I => \N__36928\
        );

    \I__7499\ : InMux
    port map (
            O => \N__36933\,
            I => \N__36925\
        );

    \I__7498\ : Span4Mux_v
    port map (
            O => \N__36928\,
            I => \N__36922\
        );

    \I__7497\ : LocalMux
    port map (
            O => \N__36925\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__7496\ : Odrv4
    port map (
            O => \N__36922\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__7495\ : InMux
    port map (
            O => \N__36917\,
            I => \N__36913\
        );

    \I__7494\ : InMux
    port map (
            O => \N__36916\,
            I => \N__36910\
        );

    \I__7493\ : LocalMux
    port map (
            O => \N__36913\,
            I => \N__36905\
        );

    \I__7492\ : LocalMux
    port map (
            O => \N__36910\,
            I => \N__36905\
        );

    \I__7491\ : Odrv4
    port map (
            O => \N__36905\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_21\
        );

    \I__7490\ : InMux
    port map (
            O => \N__36902\,
            I => \N__36896\
        );

    \I__7489\ : InMux
    port map (
            O => \N__36901\,
            I => \N__36896\
        );

    \I__7488\ : LocalMux
    port map (
            O => \N__36896\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_20\
        );

    \I__7487\ : InMux
    port map (
            O => \N__36893\,
            I => \N__36889\
        );

    \I__7486\ : InMux
    port map (
            O => \N__36892\,
            I => \N__36886\
        );

    \I__7485\ : LocalMux
    port map (
            O => \N__36889\,
            I => \N__36880\
        );

    \I__7484\ : LocalMux
    port map (
            O => \N__36886\,
            I => \N__36880\
        );

    \I__7483\ : InMux
    port map (
            O => \N__36885\,
            I => \N__36877\
        );

    \I__7482\ : Span4Mux_v
    port map (
            O => \N__36880\,
            I => \N__36874\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__36877\,
            I => \elapsed_time_ns_1_RNIL73T9_0_9\
        );

    \I__7480\ : Odrv4
    port map (
            O => \N__36874\,
            I => \elapsed_time_ns_1_RNIL73T9_0_9\
        );

    \I__7479\ : CascadeMux
    port map (
            O => \N__36869\,
            I => \N__36865\
        );

    \I__7478\ : InMux
    port map (
            O => \N__36868\,
            I => \N__36860\
        );

    \I__7477\ : InMux
    port map (
            O => \N__36865\,
            I => \N__36860\
        );

    \I__7476\ : LocalMux
    port map (
            O => \N__36860\,
            I => \N__36857\
        );

    \I__7475\ : Span4Mux_v
    port map (
            O => \N__36857\,
            I => \N__36854\
        );

    \I__7474\ : Odrv4
    port map (
            O => \N__36854\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\
        );

    \I__7473\ : CascadeMux
    port map (
            O => \N__36851\,
            I => \N__36846\
        );

    \I__7472\ : InMux
    port map (
            O => \N__36850\,
            I => \N__36843\
        );

    \I__7471\ : InMux
    port map (
            O => \N__36849\,
            I => \N__36838\
        );

    \I__7470\ : InMux
    port map (
            O => \N__36846\,
            I => \N__36838\
        );

    \I__7469\ : LocalMux
    port map (
            O => \N__36843\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__7468\ : LocalMux
    port map (
            O => \N__36838\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__7467\ : InMux
    port map (
            O => \N__36833\,
            I => \N__36828\
        );

    \I__7466\ : InMux
    port map (
            O => \N__36832\,
            I => \N__36823\
        );

    \I__7465\ : InMux
    port map (
            O => \N__36831\,
            I => \N__36823\
        );

    \I__7464\ : LocalMux
    port map (
            O => \N__36828\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__7463\ : LocalMux
    port map (
            O => \N__36823\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__7462\ : InMux
    port map (
            O => \N__36818\,
            I => \N__36815\
        );

    \I__7461\ : LocalMux
    port map (
            O => \N__36815\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\
        );

    \I__7460\ : CascadeMux
    port map (
            O => \N__36812\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20_cascade_\
        );

    \I__7459\ : InMux
    port map (
            O => \N__36809\,
            I => \N__36806\
        );

    \I__7458\ : LocalMux
    port map (
            O => \N__36806\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\
        );

    \I__7457\ : InMux
    port map (
            O => \N__36803\,
            I => \N__36800\
        );

    \I__7456\ : LocalMux
    port map (
            O => \N__36800\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19\
        );

    \I__7455\ : CascadeMux
    port map (
            O => \N__36797\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_\
        );

    \I__7454\ : InMux
    port map (
            O => \N__36794\,
            I => \N__36791\
        );

    \I__7453\ : LocalMux
    port map (
            O => \N__36791\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3\
        );

    \I__7452\ : InMux
    port map (
            O => \N__36788\,
            I => \N__36785\
        );

    \I__7451\ : LocalMux
    port map (
            O => \N__36785\,
            I => \N__36782\
        );

    \I__7450\ : Span4Mux_v
    port map (
            O => \N__36782\,
            I => \N__36778\
        );

    \I__7449\ : InMux
    port map (
            O => \N__36781\,
            I => \N__36775\
        );

    \I__7448\ : Odrv4
    port map (
            O => \N__36778\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10\
        );

    \I__7447\ : LocalMux
    port map (
            O => \N__36775\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10\
        );

    \I__7446\ : CascadeMux
    port map (
            O => \N__36770\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10_cascade_\
        );

    \I__7445\ : CascadeMux
    port map (
            O => \N__36767\,
            I => \N__36764\
        );

    \I__7444\ : InMux
    port map (
            O => \N__36764\,
            I => \N__36761\
        );

    \I__7443\ : LocalMux
    port map (
            O => \N__36761\,
            I => \N__36758\
        );

    \I__7442\ : Span4Mux_v
    port map (
            O => \N__36758\,
            I => \N__36755\
        );

    \I__7441\ : Odrv4
    port map (
            O => \N__36755\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\
        );

    \I__7440\ : InMux
    port map (
            O => \N__36752\,
            I => \N__36744\
        );

    \I__7439\ : InMux
    port map (
            O => \N__36751\,
            I => \N__36744\
        );

    \I__7438\ : InMux
    port map (
            O => \N__36750\,
            I => \N__36741\
        );

    \I__7437\ : InMux
    port map (
            O => \N__36749\,
            I => \N__36738\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__36744\,
            I => \N__36733\
        );

    \I__7435\ : LocalMux
    port map (
            O => \N__36741\,
            I => \N__36733\
        );

    \I__7434\ : LocalMux
    port map (
            O => \N__36738\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__7433\ : Odrv4
    port map (
            O => \N__36733\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__7432\ : InMux
    port map (
            O => \N__36728\,
            I => \N__36720\
        );

    \I__7431\ : InMux
    port map (
            O => \N__36727\,
            I => \N__36720\
        );

    \I__7430\ : InMux
    port map (
            O => \N__36726\,
            I => \N__36717\
        );

    \I__7429\ : InMux
    port map (
            O => \N__36725\,
            I => \N__36714\
        );

    \I__7428\ : LocalMux
    port map (
            O => \N__36720\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__7427\ : LocalMux
    port map (
            O => \N__36717\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__7426\ : LocalMux
    port map (
            O => \N__36714\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__7425\ : CascadeMux
    port map (
            O => \N__36707\,
            I => \N__36704\
        );

    \I__7424\ : InMux
    port map (
            O => \N__36704\,
            I => \N__36701\
        );

    \I__7423\ : LocalMux
    port map (
            O => \N__36701\,
            I => \N__36698\
        );

    \I__7422\ : Span4Mux_v
    port map (
            O => \N__36698\,
            I => \N__36695\
        );

    \I__7421\ : Odrv4
    port map (
            O => \N__36695\,
            I => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\
        );

    \I__7420\ : InMux
    port map (
            O => \N__36692\,
            I => \N__36689\
        );

    \I__7419\ : LocalMux
    port map (
            O => \N__36689\,
            I => \N__36686\
        );

    \I__7418\ : Span4Mux_v
    port map (
            O => \N__36686\,
            I => \N__36681\
        );

    \I__7417\ : InMux
    port map (
            O => \N__36685\,
            I => \N__36678\
        );

    \I__7416\ : InMux
    port map (
            O => \N__36684\,
            I => \N__36675\
        );

    \I__7415\ : Span4Mux_v
    port map (
            O => \N__36681\,
            I => \N__36670\
        );

    \I__7414\ : LocalMux
    port map (
            O => \N__36678\,
            I => \N__36670\
        );

    \I__7413\ : LocalMux
    port map (
            O => \N__36675\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__7412\ : Odrv4
    port map (
            O => \N__36670\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__7411\ : InMux
    port map (
            O => \N__36665\,
            I => \N__36662\
        );

    \I__7410\ : LocalMux
    port map (
            O => \N__36662\,
            I => \current_shift_inst.un38_control_input_0_s1_27\
        );

    \I__7409\ : InMux
    port map (
            O => \N__36659\,
            I => \current_shift_inst.un38_control_input_cry_26_s1\
        );

    \I__7408\ : InMux
    port map (
            O => \N__36656\,
            I => \N__36653\
        );

    \I__7407\ : LocalMux
    port map (
            O => \N__36653\,
            I => \current_shift_inst.un38_control_input_0_s1_28\
        );

    \I__7406\ : InMux
    port map (
            O => \N__36650\,
            I => \current_shift_inst.un38_control_input_cry_27_s1\
        );

    \I__7405\ : InMux
    port map (
            O => \N__36647\,
            I => \N__36644\
        );

    \I__7404\ : LocalMux
    port map (
            O => \N__36644\,
            I => \current_shift_inst.un38_control_input_0_s1_29\
        );

    \I__7403\ : InMux
    port map (
            O => \N__36641\,
            I => \current_shift_inst.un38_control_input_cry_28_s1\
        );

    \I__7402\ : InMux
    port map (
            O => \N__36638\,
            I => \N__36635\
        );

    \I__7401\ : LocalMux
    port map (
            O => \N__36635\,
            I => \N__36632\
        );

    \I__7400\ : Odrv4
    port map (
            O => \N__36632\,
            I => \current_shift_inst.un38_control_input_0_s1_30\
        );

    \I__7399\ : InMux
    port map (
            O => \N__36629\,
            I => \current_shift_inst.un38_control_input_cry_29_s1\
        );

    \I__7398\ : InMux
    port map (
            O => \N__36626\,
            I => \current_shift_inst.un38_control_input_cry_30_s1\
        );

    \I__7397\ : InMux
    port map (
            O => \N__36623\,
            I => \N__36620\
        );

    \I__7396\ : LocalMux
    port map (
            O => \N__36620\,
            I => \N__36617\
        );

    \I__7395\ : Span4Mux_h
    port map (
            O => \N__36617\,
            I => \N__36614\
        );

    \I__7394\ : Odrv4
    port map (
            O => \N__36614\,
            I => \current_shift_inst.un38_control_input_0_s1_31\
        );

    \I__7393\ : InMux
    port map (
            O => \N__36611\,
            I => \N__36608\
        );

    \I__7392\ : LocalMux
    port map (
            O => \N__36608\,
            I => \N__36605\
        );

    \I__7391\ : Span4Mux_v
    port map (
            O => \N__36605\,
            I => \N__36602\
        );

    \I__7390\ : Odrv4
    port map (
            O => \N__36602\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4\
        );

    \I__7389\ : InMux
    port map (
            O => \N__36599\,
            I => \N__36596\
        );

    \I__7388\ : LocalMux
    port map (
            O => \N__36596\,
            I => \N__36593\
        );

    \I__7387\ : Span4Mux_v
    port map (
            O => \N__36593\,
            I => \N__36590\
        );

    \I__7386\ : Odrv4
    port map (
            O => \N__36590\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI00M61_4\
        );

    \I__7385\ : InMux
    port map (
            O => \N__36587\,
            I => \N__36584\
        );

    \I__7384\ : LocalMux
    port map (
            O => \N__36584\,
            I => \current_shift_inst.un38_control_input_0_s1_18\
        );

    \I__7383\ : InMux
    port map (
            O => \N__36581\,
            I => \current_shift_inst.un38_control_input_cry_17_s1\
        );

    \I__7382\ : InMux
    port map (
            O => \N__36578\,
            I => \N__36575\
        );

    \I__7381\ : LocalMux
    port map (
            O => \N__36575\,
            I => \current_shift_inst.un38_control_input_0_s1_19\
        );

    \I__7380\ : InMux
    port map (
            O => \N__36572\,
            I => \current_shift_inst.un38_control_input_cry_18_s1\
        );

    \I__7379\ : InMux
    port map (
            O => \N__36569\,
            I => \N__36566\
        );

    \I__7378\ : LocalMux
    port map (
            O => \N__36566\,
            I => \N__36563\
        );

    \I__7377\ : Span4Mux_h
    port map (
            O => \N__36563\,
            I => \N__36560\
        );

    \I__7376\ : Odrv4
    port map (
            O => \N__36560\,
            I => \current_shift_inst.un38_control_input_0_s1_20\
        );

    \I__7375\ : InMux
    port map (
            O => \N__36557\,
            I => \current_shift_inst.un38_control_input_cry_19_s1\
        );

    \I__7374\ : InMux
    port map (
            O => \N__36554\,
            I => \N__36551\
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__36551\,
            I => \N__36548\
        );

    \I__7372\ : Span4Mux_h
    port map (
            O => \N__36548\,
            I => \N__36545\
        );

    \I__7371\ : Odrv4
    port map (
            O => \N__36545\,
            I => \current_shift_inst.un38_control_input_0_s1_21\
        );

    \I__7370\ : InMux
    port map (
            O => \N__36542\,
            I => \current_shift_inst.un38_control_input_cry_20_s1\
        );

    \I__7369\ : CascadeMux
    port map (
            O => \N__36539\,
            I => \N__36536\
        );

    \I__7368\ : InMux
    port map (
            O => \N__36536\,
            I => \N__36533\
        );

    \I__7367\ : LocalMux
    port map (
            O => \N__36533\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\
        );

    \I__7366\ : InMux
    port map (
            O => \N__36530\,
            I => \N__36527\
        );

    \I__7365\ : LocalMux
    port map (
            O => \N__36527\,
            I => \N__36524\
        );

    \I__7364\ : Odrv12
    port map (
            O => \N__36524\,
            I => \current_shift_inst.un38_control_input_0_s1_22\
        );

    \I__7363\ : InMux
    port map (
            O => \N__36521\,
            I => \current_shift_inst.un38_control_input_cry_21_s1\
        );

    \I__7362\ : InMux
    port map (
            O => \N__36518\,
            I => \N__36515\
        );

    \I__7361\ : LocalMux
    port map (
            O => \N__36515\,
            I => \N__36512\
        );

    \I__7360\ : Odrv4
    port map (
            O => \N__36512\,
            I => \current_shift_inst.un38_control_input_0_s1_23\
        );

    \I__7359\ : InMux
    port map (
            O => \N__36509\,
            I => \current_shift_inst.un38_control_input_cry_22_s1\
        );

    \I__7358\ : InMux
    port map (
            O => \N__36506\,
            I => \N__36503\
        );

    \I__7357\ : LocalMux
    port map (
            O => \N__36503\,
            I => \N__36500\
        );

    \I__7356\ : Span4Mux_h
    port map (
            O => \N__36500\,
            I => \N__36497\
        );

    \I__7355\ : Odrv4
    port map (
            O => \N__36497\,
            I => \current_shift_inst.un38_control_input_0_s1_24\
        );

    \I__7354\ : InMux
    port map (
            O => \N__36494\,
            I => \bfn_14_18_0_\
        );

    \I__7353\ : InMux
    port map (
            O => \N__36491\,
            I => \N__36488\
        );

    \I__7352\ : LocalMux
    port map (
            O => \N__36488\,
            I => \current_shift_inst.un38_control_input_0_s1_25\
        );

    \I__7351\ : InMux
    port map (
            O => \N__36485\,
            I => \current_shift_inst.un38_control_input_cry_24_s1\
        );

    \I__7350\ : InMux
    port map (
            O => \N__36482\,
            I => \N__36479\
        );

    \I__7349\ : LocalMux
    port map (
            O => \N__36479\,
            I => \current_shift_inst.un38_control_input_0_s1_26\
        );

    \I__7348\ : InMux
    port map (
            O => \N__36476\,
            I => \current_shift_inst.un38_control_input_cry_25_s1\
        );

    \I__7347\ : InMux
    port map (
            O => \N__36473\,
            I => \N__36470\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__36470\,
            I => \current_shift_inst.un38_control_input_0_s1_10\
        );

    \I__7345\ : InMux
    port map (
            O => \N__36467\,
            I => \current_shift_inst.un38_control_input_cry_9_s1\
        );

    \I__7344\ : InMux
    port map (
            O => \N__36464\,
            I => \N__36461\
        );

    \I__7343\ : LocalMux
    port map (
            O => \N__36461\,
            I => \N__36458\
        );

    \I__7342\ : Span4Mux_v
    port map (
            O => \N__36458\,
            I => \N__36455\
        );

    \I__7341\ : Odrv4
    port map (
            O => \N__36455\,
            I => \current_shift_inst.un38_control_input_0_s1_11\
        );

    \I__7340\ : InMux
    port map (
            O => \N__36452\,
            I => \current_shift_inst.un38_control_input_cry_10_s1\
        );

    \I__7339\ : InMux
    port map (
            O => \N__36449\,
            I => \N__36446\
        );

    \I__7338\ : LocalMux
    port map (
            O => \N__36446\,
            I => \N__36443\
        );

    \I__7337\ : Span4Mux_h
    port map (
            O => \N__36443\,
            I => \N__36440\
        );

    \I__7336\ : Odrv4
    port map (
            O => \N__36440\,
            I => \current_shift_inst.un38_control_input_0_s1_12\
        );

    \I__7335\ : InMux
    port map (
            O => \N__36437\,
            I => \current_shift_inst.un38_control_input_cry_11_s1\
        );

    \I__7334\ : InMux
    port map (
            O => \N__36434\,
            I => \N__36431\
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__36431\,
            I => \N__36428\
        );

    \I__7332\ : Odrv12
    port map (
            O => \N__36428\,
            I => \current_shift_inst.un38_control_input_0_s1_13\
        );

    \I__7331\ : InMux
    port map (
            O => \N__36425\,
            I => \current_shift_inst.un38_control_input_cry_12_s1\
        );

    \I__7330\ : InMux
    port map (
            O => \N__36422\,
            I => \N__36419\
        );

    \I__7329\ : LocalMux
    port map (
            O => \N__36419\,
            I => \current_shift_inst.un38_control_input_0_s1_14\
        );

    \I__7328\ : InMux
    port map (
            O => \N__36416\,
            I => \current_shift_inst.un38_control_input_cry_13_s1\
        );

    \I__7327\ : InMux
    port map (
            O => \N__36413\,
            I => \N__36410\
        );

    \I__7326\ : LocalMux
    port map (
            O => \N__36410\,
            I => \current_shift_inst.un38_control_input_0_s1_15\
        );

    \I__7325\ : InMux
    port map (
            O => \N__36407\,
            I => \current_shift_inst.un38_control_input_cry_14_s1\
        );

    \I__7324\ : InMux
    port map (
            O => \N__36404\,
            I => \N__36401\
        );

    \I__7323\ : LocalMux
    port map (
            O => \N__36401\,
            I => \current_shift_inst.un38_control_input_0_s1_16\
        );

    \I__7322\ : InMux
    port map (
            O => \N__36398\,
            I => \bfn_14_17_0_\
        );

    \I__7321\ : InMux
    port map (
            O => \N__36395\,
            I => \N__36392\
        );

    \I__7320\ : LocalMux
    port map (
            O => \N__36392\,
            I => \current_shift_inst.un38_control_input_0_s1_17\
        );

    \I__7319\ : InMux
    port map (
            O => \N__36389\,
            I => \current_shift_inst.un38_control_input_cry_16_s1\
        );

    \I__7318\ : InMux
    port map (
            O => \N__36386\,
            I => \N__36383\
        );

    \I__7317\ : LocalMux
    port map (
            O => \N__36383\,
            I => \N__36380\
        );

    \I__7316\ : Odrv12
    port map (
            O => \N__36380\,
            I => \current_shift_inst.un38_control_input_0_s1_3\
        );

    \I__7315\ : InMux
    port map (
            O => \N__36377\,
            I => \current_shift_inst.un38_control_input_cry_2_s1\
        );

    \I__7314\ : InMux
    port map (
            O => \N__36374\,
            I => \N__36371\
        );

    \I__7313\ : LocalMux
    port map (
            O => \N__36371\,
            I => \N__36368\
        );

    \I__7312\ : Odrv4
    port map (
            O => \N__36368\,
            I => \current_shift_inst.un38_control_input_0_s1_4\
        );

    \I__7311\ : InMux
    port map (
            O => \N__36365\,
            I => \current_shift_inst.un38_control_input_cry_3_s1\
        );

    \I__7310\ : InMux
    port map (
            O => \N__36362\,
            I => \N__36359\
        );

    \I__7309\ : LocalMux
    port map (
            O => \N__36359\,
            I => \N__36356\
        );

    \I__7308\ : Odrv4
    port map (
            O => \N__36356\,
            I => \current_shift_inst.un38_control_input_0_s1_5\
        );

    \I__7307\ : InMux
    port map (
            O => \N__36353\,
            I => \current_shift_inst.un38_control_input_cry_4_s1\
        );

    \I__7306\ : CascadeMux
    port map (
            O => \N__36350\,
            I => \N__36347\
        );

    \I__7305\ : InMux
    port map (
            O => \N__36347\,
            I => \N__36344\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__36344\,
            I => \N__36341\
        );

    \I__7303\ : Span4Mux_h
    port map (
            O => \N__36341\,
            I => \N__36338\
        );

    \I__7302\ : Odrv4
    port map (
            O => \N__36338\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\
        );

    \I__7301\ : InMux
    port map (
            O => \N__36335\,
            I => \N__36332\
        );

    \I__7300\ : LocalMux
    port map (
            O => \N__36332\,
            I => \N__36329\
        );

    \I__7299\ : Odrv12
    port map (
            O => \N__36329\,
            I => \current_shift_inst.un38_control_input_0_s1_6\
        );

    \I__7298\ : InMux
    port map (
            O => \N__36326\,
            I => \current_shift_inst.un38_control_input_cry_5_s1\
        );

    \I__7297\ : InMux
    port map (
            O => \N__36323\,
            I => \N__36320\
        );

    \I__7296\ : LocalMux
    port map (
            O => \N__36320\,
            I => \N__36317\
        );

    \I__7295\ : Odrv4
    port map (
            O => \N__36317\,
            I => \current_shift_inst.un38_control_input_0_s1_7\
        );

    \I__7294\ : InMux
    port map (
            O => \N__36314\,
            I => \current_shift_inst.un38_control_input_cry_6_s1\
        );

    \I__7293\ : InMux
    port map (
            O => \N__36311\,
            I => \N__36308\
        );

    \I__7292\ : LocalMux
    port map (
            O => \N__36308\,
            I => \N__36305\
        );

    \I__7291\ : Span4Mux_v
    port map (
            O => \N__36305\,
            I => \N__36302\
        );

    \I__7290\ : Odrv4
    port map (
            O => \N__36302\,
            I => \current_shift_inst.un38_control_input_0_s1_8\
        );

    \I__7289\ : InMux
    port map (
            O => \N__36299\,
            I => \bfn_14_16_0_\
        );

    \I__7288\ : InMux
    port map (
            O => \N__36296\,
            I => \N__36293\
        );

    \I__7287\ : LocalMux
    port map (
            O => \N__36293\,
            I => \N__36290\
        );

    \I__7286\ : Span4Mux_v
    port map (
            O => \N__36290\,
            I => \N__36287\
        );

    \I__7285\ : Span4Mux_h
    port map (
            O => \N__36287\,
            I => \N__36284\
        );

    \I__7284\ : Odrv4
    port map (
            O => \N__36284\,
            I => \current_shift_inst.un38_control_input_0_s1_9\
        );

    \I__7283\ : InMux
    port map (
            O => \N__36281\,
            I => \current_shift_inst.un38_control_input_cry_8_s1\
        );

    \I__7282\ : InMux
    port map (
            O => \N__36278\,
            I => \N__36273\
        );

    \I__7281\ : InMux
    port map (
            O => \N__36277\,
            I => \N__36268\
        );

    \I__7280\ : InMux
    port map (
            O => \N__36276\,
            I => \N__36268\
        );

    \I__7279\ : LocalMux
    port map (
            O => \N__36273\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__7278\ : LocalMux
    port map (
            O => \N__36268\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__7277\ : InMux
    port map (
            O => \N__36263\,
            I => \bfn_14_14_0_\
        );

    \I__7276\ : InMux
    port map (
            O => \N__36260\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\
        );

    \I__7275\ : InMux
    port map (
            O => \N__36257\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\
        );

    \I__7274\ : InMux
    port map (
            O => \N__36254\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\
        );

    \I__7273\ : InMux
    port map (
            O => \N__36251\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\
        );

    \I__7272\ : InMux
    port map (
            O => \N__36248\,
            I => \N__36243\
        );

    \I__7271\ : InMux
    port map (
            O => \N__36247\,
            I => \N__36238\
        );

    \I__7270\ : InMux
    port map (
            O => \N__36246\,
            I => \N__36238\
        );

    \I__7269\ : LocalMux
    port map (
            O => \N__36243\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__7268\ : LocalMux
    port map (
            O => \N__36238\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__7267\ : InMux
    port map (
            O => \N__36233\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\
        );

    \I__7266\ : IoInMux
    port map (
            O => \N__36230\,
            I => \N__36213\
        );

    \I__7265\ : InMux
    port map (
            O => \N__36229\,
            I => \N__36206\
        );

    \I__7264\ : InMux
    port map (
            O => \N__36228\,
            I => \N__36206\
        );

    \I__7263\ : InMux
    port map (
            O => \N__36227\,
            I => \N__36206\
        );

    \I__7262\ : InMux
    port map (
            O => \N__36226\,
            I => \N__36197\
        );

    \I__7261\ : InMux
    port map (
            O => \N__36225\,
            I => \N__36197\
        );

    \I__7260\ : InMux
    port map (
            O => \N__36224\,
            I => \N__36197\
        );

    \I__7259\ : InMux
    port map (
            O => \N__36223\,
            I => \N__36197\
        );

    \I__7258\ : InMux
    port map (
            O => \N__36222\,
            I => \N__36186\
        );

    \I__7257\ : InMux
    port map (
            O => \N__36221\,
            I => \N__36186\
        );

    \I__7256\ : InMux
    port map (
            O => \N__36220\,
            I => \N__36186\
        );

    \I__7255\ : InMux
    port map (
            O => \N__36219\,
            I => \N__36177\
        );

    \I__7254\ : InMux
    port map (
            O => \N__36218\,
            I => \N__36177\
        );

    \I__7253\ : InMux
    port map (
            O => \N__36217\,
            I => \N__36177\
        );

    \I__7252\ : InMux
    port map (
            O => \N__36216\,
            I => \N__36177\
        );

    \I__7251\ : LocalMux
    port map (
            O => \N__36213\,
            I => \N__36170\
        );

    \I__7250\ : LocalMux
    port map (
            O => \N__36206\,
            I => \N__36158\
        );

    \I__7249\ : LocalMux
    port map (
            O => \N__36197\,
            I => \N__36155\
        );

    \I__7248\ : InMux
    port map (
            O => \N__36196\,
            I => \N__36146\
        );

    \I__7247\ : InMux
    port map (
            O => \N__36195\,
            I => \N__36146\
        );

    \I__7246\ : InMux
    port map (
            O => \N__36194\,
            I => \N__36146\
        );

    \I__7245\ : InMux
    port map (
            O => \N__36193\,
            I => \N__36146\
        );

    \I__7244\ : LocalMux
    port map (
            O => \N__36186\,
            I => \N__36141\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__36177\,
            I => \N__36141\
        );

    \I__7242\ : InMux
    port map (
            O => \N__36176\,
            I => \N__36132\
        );

    \I__7241\ : InMux
    port map (
            O => \N__36175\,
            I => \N__36132\
        );

    \I__7240\ : InMux
    port map (
            O => \N__36174\,
            I => \N__36132\
        );

    \I__7239\ : InMux
    port map (
            O => \N__36173\,
            I => \N__36132\
        );

    \I__7238\ : IoSpan4Mux
    port map (
            O => \N__36170\,
            I => \N__36129\
        );

    \I__7237\ : InMux
    port map (
            O => \N__36169\,
            I => \N__36126\
        );

    \I__7236\ : InMux
    port map (
            O => \N__36168\,
            I => \N__36117\
        );

    \I__7235\ : InMux
    port map (
            O => \N__36167\,
            I => \N__36117\
        );

    \I__7234\ : InMux
    port map (
            O => \N__36166\,
            I => \N__36117\
        );

    \I__7233\ : InMux
    port map (
            O => \N__36165\,
            I => \N__36117\
        );

    \I__7232\ : InMux
    port map (
            O => \N__36164\,
            I => \N__36108\
        );

    \I__7231\ : InMux
    port map (
            O => \N__36163\,
            I => \N__36108\
        );

    \I__7230\ : InMux
    port map (
            O => \N__36162\,
            I => \N__36108\
        );

    \I__7229\ : InMux
    port map (
            O => \N__36161\,
            I => \N__36108\
        );

    \I__7228\ : Span4Mux_v
    port map (
            O => \N__36158\,
            I => \N__36097\
        );

    \I__7227\ : Span4Mux_v
    port map (
            O => \N__36155\,
            I => \N__36097\
        );

    \I__7226\ : LocalMux
    port map (
            O => \N__36146\,
            I => \N__36097\
        );

    \I__7225\ : Span4Mux_v
    port map (
            O => \N__36141\,
            I => \N__36097\
        );

    \I__7224\ : LocalMux
    port map (
            O => \N__36132\,
            I => \N__36097\
        );

    \I__7223\ : Span4Mux_s1_v
    port map (
            O => \N__36129\,
            I => \N__36094\
        );

    \I__7222\ : LocalMux
    port map (
            O => \N__36126\,
            I => \N__36087\
        );

    \I__7221\ : LocalMux
    port map (
            O => \N__36117\,
            I => \N__36087\
        );

    \I__7220\ : LocalMux
    port map (
            O => \N__36108\,
            I => \N__36087\
        );

    \I__7219\ : Span4Mux_h
    port map (
            O => \N__36097\,
            I => \N__36084\
        );

    \I__7218\ : Sp12to4
    port map (
            O => \N__36094\,
            I => \N__36081\
        );

    \I__7217\ : Span12Mux_h
    port map (
            O => \N__36087\,
            I => \N__36078\
        );

    \I__7216\ : Span4Mux_h
    port map (
            O => \N__36084\,
            I => \N__36075\
        );

    \I__7215\ : Span12Mux_s9_v
    port map (
            O => \N__36081\,
            I => \N__36072\
        );

    \I__7214\ : Odrv12
    port map (
            O => \N__36078\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__7213\ : Odrv4
    port map (
            O => \N__36075\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__7212\ : Odrv12
    port map (
            O => \N__36072\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__7211\ : InMux
    port map (
            O => \N__36065\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\
        );

    \I__7210\ : CascadeMux
    port map (
            O => \N__36062\,
            I => \N__36058\
        );

    \I__7209\ : InMux
    port map (
            O => \N__36061\,
            I => \N__36054\
        );

    \I__7208\ : InMux
    port map (
            O => \N__36058\,
            I => \N__36049\
        );

    \I__7207\ : InMux
    port map (
            O => \N__36057\,
            I => \N__36049\
        );

    \I__7206\ : LocalMux
    port map (
            O => \N__36054\,
            I => \N__36044\
        );

    \I__7205\ : LocalMux
    port map (
            O => \N__36049\,
            I => \N__36044\
        );

    \I__7204\ : Odrv4
    port map (
            O => \N__36044\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__7203\ : InMux
    port map (
            O => \N__36041\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\
        );

    \I__7202\ : InMux
    port map (
            O => \N__36038\,
            I => \bfn_14_13_0_\
        );

    \I__7201\ : InMux
    port map (
            O => \N__36035\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\
        );

    \I__7200\ : InMux
    port map (
            O => \N__36032\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\
        );

    \I__7199\ : InMux
    port map (
            O => \N__36029\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\
        );

    \I__7198\ : InMux
    port map (
            O => \N__36026\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__7197\ : CascadeMux
    port map (
            O => \N__36023\,
            I => \N__36018\
        );

    \I__7196\ : InMux
    port map (
            O => \N__36022\,
            I => \N__36015\
        );

    \I__7195\ : InMux
    port map (
            O => \N__36021\,
            I => \N__36010\
        );

    \I__7194\ : InMux
    port map (
            O => \N__36018\,
            I => \N__36010\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__36015\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__7192\ : LocalMux
    port map (
            O => \N__36010\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__7191\ : InMux
    port map (
            O => \N__36005\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\
        );

    \I__7190\ : CascadeMux
    port map (
            O => \N__36002\,
            I => \N__35997\
        );

    \I__7189\ : InMux
    port map (
            O => \N__36001\,
            I => \N__35994\
        );

    \I__7188\ : InMux
    port map (
            O => \N__36000\,
            I => \N__35989\
        );

    \I__7187\ : InMux
    port map (
            O => \N__35997\,
            I => \N__35989\
        );

    \I__7186\ : LocalMux
    port map (
            O => \N__35994\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__7185\ : LocalMux
    port map (
            O => \N__35989\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__7184\ : InMux
    port map (
            O => \N__35984\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\
        );

    \I__7183\ : CascadeMux
    port map (
            O => \N__35981\,
            I => \N__35977\
        );

    \I__7182\ : InMux
    port map (
            O => \N__35980\,
            I => \N__35973\
        );

    \I__7181\ : InMux
    port map (
            O => \N__35977\,
            I => \N__35968\
        );

    \I__7180\ : InMux
    port map (
            O => \N__35976\,
            I => \N__35968\
        );

    \I__7179\ : LocalMux
    port map (
            O => \N__35973\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__7178\ : LocalMux
    port map (
            O => \N__35968\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__7177\ : InMux
    port map (
            O => \N__35963\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\
        );

    \I__7176\ : InMux
    port map (
            O => \N__35960\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\
        );

    \I__7175\ : InMux
    port map (
            O => \N__35957\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\
        );

    \I__7174\ : InMux
    port map (
            O => \N__35954\,
            I => \bfn_14_12_0_\
        );

    \I__7173\ : InMux
    port map (
            O => \N__35951\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\
        );

    \I__7172\ : InMux
    port map (
            O => \N__35948\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\
        );

    \I__7171\ : InMux
    port map (
            O => \N__35945\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\
        );

    \I__7170\ : InMux
    port map (
            O => \N__35942\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\
        );

    \I__7169\ : InMux
    port map (
            O => \N__35939\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\
        );

    \I__7168\ : InMux
    port map (
            O => \N__35936\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\
        );

    \I__7167\ : InMux
    port map (
            O => \N__35933\,
            I => \N__35929\
        );

    \I__7166\ : InMux
    port map (
            O => \N__35932\,
            I => \N__35925\
        );

    \I__7165\ : LocalMux
    port map (
            O => \N__35929\,
            I => \N__35922\
        );

    \I__7164\ : InMux
    port map (
            O => \N__35928\,
            I => \N__35919\
        );

    \I__7163\ : LocalMux
    port map (
            O => \N__35925\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13\
        );

    \I__7162\ : Odrv4
    port map (
            O => \N__35922\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13\
        );

    \I__7161\ : LocalMux
    port map (
            O => \N__35919\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13\
        );

    \I__7160\ : InMux
    port map (
            O => \N__35912\,
            I => \N__35909\
        );

    \I__7159\ : LocalMux
    port map (
            O => \N__35909\,
            I => \N__35906\
        );

    \I__7158\ : Span4Mux_h
    port map (
            O => \N__35906\,
            I => \N__35903\
        );

    \I__7157\ : Odrv4
    port map (
            O => \N__35903\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\
        );

    \I__7156\ : InMux
    port map (
            O => \N__35900\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\
        );

    \I__7155\ : CascadeMux
    port map (
            O => \N__35897\,
            I => \N__35894\
        );

    \I__7154\ : InMux
    port map (
            O => \N__35894\,
            I => \N__35891\
        );

    \I__7153\ : LocalMux
    port map (
            O => \N__35891\,
            I => \N__35888\
        );

    \I__7152\ : Span4Mux_h
    port map (
            O => \N__35888\,
            I => \N__35885\
        );

    \I__7151\ : Odrv4
    port map (
            O => \N__35885\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1Z0Z_30\
        );

    \I__7150\ : InMux
    port map (
            O => \N__35882\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\
        );

    \I__7149\ : InMux
    port map (
            O => \N__35879\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\
        );

    \I__7148\ : InMux
    port map (
            O => \N__35876\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\
        );

    \I__7147\ : InMux
    port map (
            O => \N__35873\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\
        );

    \I__7146\ : IoInMux
    port map (
            O => \N__35870\,
            I => \N__35867\
        );

    \I__7145\ : LocalMux
    port map (
            O => \N__35867\,
            I => s2_phy_c
        );

    \I__7144\ : InMux
    port map (
            O => \N__35864\,
            I => \N__35861\
        );

    \I__7143\ : LocalMux
    port map (
            O => \N__35861\,
            I => \N__35857\
        );

    \I__7142\ : InMux
    port map (
            O => \N__35860\,
            I => \N__35854\
        );

    \I__7141\ : Span4Mux_v
    port map (
            O => \N__35857\,
            I => \N__35847\
        );

    \I__7140\ : LocalMux
    port map (
            O => \N__35854\,
            I => \N__35847\
        );

    \I__7139\ : InMux
    port map (
            O => \N__35853\,
            I => \N__35844\
        );

    \I__7138\ : InMux
    port map (
            O => \N__35852\,
            I => \N__35841\
        );

    \I__7137\ : Span4Mux_v
    port map (
            O => \N__35847\,
            I => \N__35838\
        );

    \I__7136\ : LocalMux
    port map (
            O => \N__35844\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__7135\ : LocalMux
    port map (
            O => \N__35841\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__7134\ : Odrv4
    port map (
            O => \N__35838\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__7133\ : InMux
    port map (
            O => \N__35831\,
            I => \N__35828\
        );

    \I__7132\ : LocalMux
    port map (
            O => \N__35828\,
            I => \N__35823\
        );

    \I__7131\ : InMux
    port map (
            O => \N__35827\,
            I => \N__35818\
        );

    \I__7130\ : InMux
    port map (
            O => \N__35826\,
            I => \N__35818\
        );

    \I__7129\ : Span4Mux_h
    port map (
            O => \N__35823\,
            I => \N__35812\
        );

    \I__7128\ : LocalMux
    port map (
            O => \N__35818\,
            I => \N__35812\
        );

    \I__7127\ : InMux
    port map (
            O => \N__35817\,
            I => \N__35809\
        );

    \I__7126\ : Span4Mux_v
    port map (
            O => \N__35812\,
            I => \N__35806\
        );

    \I__7125\ : LocalMux
    port map (
            O => \N__35809\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__7124\ : Odrv4
    port map (
            O => \N__35806\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__7123\ : InMux
    port map (
            O => \N__35801\,
            I => \N__35798\
        );

    \I__7122\ : LocalMux
    port map (
            O => \N__35798\,
            I => \N__35793\
        );

    \I__7121\ : InMux
    port map (
            O => \N__35797\,
            I => \N__35790\
        );

    \I__7120\ : InMux
    port map (
            O => \N__35796\,
            I => \N__35787\
        );

    \I__7119\ : Span4Mux_v
    port map (
            O => \N__35793\,
            I => \N__35782\
        );

    \I__7118\ : LocalMux
    port map (
            O => \N__35790\,
            I => \N__35782\
        );

    \I__7117\ : LocalMux
    port map (
            O => \N__35787\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__7116\ : Odrv4
    port map (
            O => \N__35782\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__7115\ : InMux
    port map (
            O => \N__35777\,
            I => \N__35774\
        );

    \I__7114\ : LocalMux
    port map (
            O => \N__35774\,
            I => \N__35770\
        );

    \I__7113\ : InMux
    port map (
            O => \N__35773\,
            I => \N__35766\
        );

    \I__7112\ : Span4Mux_v
    port map (
            O => \N__35770\,
            I => \N__35763\
        );

    \I__7111\ : InMux
    port map (
            O => \N__35769\,
            I => \N__35760\
        );

    \I__7110\ : LocalMux
    port map (
            O => \N__35766\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30\
        );

    \I__7109\ : Odrv4
    port map (
            O => \N__35763\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30\
        );

    \I__7108\ : LocalMux
    port map (
            O => \N__35760\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30\
        );

    \I__7107\ : InMux
    port map (
            O => \N__35753\,
            I => \N__35750\
        );

    \I__7106\ : LocalMux
    port map (
            O => \N__35750\,
            I => \current_shift_inst.un38_control_input_0_s0_24\
        );

    \I__7105\ : InMux
    port map (
            O => \N__35747\,
            I => \N__35744\
        );

    \I__7104\ : LocalMux
    port map (
            O => \N__35744\,
            I => \N__35741\
        );

    \I__7103\ : Span4Mux_v
    port map (
            O => \N__35741\,
            I => \N__35738\
        );

    \I__7102\ : Odrv4
    port map (
            O => \N__35738\,
            I => \current_shift_inst.control_input_axb_21\
        );

    \I__7101\ : InMux
    port map (
            O => \N__35735\,
            I => \N__35732\
        );

    \I__7100\ : LocalMux
    port map (
            O => \N__35732\,
            I => \current_shift_inst.un38_control_input_0_s0_25\
        );

    \I__7099\ : InMux
    port map (
            O => \N__35729\,
            I => \N__35726\
        );

    \I__7098\ : LocalMux
    port map (
            O => \N__35726\,
            I => \N__35723\
        );

    \I__7097\ : Span4Mux_h
    port map (
            O => \N__35723\,
            I => \N__35720\
        );

    \I__7096\ : Odrv4
    port map (
            O => \N__35720\,
            I => \current_shift_inst.control_input_axb_22\
        );

    \I__7095\ : CascadeMux
    port map (
            O => \N__35717\,
            I => \N__35714\
        );

    \I__7094\ : InMux
    port map (
            O => \N__35714\,
            I => \N__35711\
        );

    \I__7093\ : LocalMux
    port map (
            O => \N__35711\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\
        );

    \I__7092\ : InMux
    port map (
            O => \N__35708\,
            I => \N__35705\
        );

    \I__7091\ : LocalMux
    port map (
            O => \N__35705\,
            I => \current_shift_inst.un38_control_input_0_s0_26\
        );

    \I__7090\ : InMux
    port map (
            O => \N__35702\,
            I => \N__35699\
        );

    \I__7089\ : LocalMux
    port map (
            O => \N__35699\,
            I => \N__35696\
        );

    \I__7088\ : Span4Mux_h
    port map (
            O => \N__35696\,
            I => \N__35693\
        );

    \I__7087\ : Odrv4
    port map (
            O => \N__35693\,
            I => \current_shift_inst.control_input_axb_23\
        );

    \I__7086\ : CascadeMux
    port map (
            O => \N__35690\,
            I => \N__35687\
        );

    \I__7085\ : InMux
    port map (
            O => \N__35687\,
            I => \N__35684\
        );

    \I__7084\ : LocalMux
    port map (
            O => \N__35684\,
            I => \N__35681\
        );

    \I__7083\ : Span4Mux_h
    port map (
            O => \N__35681\,
            I => \N__35677\
        );

    \I__7082\ : InMux
    port map (
            O => \N__35680\,
            I => \N__35673\
        );

    \I__7081\ : Sp12to4
    port map (
            O => \N__35677\,
            I => \N__35670\
        );

    \I__7080\ : InMux
    port map (
            O => \N__35676\,
            I => \N__35667\
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__35673\,
            I => \N__35660\
        );

    \I__7078\ : Span12Mux_v
    port map (
            O => \N__35670\,
            I => \N__35660\
        );

    \I__7077\ : LocalMux
    port map (
            O => \N__35667\,
            I => \N__35660\
        );

    \I__7076\ : Span12Mux_v
    port map (
            O => \N__35660\,
            I => \N__35657\
        );

    \I__7075\ : Odrv12
    port map (
            O => \N__35657\,
            I => \il_max_comp1_D2\
        );

    \I__7074\ : IoInMux
    port map (
            O => \N__35654\,
            I => \N__35651\
        );

    \I__7073\ : LocalMux
    port map (
            O => \N__35651\,
            I => \N__35648\
        );

    \I__7072\ : Span4Mux_s3_v
    port map (
            O => \N__35648\,
            I => \N__35645\
        );

    \I__7071\ : Sp12to4
    port map (
            O => \N__35645\,
            I => \N__35642\
        );

    \I__7070\ : Span12Mux_h
    port map (
            O => \N__35642\,
            I => \N__35638\
        );

    \I__7069\ : InMux
    port map (
            O => \N__35641\,
            I => \N__35635\
        );

    \I__7068\ : Odrv12
    port map (
            O => \N__35638\,
            I => \T01_c\
        );

    \I__7067\ : LocalMux
    port map (
            O => \N__35635\,
            I => \T01_c\
        );

    \I__7066\ : CascadeMux
    port map (
            O => \N__35630\,
            I => \N__35625\
        );

    \I__7065\ : InMux
    port map (
            O => \N__35629\,
            I => \N__35618\
        );

    \I__7064\ : InMux
    port map (
            O => \N__35628\,
            I => \N__35618\
        );

    \I__7063\ : InMux
    port map (
            O => \N__35625\,
            I => \N__35615\
        );

    \I__7062\ : InMux
    port map (
            O => \N__35624\,
            I => \N__35610\
        );

    \I__7061\ : InMux
    port map (
            O => \N__35623\,
            I => \N__35610\
        );

    \I__7060\ : LocalMux
    port map (
            O => \N__35618\,
            I => \N__35603\
        );

    \I__7059\ : LocalMux
    port map (
            O => \N__35615\,
            I => \N__35603\
        );

    \I__7058\ : LocalMux
    port map (
            O => \N__35610\,
            I => \N__35603\
        );

    \I__7057\ : Span4Mux_v
    port map (
            O => \N__35603\,
            I => \N__35598\
        );

    \I__7056\ : InMux
    port map (
            O => \N__35602\,
            I => \N__35593\
        );

    \I__7055\ : InMux
    port map (
            O => \N__35601\,
            I => \N__35593\
        );

    \I__7054\ : Odrv4
    port map (
            O => \N__35598\,
            I => state_3
        );

    \I__7053\ : LocalMux
    port map (
            O => \N__35593\,
            I => state_3
        );

    \I__7052\ : IoInMux
    port map (
            O => \N__35588\,
            I => \N__35585\
        );

    \I__7051\ : LocalMux
    port map (
            O => \N__35585\,
            I => \N__35582\
        );

    \I__7050\ : Span4Mux_s2_v
    port map (
            O => \N__35582\,
            I => \N__35579\
        );

    \I__7049\ : Span4Mux_h
    port map (
            O => \N__35579\,
            I => \N__35576\
        );

    \I__7048\ : Span4Mux_v
    port map (
            O => \N__35576\,
            I => \N__35571\
        );

    \I__7047\ : InMux
    port map (
            O => \N__35575\,
            I => \N__35568\
        );

    \I__7046\ : InMux
    port map (
            O => \N__35574\,
            I => \N__35565\
        );

    \I__7045\ : Odrv4
    port map (
            O => \N__35571\,
            I => s1_phy_c
        );

    \I__7044\ : LocalMux
    port map (
            O => \N__35568\,
            I => s1_phy_c
        );

    \I__7043\ : LocalMux
    port map (
            O => \N__35565\,
            I => s1_phy_c
        );

    \I__7042\ : IoInMux
    port map (
            O => \N__35558\,
            I => \N__35555\
        );

    \I__7041\ : LocalMux
    port map (
            O => \N__35555\,
            I => \N__35552\
        );

    \I__7040\ : Span12Mux_s0_v
    port map (
            O => \N__35552\,
            I => \N__35549\
        );

    \I__7039\ : Odrv12
    port map (
            O => \N__35549\,
            I => \current_shift_inst.timer_s1.N_162_i\
        );

    \I__7038\ : InMux
    port map (
            O => \N__35546\,
            I => \N__35543\
        );

    \I__7037\ : LocalMux
    port map (
            O => \N__35543\,
            I => \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\
        );

    \I__7036\ : InMux
    port map (
            O => \N__35540\,
            I => \N__35537\
        );

    \I__7035\ : LocalMux
    port map (
            O => \N__35537\,
            I => \current_shift_inst.un38_control_input_0_s0_27\
        );

    \I__7034\ : InMux
    port map (
            O => \N__35534\,
            I => \N__35531\
        );

    \I__7033\ : LocalMux
    port map (
            O => \N__35531\,
            I => \N__35528\
        );

    \I__7032\ : Odrv4
    port map (
            O => \N__35528\,
            I => \current_shift_inst.control_input_axb_24\
        );

    \I__7031\ : InMux
    port map (
            O => \N__35525\,
            I => \N__35522\
        );

    \I__7030\ : LocalMux
    port map (
            O => \N__35522\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\
        );

    \I__7029\ : CascadeMux
    port map (
            O => \N__35519\,
            I => \N__35516\
        );

    \I__7028\ : InMux
    port map (
            O => \N__35516\,
            I => \N__35513\
        );

    \I__7027\ : LocalMux
    port map (
            O => \N__35513\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\
        );

    \I__7026\ : CascadeMux
    port map (
            O => \N__35510\,
            I => \N__35507\
        );

    \I__7025\ : InMux
    port map (
            O => \N__35507\,
            I => \N__35504\
        );

    \I__7024\ : LocalMux
    port map (
            O => \N__35504\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\
        );

    \I__7023\ : InMux
    port map (
            O => \N__35501\,
            I => \N__35498\
        );

    \I__7022\ : LocalMux
    port map (
            O => \N__35498\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\
        );

    \I__7021\ : CascadeMux
    port map (
            O => \N__35495\,
            I => \N__35492\
        );

    \I__7020\ : InMux
    port map (
            O => \N__35492\,
            I => \N__35489\
        );

    \I__7019\ : LocalMux
    port map (
            O => \N__35489\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\
        );

    \I__7018\ : InMux
    port map (
            O => \N__35486\,
            I => \N__35483\
        );

    \I__7017\ : LocalMux
    port map (
            O => \N__35483\,
            I => \current_shift_inst.un38_control_input_0_s0_29\
        );

    \I__7016\ : InMux
    port map (
            O => \N__35480\,
            I => \N__35477\
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__35477\,
            I => \N__35474\
        );

    \I__7014\ : Span4Mux_v
    port map (
            O => \N__35474\,
            I => \N__35471\
        );

    \I__7013\ : Odrv4
    port map (
            O => \N__35471\,
            I => \current_shift_inst.control_input_axb_26\
        );

    \I__7012\ : InMux
    port map (
            O => \N__35468\,
            I => \N__35465\
        );

    \I__7011\ : LocalMux
    port map (
            O => \N__35465\,
            I => \current_shift_inst.un38_control_input_0_s0_23\
        );

    \I__7010\ : InMux
    port map (
            O => \N__35462\,
            I => \N__35459\
        );

    \I__7009\ : LocalMux
    port map (
            O => \N__35459\,
            I => \N__35456\
        );

    \I__7008\ : Span4Mux_v
    port map (
            O => \N__35456\,
            I => \N__35453\
        );

    \I__7007\ : Odrv4
    port map (
            O => \N__35453\,
            I => \current_shift_inst.control_input_axb_20\
        );

    \I__7006\ : CascadeMux
    port map (
            O => \N__35450\,
            I => \N__35447\
        );

    \I__7005\ : InMux
    port map (
            O => \N__35447\,
            I => \N__35444\
        );

    \I__7004\ : LocalMux
    port map (
            O => \N__35444\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\
        );

    \I__7003\ : CascadeMux
    port map (
            O => \N__35441\,
            I => \N__35438\
        );

    \I__7002\ : InMux
    port map (
            O => \N__35438\,
            I => \N__35435\
        );

    \I__7001\ : LocalMux
    port map (
            O => \N__35435\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\
        );

    \I__7000\ : CascadeMux
    port map (
            O => \N__35432\,
            I => \N__35429\
        );

    \I__6999\ : InMux
    port map (
            O => \N__35429\,
            I => \N__35426\
        );

    \I__6998\ : LocalMux
    port map (
            O => \N__35426\,
            I => \N__35423\
        );

    \I__6997\ : Odrv12
    port map (
            O => \N__35423\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\
        );

    \I__6996\ : CascadeMux
    port map (
            O => \N__35420\,
            I => \N__35417\
        );

    \I__6995\ : InMux
    port map (
            O => \N__35417\,
            I => \N__35414\
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__35414\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\
        );

    \I__6993\ : InMux
    port map (
            O => \N__35411\,
            I => \N__35408\
        );

    \I__6992\ : LocalMux
    port map (
            O => \N__35408\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\
        );

    \I__6991\ : InMux
    port map (
            O => \N__35405\,
            I => \N__35402\
        );

    \I__6990\ : LocalMux
    port map (
            O => \N__35402\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\
        );

    \I__6989\ : InMux
    port map (
            O => \N__35399\,
            I => \N__35396\
        );

    \I__6988\ : LocalMux
    port map (
            O => \N__35396\,
            I => \current_shift_inst.un38_control_input_0_s0_19\
        );

    \I__6987\ : InMux
    port map (
            O => \N__35393\,
            I => \N__35390\
        );

    \I__6986\ : LocalMux
    port map (
            O => \N__35390\,
            I => \N__35387\
        );

    \I__6985\ : Odrv4
    port map (
            O => \N__35387\,
            I => \current_shift_inst.control_input_axb_16\
        );

    \I__6984\ : InMux
    port map (
            O => \N__35384\,
            I => \N__35381\
        );

    \I__6983\ : LocalMux
    port map (
            O => \N__35381\,
            I => \current_shift_inst.un38_control_input_0_s0_28\
        );

    \I__6982\ : InMux
    port map (
            O => \N__35378\,
            I => \N__35375\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__35375\,
            I => \N__35372\
        );

    \I__6980\ : Odrv4
    port map (
            O => \N__35372\,
            I => \current_shift_inst.control_input_axb_25\
        );

    \I__6979\ : InMux
    port map (
            O => \N__35369\,
            I => \N__35366\
        );

    \I__6978\ : LocalMux
    port map (
            O => \N__35366\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6\
        );

    \I__6977\ : InMux
    port map (
            O => \N__35363\,
            I => \N__35360\
        );

    \I__6976\ : LocalMux
    port map (
            O => \N__35360\,
            I => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\
        );

    \I__6975\ : CascadeMux
    port map (
            O => \N__35357\,
            I => \N__35354\
        );

    \I__6974\ : InMux
    port map (
            O => \N__35354\,
            I => \N__35351\
        );

    \I__6973\ : LocalMux
    port map (
            O => \N__35351\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\
        );

    \I__6972\ : CascadeMux
    port map (
            O => \N__35348\,
            I => \N__35345\
        );

    \I__6971\ : InMux
    port map (
            O => \N__35345\,
            I => \N__35342\
        );

    \I__6970\ : LocalMux
    port map (
            O => \N__35342\,
            I => \current_shift_inst.un38_control_input_0_s0_14\
        );

    \I__6969\ : CascadeMux
    port map (
            O => \N__35339\,
            I => \N__35336\
        );

    \I__6968\ : InMux
    port map (
            O => \N__35336\,
            I => \N__35333\
        );

    \I__6967\ : LocalMux
    port map (
            O => \N__35333\,
            I => \N__35330\
        );

    \I__6966\ : Odrv4
    port map (
            O => \N__35330\,
            I => \current_shift_inst.control_input_axb_11\
        );

    \I__6965\ : InMux
    port map (
            O => \N__35327\,
            I => \N__35324\
        );

    \I__6964\ : LocalMux
    port map (
            O => \N__35324\,
            I => \current_shift_inst.un38_control_input_0_s0_15\
        );

    \I__6963\ : InMux
    port map (
            O => \N__35321\,
            I => \N__35318\
        );

    \I__6962\ : LocalMux
    port map (
            O => \N__35318\,
            I => \N__35315\
        );

    \I__6961\ : Odrv4
    port map (
            O => \N__35315\,
            I => \current_shift_inst.control_input_axb_12\
        );

    \I__6960\ : InMux
    port map (
            O => \N__35312\,
            I => \N__35309\
        );

    \I__6959\ : LocalMux
    port map (
            O => \N__35309\,
            I => \N__35306\
        );

    \I__6958\ : Odrv4
    port map (
            O => \N__35306\,
            I => \current_shift_inst.un38_control_input_0_s0_16\
        );

    \I__6957\ : InMux
    port map (
            O => \N__35303\,
            I => \N__35300\
        );

    \I__6956\ : LocalMux
    port map (
            O => \N__35300\,
            I => \N__35297\
        );

    \I__6955\ : Odrv4
    port map (
            O => \N__35297\,
            I => \current_shift_inst.control_input_axb_13\
        );

    \I__6954\ : InMux
    port map (
            O => \N__35294\,
            I => \N__35291\
        );

    \I__6953\ : LocalMux
    port map (
            O => \N__35291\,
            I => \N__35288\
        );

    \I__6952\ : Odrv4
    port map (
            O => \N__35288\,
            I => \current_shift_inst.un38_control_input_0_s0_17\
        );

    \I__6951\ : InMux
    port map (
            O => \N__35285\,
            I => \N__35282\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__35282\,
            I => \N__35279\
        );

    \I__6949\ : Odrv4
    port map (
            O => \N__35279\,
            I => \current_shift_inst.control_input_axb_14\
        );

    \I__6948\ : InMux
    port map (
            O => \N__35276\,
            I => \N__35273\
        );

    \I__6947\ : LocalMux
    port map (
            O => \N__35273\,
            I => \N__35270\
        );

    \I__6946\ : Odrv4
    port map (
            O => \N__35270\,
            I => \current_shift_inst.un38_control_input_0_s0_18\
        );

    \I__6945\ : InMux
    port map (
            O => \N__35267\,
            I => \N__35264\
        );

    \I__6944\ : LocalMux
    port map (
            O => \N__35264\,
            I => \N__35261\
        );

    \I__6943\ : Odrv4
    port map (
            O => \N__35261\,
            I => \current_shift_inst.control_input_axb_15\
        );

    \I__6942\ : InMux
    port map (
            O => \N__35258\,
            I => \N__35255\
        );

    \I__6941\ : LocalMux
    port map (
            O => \N__35255\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\
        );

    \I__6940\ : InMux
    port map (
            O => \N__35252\,
            I => \N__35246\
        );

    \I__6939\ : InMux
    port map (
            O => \N__35251\,
            I => \N__35246\
        );

    \I__6938\ : LocalMux
    port map (
            O => \N__35246\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_24\
        );

    \I__6937\ : CascadeMux
    port map (
            O => \N__35243\,
            I => \N__35240\
        );

    \I__6936\ : InMux
    port map (
            O => \N__35240\,
            I => \N__35234\
        );

    \I__6935\ : InMux
    port map (
            O => \N__35239\,
            I => \N__35234\
        );

    \I__6934\ : LocalMux
    port map (
            O => \N__35234\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_25\
        );

    \I__6933\ : CascadeMux
    port map (
            O => \N__35231\,
            I => \N__35228\
        );

    \I__6932\ : InMux
    port map (
            O => \N__35228\,
            I => \N__35222\
        );

    \I__6931\ : InMux
    port map (
            O => \N__35227\,
            I => \N__35222\
        );

    \I__6930\ : LocalMux
    port map (
            O => \N__35222\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\
        );

    \I__6929\ : InMux
    port map (
            O => \N__35219\,
            I => \N__35213\
        );

    \I__6928\ : InMux
    port map (
            O => \N__35218\,
            I => \N__35213\
        );

    \I__6927\ : LocalMux
    port map (
            O => \N__35213\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_30\
        );

    \I__6926\ : InMux
    port map (
            O => \N__35210\,
            I => \N__35207\
        );

    \I__6925\ : LocalMux
    port map (
            O => \N__35207\,
            I => \N__35204\
        );

    \I__6924\ : Odrv4
    port map (
            O => \N__35204\,
            I => \current_shift_inst.un38_control_input_0_s0_10\
        );

    \I__6923\ : InMux
    port map (
            O => \N__35201\,
            I => \N__35198\
        );

    \I__6922\ : LocalMux
    port map (
            O => \N__35198\,
            I => \N__35195\
        );

    \I__6921\ : Odrv4
    port map (
            O => \N__35195\,
            I => \current_shift_inst.control_input_axb_7\
        );

    \I__6920\ : CascadeMux
    port map (
            O => \N__35192\,
            I => \N__35189\
        );

    \I__6919\ : InMux
    port map (
            O => \N__35189\,
            I => \N__35186\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__35186\,
            I => \N__35183\
        );

    \I__6917\ : Odrv4
    port map (
            O => \N__35183\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\
        );

    \I__6916\ : InMux
    port map (
            O => \N__35180\,
            I => \N__35174\
        );

    \I__6915\ : InMux
    port map (
            O => \N__35179\,
            I => \N__35174\
        );

    \I__6914\ : LocalMux
    port map (
            O => \N__35174\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_23\
        );

    \I__6913\ : CascadeMux
    port map (
            O => \N__35171\,
            I => \N__35165\
        );

    \I__6912\ : InMux
    port map (
            O => \N__35170\,
            I => \N__35161\
        );

    \I__6911\ : InMux
    port map (
            O => \N__35169\,
            I => \N__35158\
        );

    \I__6910\ : InMux
    port map (
            O => \N__35168\,
            I => \N__35155\
        );

    \I__6909\ : InMux
    port map (
            O => \N__35165\,
            I => \N__35152\
        );

    \I__6908\ : InMux
    port map (
            O => \N__35164\,
            I => \N__35149\
        );

    \I__6907\ : LocalMux
    port map (
            O => \N__35161\,
            I => \N__35146\
        );

    \I__6906\ : LocalMux
    port map (
            O => \N__35158\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__6905\ : LocalMux
    port map (
            O => \N__35155\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__6904\ : LocalMux
    port map (
            O => \N__35152\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__6903\ : LocalMux
    port map (
            O => \N__35149\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__6902\ : Odrv12
    port map (
            O => \N__35146\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__6901\ : InMux
    port map (
            O => \N__35135\,
            I => \N__35131\
        );

    \I__6900\ : InMux
    port map (
            O => \N__35134\,
            I => \N__35128\
        );

    \I__6899\ : LocalMux
    port map (
            O => \N__35131\,
            I => \N__35124\
        );

    \I__6898\ : LocalMux
    port map (
            O => \N__35128\,
            I => \N__35121\
        );

    \I__6897\ : InMux
    port map (
            O => \N__35127\,
            I => \N__35118\
        );

    \I__6896\ : Span4Mux_h
    port map (
            O => \N__35124\,
            I => \N__35111\
        );

    \I__6895\ : Span4Mux_v
    port map (
            O => \N__35121\,
            I => \N__35111\
        );

    \I__6894\ : LocalMux
    port map (
            O => \N__35118\,
            I => \N__35111\
        );

    \I__6893\ : Odrv4
    port map (
            O => \N__35111\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__6892\ : InMux
    port map (
            O => \N__35108\,
            I => \N__35104\
        );

    \I__6891\ : InMux
    port map (
            O => \N__35107\,
            I => \N__35101\
        );

    \I__6890\ : LocalMux
    port map (
            O => \N__35104\,
            I => \phase_controller_inst1.stoper_tr.runningZ0\
        );

    \I__6889\ : LocalMux
    port map (
            O => \N__35101\,
            I => \phase_controller_inst1.stoper_tr.runningZ0\
        );

    \I__6888\ : InMux
    port map (
            O => \N__35096\,
            I => \N__35093\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__35093\,
            I => \N__35088\
        );

    \I__6886\ : InMux
    port map (
            O => \N__35092\,
            I => \N__35083\
        );

    \I__6885\ : InMux
    port map (
            O => \N__35091\,
            I => \N__35083\
        );

    \I__6884\ : Odrv4
    port map (
            O => \N__35088\,
            I => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\
        );

    \I__6883\ : LocalMux
    port map (
            O => \N__35083\,
            I => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\
        );

    \I__6882\ : CascadeMux
    port map (
            O => \N__35078\,
            I => \N__35075\
        );

    \I__6881\ : InMux
    port map (
            O => \N__35075\,
            I => \N__35071\
        );

    \I__6880\ : InMux
    port map (
            O => \N__35074\,
            I => \N__35068\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__35071\,
            I => \N__35061\
        );

    \I__6878\ : LocalMux
    port map (
            O => \N__35068\,
            I => \N__35061\
        );

    \I__6877\ : InMux
    port map (
            O => \N__35067\,
            I => \N__35056\
        );

    \I__6876\ : InMux
    port map (
            O => \N__35066\,
            I => \N__35056\
        );

    \I__6875\ : Odrv12
    port map (
            O => \N__35061\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__6874\ : LocalMux
    port map (
            O => \N__35056\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__6873\ : InMux
    port map (
            O => \N__35051\,
            I => \N__35048\
        );

    \I__6872\ : LocalMux
    port map (
            O => \N__35048\,
            I => \phase_controller_inst1.state_RNI7NN7Z0Z_0\
        );

    \I__6871\ : InMux
    port map (
            O => \N__35045\,
            I => \N__35042\
        );

    \I__6870\ : LocalMux
    port map (
            O => \N__35042\,
            I => \phase_controller_inst1.start_timer_tr_RNOZ0Z_0\
        );

    \I__6869\ : InMux
    port map (
            O => \N__35039\,
            I => \N__35031\
        );

    \I__6868\ : InMux
    port map (
            O => \N__35038\,
            I => \N__35031\
        );

    \I__6867\ : InMux
    port map (
            O => \N__35037\,
            I => \N__35026\
        );

    \I__6866\ : InMux
    port map (
            O => \N__35036\,
            I => \N__35026\
        );

    \I__6865\ : LocalMux
    port map (
            O => \N__35031\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__6864\ : LocalMux
    port map (
            O => \N__35026\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__6863\ : CascadeMux
    port map (
            O => \N__35021\,
            I => \N__35017\
        );

    \I__6862\ : CascadeMux
    port map (
            O => \N__35020\,
            I => \N__35014\
        );

    \I__6861\ : InMux
    port map (
            O => \N__35017\,
            I => \N__35008\
        );

    \I__6860\ : InMux
    port map (
            O => \N__35014\,
            I => \N__35005\
        );

    \I__6859\ : InMux
    port map (
            O => \N__35013\,
            I => \N__35000\
        );

    \I__6858\ : InMux
    port map (
            O => \N__35012\,
            I => \N__35000\
        );

    \I__6857\ : InMux
    port map (
            O => \N__35011\,
            I => \N__34997\
        );

    \I__6856\ : LocalMux
    port map (
            O => \N__35008\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__6855\ : LocalMux
    port map (
            O => \N__35005\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__6854\ : LocalMux
    port map (
            O => \N__35000\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__6853\ : LocalMux
    port map (
            O => \N__34997\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__6852\ : InMux
    port map (
            O => \N__34988\,
            I => \N__34983\
        );

    \I__6851\ : InMux
    port map (
            O => \N__34987\,
            I => \N__34980\
        );

    \I__6850\ : InMux
    port map (
            O => \N__34986\,
            I => \N__34977\
        );

    \I__6849\ : LocalMux
    port map (
            O => \N__34983\,
            I => \N__34974\
        );

    \I__6848\ : LocalMux
    port map (
            O => \N__34980\,
            I => \N__34969\
        );

    \I__6847\ : LocalMux
    port map (
            O => \N__34977\,
            I => \N__34969\
        );

    \I__6846\ : Sp12to4
    port map (
            O => \N__34974\,
            I => \N__34964\
        );

    \I__6845\ : Sp12to4
    port map (
            O => \N__34969\,
            I => \N__34964\
        );

    \I__6844\ : Span12Mux_v
    port map (
            O => \N__34964\,
            I => \N__34961\
        );

    \I__6843\ : Odrv12
    port map (
            O => \N__34961\,
            I => \il_min_comp1_D2\
        );

    \I__6842\ : CascadeMux
    port map (
            O => \N__34958\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24_cascade_\
        );

    \I__6841\ : InMux
    port map (
            O => \N__34955\,
            I => \N__34949\
        );

    \I__6840\ : InMux
    port map (
            O => \N__34954\,
            I => \N__34949\
        );

    \I__6839\ : LocalMux
    port map (
            O => \N__34949\,
            I => \N__34945\
        );

    \I__6838\ : InMux
    port map (
            O => \N__34948\,
            I => \N__34942\
        );

    \I__6837\ : Span4Mux_h
    port map (
            O => \N__34945\,
            I => \N__34939\
        );

    \I__6836\ : LocalMux
    port map (
            O => \N__34942\,
            I => \N__34935\
        );

    \I__6835\ : Span4Mux_h
    port map (
            O => \N__34939\,
            I => \N__34932\
        );

    \I__6834\ : InMux
    port map (
            O => \N__34938\,
            I => \N__34929\
        );

    \I__6833\ : Odrv4
    port map (
            O => \N__34935\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__6832\ : Odrv4
    port map (
            O => \N__34932\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__6831\ : LocalMux
    port map (
            O => \N__34929\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__6830\ : InMux
    port map (
            O => \N__34922\,
            I => \N__34916\
        );

    \I__6829\ : InMux
    port map (
            O => \N__34921\,
            I => \N__34916\
        );

    \I__6828\ : LocalMux
    port map (
            O => \N__34916\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_24\
        );

    \I__6827\ : InMux
    port map (
            O => \N__34913\,
            I => \N__34910\
        );

    \I__6826\ : LocalMux
    port map (
            O => \N__34910\,
            I => \N__34906\
        );

    \I__6825\ : InMux
    port map (
            O => \N__34909\,
            I => \N__34902\
        );

    \I__6824\ : Span4Mux_h
    port map (
            O => \N__34906\,
            I => \N__34899\
        );

    \I__6823\ : InMux
    port map (
            O => \N__34905\,
            I => \N__34896\
        );

    \I__6822\ : LocalMux
    port map (
            O => \N__34902\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7\
        );

    \I__6821\ : Odrv4
    port map (
            O => \N__34899\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7\
        );

    \I__6820\ : LocalMux
    port map (
            O => \N__34896\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7\
        );

    \I__6819\ : InMux
    port map (
            O => \N__34889\,
            I => \N__34886\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__34886\,
            I => \N__34882\
        );

    \I__6817\ : InMux
    port map (
            O => \N__34885\,
            I => \N__34878\
        );

    \I__6816\ : Span4Mux_v
    port map (
            O => \N__34882\,
            I => \N__34875\
        );

    \I__6815\ : InMux
    port map (
            O => \N__34881\,
            I => \N__34872\
        );

    \I__6814\ : LocalMux
    port map (
            O => \N__34878\,
            I => \N__34868\
        );

    \I__6813\ : Sp12to4
    port map (
            O => \N__34875\,
            I => \N__34863\
        );

    \I__6812\ : LocalMux
    port map (
            O => \N__34872\,
            I => \N__34863\
        );

    \I__6811\ : InMux
    port map (
            O => \N__34871\,
            I => \N__34860\
        );

    \I__6810\ : Odrv4
    port map (
            O => \N__34868\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__6809\ : Odrv12
    port map (
            O => \N__34863\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__6808\ : LocalMux
    port map (
            O => \N__34860\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__6807\ : InMux
    port map (
            O => \N__34853\,
            I => \N__34850\
        );

    \I__6806\ : LocalMux
    port map (
            O => \N__34850\,
            I => \N__34847\
        );

    \I__6805\ : Odrv12
    port map (
            O => \N__34847\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\
        );

    \I__6804\ : InMux
    port map (
            O => \N__34844\,
            I => \N__34825\
        );

    \I__6803\ : InMux
    port map (
            O => \N__34843\,
            I => \N__34818\
        );

    \I__6802\ : InMux
    port map (
            O => \N__34842\,
            I => \N__34818\
        );

    \I__6801\ : InMux
    port map (
            O => \N__34841\,
            I => \N__34818\
        );

    \I__6800\ : InMux
    port map (
            O => \N__34840\,
            I => \N__34810\
        );

    \I__6799\ : InMux
    port map (
            O => \N__34839\,
            I => \N__34810\
        );

    \I__6798\ : InMux
    port map (
            O => \N__34838\,
            I => \N__34795\
        );

    \I__6797\ : InMux
    port map (
            O => \N__34837\,
            I => \N__34795\
        );

    \I__6796\ : InMux
    port map (
            O => \N__34836\,
            I => \N__34795\
        );

    \I__6795\ : InMux
    port map (
            O => \N__34835\,
            I => \N__34795\
        );

    \I__6794\ : InMux
    port map (
            O => \N__34834\,
            I => \N__34795\
        );

    \I__6793\ : InMux
    port map (
            O => \N__34833\,
            I => \N__34795\
        );

    \I__6792\ : InMux
    port map (
            O => \N__34832\,
            I => \N__34795\
        );

    \I__6791\ : InMux
    port map (
            O => \N__34831\,
            I => \N__34786\
        );

    \I__6790\ : InMux
    port map (
            O => \N__34830\,
            I => \N__34786\
        );

    \I__6789\ : InMux
    port map (
            O => \N__34829\,
            I => \N__34786\
        );

    \I__6788\ : InMux
    port map (
            O => \N__34828\,
            I => \N__34786\
        );

    \I__6787\ : LocalMux
    port map (
            O => \N__34825\,
            I => \N__34781\
        );

    \I__6786\ : LocalMux
    port map (
            O => \N__34818\,
            I => \N__34781\
        );

    \I__6785\ : InMux
    port map (
            O => \N__34817\,
            I => \N__34762\
        );

    \I__6784\ : InMux
    port map (
            O => \N__34816\,
            I => \N__34759\
        );

    \I__6783\ : InMux
    port map (
            O => \N__34815\,
            I => \N__34743\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__34810\,
            I => \N__34723\
        );

    \I__6781\ : LocalMux
    port map (
            O => \N__34795\,
            I => \N__34723\
        );

    \I__6780\ : LocalMux
    port map (
            O => \N__34786\,
            I => \N__34723\
        );

    \I__6779\ : Span4Mux_v
    port map (
            O => \N__34781\,
            I => \N__34723\
        );

    \I__6778\ : InMux
    port map (
            O => \N__34780\,
            I => \N__34712\
        );

    \I__6777\ : InMux
    port map (
            O => \N__34779\,
            I => \N__34712\
        );

    \I__6776\ : InMux
    port map (
            O => \N__34778\,
            I => \N__34712\
        );

    \I__6775\ : InMux
    port map (
            O => \N__34777\,
            I => \N__34712\
        );

    \I__6774\ : InMux
    port map (
            O => \N__34776\,
            I => \N__34712\
        );

    \I__6773\ : InMux
    port map (
            O => \N__34775\,
            I => \N__34704\
        );

    \I__6772\ : InMux
    port map (
            O => \N__34774\,
            I => \N__34704\
        );

    \I__6771\ : InMux
    port map (
            O => \N__34773\,
            I => \N__34691\
        );

    \I__6770\ : InMux
    port map (
            O => \N__34772\,
            I => \N__34691\
        );

    \I__6769\ : InMux
    port map (
            O => \N__34771\,
            I => \N__34691\
        );

    \I__6768\ : InMux
    port map (
            O => \N__34770\,
            I => \N__34691\
        );

    \I__6767\ : InMux
    port map (
            O => \N__34769\,
            I => \N__34691\
        );

    \I__6766\ : InMux
    port map (
            O => \N__34768\,
            I => \N__34691\
        );

    \I__6765\ : InMux
    port map (
            O => \N__34767\,
            I => \N__34686\
        );

    \I__6764\ : InMux
    port map (
            O => \N__34766\,
            I => \N__34686\
        );

    \I__6763\ : CascadeMux
    port map (
            O => \N__34765\,
            I => \N__34680\
        );

    \I__6762\ : LocalMux
    port map (
            O => \N__34762\,
            I => \N__34674\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__34759\,
            I => \N__34674\
        );

    \I__6760\ : InMux
    port map (
            O => \N__34758\,
            I => \N__34663\
        );

    \I__6759\ : InMux
    port map (
            O => \N__34757\,
            I => \N__34660\
        );

    \I__6758\ : InMux
    port map (
            O => \N__34756\,
            I => \N__34647\
        );

    \I__6757\ : InMux
    port map (
            O => \N__34755\,
            I => \N__34647\
        );

    \I__6756\ : InMux
    port map (
            O => \N__34754\,
            I => \N__34647\
        );

    \I__6755\ : InMux
    port map (
            O => \N__34753\,
            I => \N__34647\
        );

    \I__6754\ : InMux
    port map (
            O => \N__34752\,
            I => \N__34647\
        );

    \I__6753\ : InMux
    port map (
            O => \N__34751\,
            I => \N__34647\
        );

    \I__6752\ : InMux
    port map (
            O => \N__34750\,
            I => \N__34636\
        );

    \I__6751\ : InMux
    port map (
            O => \N__34749\,
            I => \N__34636\
        );

    \I__6750\ : InMux
    port map (
            O => \N__34748\,
            I => \N__34636\
        );

    \I__6749\ : InMux
    port map (
            O => \N__34747\,
            I => \N__34636\
        );

    \I__6748\ : InMux
    port map (
            O => \N__34746\,
            I => \N__34636\
        );

    \I__6747\ : LocalMux
    port map (
            O => \N__34743\,
            I => \N__34633\
        );

    \I__6746\ : InMux
    port map (
            O => \N__34742\,
            I => \N__34630\
        );

    \I__6745\ : InMux
    port map (
            O => \N__34741\,
            I => \N__34623\
        );

    \I__6744\ : InMux
    port map (
            O => \N__34740\,
            I => \N__34623\
        );

    \I__6743\ : InMux
    port map (
            O => \N__34739\,
            I => \N__34623\
        );

    \I__6742\ : InMux
    port map (
            O => \N__34738\,
            I => \N__34620\
        );

    \I__6741\ : InMux
    port map (
            O => \N__34737\,
            I => \N__34615\
        );

    \I__6740\ : InMux
    port map (
            O => \N__34736\,
            I => \N__34615\
        );

    \I__6739\ : InMux
    port map (
            O => \N__34735\,
            I => \N__34590\
        );

    \I__6738\ : InMux
    port map (
            O => \N__34734\,
            I => \N__34590\
        );

    \I__6737\ : InMux
    port map (
            O => \N__34733\,
            I => \N__34590\
        );

    \I__6736\ : InMux
    port map (
            O => \N__34732\,
            I => \N__34590\
        );

    \I__6735\ : Span4Mux_v
    port map (
            O => \N__34723\,
            I => \N__34585\
        );

    \I__6734\ : LocalMux
    port map (
            O => \N__34712\,
            I => \N__34585\
        );

    \I__6733\ : CascadeMux
    port map (
            O => \N__34711\,
            I => \N__34582\
        );

    \I__6732\ : InMux
    port map (
            O => \N__34710\,
            I => \N__34578\
        );

    \I__6731\ : InMux
    port map (
            O => \N__34709\,
            I => \N__34575\
        );

    \I__6730\ : LocalMux
    port map (
            O => \N__34704\,
            I => \N__34568\
        );

    \I__6729\ : LocalMux
    port map (
            O => \N__34691\,
            I => \N__34568\
        );

    \I__6728\ : LocalMux
    port map (
            O => \N__34686\,
            I => \N__34568\
        );

    \I__6727\ : InMux
    port map (
            O => \N__34685\,
            I => \N__34557\
        );

    \I__6726\ : InMux
    port map (
            O => \N__34684\,
            I => \N__34557\
        );

    \I__6725\ : InMux
    port map (
            O => \N__34683\,
            I => \N__34557\
        );

    \I__6724\ : InMux
    port map (
            O => \N__34680\,
            I => \N__34557\
        );

    \I__6723\ : InMux
    port map (
            O => \N__34679\,
            I => \N__34557\
        );

    \I__6722\ : Span4Mux_v
    port map (
            O => \N__34674\,
            I => \N__34554\
        );

    \I__6721\ : InMux
    port map (
            O => \N__34673\,
            I => \N__34551\
        );

    \I__6720\ : InMux
    port map (
            O => \N__34672\,
            I => \N__34536\
        );

    \I__6719\ : InMux
    port map (
            O => \N__34671\,
            I => \N__34536\
        );

    \I__6718\ : InMux
    port map (
            O => \N__34670\,
            I => \N__34536\
        );

    \I__6717\ : InMux
    port map (
            O => \N__34669\,
            I => \N__34536\
        );

    \I__6716\ : InMux
    port map (
            O => \N__34668\,
            I => \N__34536\
        );

    \I__6715\ : InMux
    port map (
            O => \N__34667\,
            I => \N__34536\
        );

    \I__6714\ : InMux
    port map (
            O => \N__34666\,
            I => \N__34536\
        );

    \I__6713\ : LocalMux
    port map (
            O => \N__34663\,
            I => \N__34533\
        );

    \I__6712\ : LocalMux
    port map (
            O => \N__34660\,
            I => \N__34530\
        );

    \I__6711\ : LocalMux
    port map (
            O => \N__34647\,
            I => \N__34525\
        );

    \I__6710\ : LocalMux
    port map (
            O => \N__34636\,
            I => \N__34525\
        );

    \I__6709\ : Span4Mux_v
    port map (
            O => \N__34633\,
            I => \N__34520\
        );

    \I__6708\ : LocalMux
    port map (
            O => \N__34630\,
            I => \N__34520\
        );

    \I__6707\ : LocalMux
    port map (
            O => \N__34623\,
            I => \N__34517\
        );

    \I__6706\ : LocalMux
    port map (
            O => \N__34620\,
            I => \N__34512\
        );

    \I__6705\ : LocalMux
    port map (
            O => \N__34615\,
            I => \N__34512\
        );

    \I__6704\ : InMux
    port map (
            O => \N__34614\,
            I => \N__34507\
        );

    \I__6703\ : InMux
    port map (
            O => \N__34613\,
            I => \N__34507\
        );

    \I__6702\ : InMux
    port map (
            O => \N__34612\,
            I => \N__34504\
        );

    \I__6701\ : InMux
    port map (
            O => \N__34611\,
            I => \N__34491\
        );

    \I__6700\ : InMux
    port map (
            O => \N__34610\,
            I => \N__34491\
        );

    \I__6699\ : InMux
    port map (
            O => \N__34609\,
            I => \N__34491\
        );

    \I__6698\ : InMux
    port map (
            O => \N__34608\,
            I => \N__34491\
        );

    \I__6697\ : InMux
    port map (
            O => \N__34607\,
            I => \N__34491\
        );

    \I__6696\ : InMux
    port map (
            O => \N__34606\,
            I => \N__34491\
        );

    \I__6695\ : InMux
    port map (
            O => \N__34605\,
            I => \N__34486\
        );

    \I__6694\ : InMux
    port map (
            O => \N__34604\,
            I => \N__34486\
        );

    \I__6693\ : InMux
    port map (
            O => \N__34603\,
            I => \N__34475\
        );

    \I__6692\ : InMux
    port map (
            O => \N__34602\,
            I => \N__34475\
        );

    \I__6691\ : InMux
    port map (
            O => \N__34601\,
            I => \N__34475\
        );

    \I__6690\ : InMux
    port map (
            O => \N__34600\,
            I => \N__34475\
        );

    \I__6689\ : InMux
    port map (
            O => \N__34599\,
            I => \N__34475\
        );

    \I__6688\ : LocalMux
    port map (
            O => \N__34590\,
            I => \N__34472\
        );

    \I__6687\ : Span4Mux_h
    port map (
            O => \N__34585\,
            I => \N__34469\
        );

    \I__6686\ : InMux
    port map (
            O => \N__34582\,
            I => \N__34464\
        );

    \I__6685\ : InMux
    port map (
            O => \N__34581\,
            I => \N__34464\
        );

    \I__6684\ : LocalMux
    port map (
            O => \N__34578\,
            I => \N__34459\
        );

    \I__6683\ : LocalMux
    port map (
            O => \N__34575\,
            I => \N__34459\
        );

    \I__6682\ : Span4Mux_v
    port map (
            O => \N__34568\,
            I => \N__34452\
        );

    \I__6681\ : LocalMux
    port map (
            O => \N__34557\,
            I => \N__34452\
        );

    \I__6680\ : Span4Mux_h
    port map (
            O => \N__34554\,
            I => \N__34452\
        );

    \I__6679\ : LocalMux
    port map (
            O => \N__34551\,
            I => \N__34435\
        );

    \I__6678\ : LocalMux
    port map (
            O => \N__34536\,
            I => \N__34435\
        );

    \I__6677\ : Span4Mux_v
    port map (
            O => \N__34533\,
            I => \N__34435\
        );

    \I__6676\ : Span4Mux_v
    port map (
            O => \N__34530\,
            I => \N__34435\
        );

    \I__6675\ : Span4Mux_v
    port map (
            O => \N__34525\,
            I => \N__34435\
        );

    \I__6674\ : Span4Mux_v
    port map (
            O => \N__34520\,
            I => \N__34435\
        );

    \I__6673\ : Span4Mux_h
    port map (
            O => \N__34517\,
            I => \N__34435\
        );

    \I__6672\ : Span4Mux_v
    port map (
            O => \N__34512\,
            I => \N__34435\
        );

    \I__6671\ : LocalMux
    port map (
            O => \N__34507\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__6670\ : LocalMux
    port map (
            O => \N__34504\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__6669\ : LocalMux
    port map (
            O => \N__34491\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__6668\ : LocalMux
    port map (
            O => \N__34486\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__6667\ : LocalMux
    port map (
            O => \N__34475\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__6666\ : Odrv4
    port map (
            O => \N__34472\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__6665\ : Odrv4
    port map (
            O => \N__34469\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__6664\ : LocalMux
    port map (
            O => \N__34464\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__6663\ : Odrv4
    port map (
            O => \N__34459\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__6662\ : Odrv4
    port map (
            O => \N__34452\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__6661\ : Odrv4
    port map (
            O => \N__34435\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__6660\ : InMux
    port map (
            O => \N__34412\,
            I => \N__34409\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__34409\,
            I => \N__34405\
        );

    \I__6658\ : InMux
    port map (
            O => \N__34408\,
            I => \N__34401\
        );

    \I__6657\ : Span4Mux_h
    port map (
            O => \N__34405\,
            I => \N__34398\
        );

    \I__6656\ : InMux
    port map (
            O => \N__34404\,
            I => \N__34395\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__34401\,
            I => \N__34390\
        );

    \I__6654\ : Span4Mux_v
    port map (
            O => \N__34398\,
            I => \N__34390\
        );

    \I__6653\ : LocalMux
    port map (
            O => \N__34395\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8\
        );

    \I__6652\ : Odrv4
    port map (
            O => \N__34390\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8\
        );

    \I__6651\ : InMux
    port map (
            O => \N__34385\,
            I => \N__34381\
        );

    \I__6650\ : InMux
    port map (
            O => \N__34384\,
            I => \N__34378\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__34381\,
            I => \N__34375\
        );

    \I__6648\ : LocalMux
    port map (
            O => \N__34378\,
            I => \N__34371\
        );

    \I__6647\ : Span4Mux_v
    port map (
            O => \N__34375\,
            I => \N__34368\
        );

    \I__6646\ : InMux
    port map (
            O => \N__34374\,
            I => \N__34365\
        );

    \I__6645\ : Span12Mux_h
    port map (
            O => \N__34371\,
            I => \N__34361\
        );

    \I__6644\ : Sp12to4
    port map (
            O => \N__34368\,
            I => \N__34356\
        );

    \I__6643\ : LocalMux
    port map (
            O => \N__34365\,
            I => \N__34356\
        );

    \I__6642\ : InMux
    port map (
            O => \N__34364\,
            I => \N__34353\
        );

    \I__6641\ : Odrv12
    port map (
            O => \N__34361\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__6640\ : Odrv12
    port map (
            O => \N__34356\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__6639\ : LocalMux
    port map (
            O => \N__34353\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__6638\ : InMux
    port map (
            O => \N__34346\,
            I => \N__34343\
        );

    \I__6637\ : LocalMux
    port map (
            O => \N__34343\,
            I => \N__34340\
        );

    \I__6636\ : Odrv4
    port map (
            O => \N__34340\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\
        );

    \I__6635\ : CEMux
    port map (
            O => \N__34337\,
            I => \N__34334\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__34334\,
            I => \N__34313\
        );

    \I__6633\ : InMux
    port map (
            O => \N__34333\,
            I => \N__34302\
        );

    \I__6632\ : InMux
    port map (
            O => \N__34332\,
            I => \N__34302\
        );

    \I__6631\ : InMux
    port map (
            O => \N__34331\,
            I => \N__34302\
        );

    \I__6630\ : InMux
    port map (
            O => \N__34330\,
            I => \N__34293\
        );

    \I__6629\ : InMux
    port map (
            O => \N__34329\,
            I => \N__34293\
        );

    \I__6628\ : InMux
    port map (
            O => \N__34328\,
            I => \N__34293\
        );

    \I__6627\ : InMux
    port map (
            O => \N__34327\,
            I => \N__34293\
        );

    \I__6626\ : InMux
    port map (
            O => \N__34326\,
            I => \N__34284\
        );

    \I__6625\ : InMux
    port map (
            O => \N__34325\,
            I => \N__34284\
        );

    \I__6624\ : InMux
    port map (
            O => \N__34324\,
            I => \N__34284\
        );

    \I__6623\ : InMux
    port map (
            O => \N__34323\,
            I => \N__34284\
        );

    \I__6622\ : CEMux
    port map (
            O => \N__34322\,
            I => \N__34281\
        );

    \I__6621\ : CEMux
    port map (
            O => \N__34321\,
            I => \N__34277\
        );

    \I__6620\ : InMux
    port map (
            O => \N__34320\,
            I => \N__34267\
        );

    \I__6619\ : InMux
    port map (
            O => \N__34319\,
            I => \N__34267\
        );

    \I__6618\ : InMux
    port map (
            O => \N__34318\,
            I => \N__34267\
        );

    \I__6617\ : InMux
    port map (
            O => \N__34317\,
            I => \N__34267\
        );

    \I__6616\ : CEMux
    port map (
            O => \N__34316\,
            I => \N__34264\
        );

    \I__6615\ : Span4Mux_v
    port map (
            O => \N__34313\,
            I => \N__34258\
        );

    \I__6614\ : CEMux
    port map (
            O => \N__34312\,
            I => \N__34255\
        );

    \I__6613\ : InMux
    port map (
            O => \N__34311\,
            I => \N__34247\
        );

    \I__6612\ : InMux
    port map (
            O => \N__34310\,
            I => \N__34247\
        );

    \I__6611\ : InMux
    port map (
            O => \N__34309\,
            I => \N__34247\
        );

    \I__6610\ : LocalMux
    port map (
            O => \N__34302\,
            I => \N__34238\
        );

    \I__6609\ : LocalMux
    port map (
            O => \N__34293\,
            I => \N__34238\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__34284\,
            I => \N__34238\
        );

    \I__6607\ : LocalMux
    port map (
            O => \N__34281\,
            I => \N__34238\
        );

    \I__6606\ : CEMux
    port map (
            O => \N__34280\,
            I => \N__34223\
        );

    \I__6605\ : LocalMux
    port map (
            O => \N__34277\,
            I => \N__34220\
        );

    \I__6604\ : CEMux
    port map (
            O => \N__34276\,
            I => \N__34217\
        );

    \I__6603\ : LocalMux
    port map (
            O => \N__34267\,
            I => \N__34212\
        );

    \I__6602\ : LocalMux
    port map (
            O => \N__34264\,
            I => \N__34212\
        );

    \I__6601\ : CEMux
    port map (
            O => \N__34263\,
            I => \N__34209\
        );

    \I__6600\ : CEMux
    port map (
            O => \N__34262\,
            I => \N__34206\
        );

    \I__6599\ : CEMux
    port map (
            O => \N__34261\,
            I => \N__34203\
        );

    \I__6598\ : Span4Mux_h
    port map (
            O => \N__34258\,
            I => \N__34197\
        );

    \I__6597\ : LocalMux
    port map (
            O => \N__34255\,
            I => \N__34197\
        );

    \I__6596\ : CEMux
    port map (
            O => \N__34254\,
            I => \N__34194\
        );

    \I__6595\ : LocalMux
    port map (
            O => \N__34247\,
            I => \N__34189\
        );

    \I__6594\ : Span4Mux_v
    port map (
            O => \N__34238\,
            I => \N__34189\
        );

    \I__6593\ : InMux
    port map (
            O => \N__34237\,
            I => \N__34180\
        );

    \I__6592\ : InMux
    port map (
            O => \N__34236\,
            I => \N__34180\
        );

    \I__6591\ : InMux
    port map (
            O => \N__34235\,
            I => \N__34180\
        );

    \I__6590\ : InMux
    port map (
            O => \N__34234\,
            I => \N__34180\
        );

    \I__6589\ : InMux
    port map (
            O => \N__34233\,
            I => \N__34171\
        );

    \I__6588\ : InMux
    port map (
            O => \N__34232\,
            I => \N__34171\
        );

    \I__6587\ : InMux
    port map (
            O => \N__34231\,
            I => \N__34171\
        );

    \I__6586\ : InMux
    port map (
            O => \N__34230\,
            I => \N__34171\
        );

    \I__6585\ : InMux
    port map (
            O => \N__34229\,
            I => \N__34162\
        );

    \I__6584\ : InMux
    port map (
            O => \N__34228\,
            I => \N__34162\
        );

    \I__6583\ : InMux
    port map (
            O => \N__34227\,
            I => \N__34162\
        );

    \I__6582\ : InMux
    port map (
            O => \N__34226\,
            I => \N__34162\
        );

    \I__6581\ : LocalMux
    port map (
            O => \N__34223\,
            I => \N__34159\
        );

    \I__6580\ : Span4Mux_v
    port map (
            O => \N__34220\,
            I => \N__34154\
        );

    \I__6579\ : LocalMux
    port map (
            O => \N__34217\,
            I => \N__34154\
        );

    \I__6578\ : Span4Mux_h
    port map (
            O => \N__34212\,
            I => \N__34151\
        );

    \I__6577\ : LocalMux
    port map (
            O => \N__34209\,
            I => \N__34148\
        );

    \I__6576\ : LocalMux
    port map (
            O => \N__34206\,
            I => \N__34145\
        );

    \I__6575\ : LocalMux
    port map (
            O => \N__34203\,
            I => \N__34142\
        );

    \I__6574\ : CEMux
    port map (
            O => \N__34202\,
            I => \N__34138\
        );

    \I__6573\ : Span4Mux_h
    port map (
            O => \N__34197\,
            I => \N__34135\
        );

    \I__6572\ : LocalMux
    port map (
            O => \N__34194\,
            I => \N__34132\
        );

    \I__6571\ : Span4Mux_h
    port map (
            O => \N__34189\,
            I => \N__34121\
        );

    \I__6570\ : LocalMux
    port map (
            O => \N__34180\,
            I => \N__34121\
        );

    \I__6569\ : LocalMux
    port map (
            O => \N__34171\,
            I => \N__34121\
        );

    \I__6568\ : LocalMux
    port map (
            O => \N__34162\,
            I => \N__34121\
        );

    \I__6567\ : Span4Mux_h
    port map (
            O => \N__34159\,
            I => \N__34121\
        );

    \I__6566\ : Span4Mux_v
    port map (
            O => \N__34154\,
            I => \N__34118\
        );

    \I__6565\ : Span4Mux_v
    port map (
            O => \N__34151\,
            I => \N__34115\
        );

    \I__6564\ : Span4Mux_h
    port map (
            O => \N__34148\,
            I => \N__34110\
        );

    \I__6563\ : Span4Mux_v
    port map (
            O => \N__34145\,
            I => \N__34110\
        );

    \I__6562\ : Span4Mux_v
    port map (
            O => \N__34142\,
            I => \N__34107\
        );

    \I__6561\ : InMux
    port map (
            O => \N__34141\,
            I => \N__34104\
        );

    \I__6560\ : LocalMux
    port map (
            O => \N__34138\,
            I => \N__34099\
        );

    \I__6559\ : Sp12to4
    port map (
            O => \N__34135\,
            I => \N__34099\
        );

    \I__6558\ : Span4Mux_h
    port map (
            O => \N__34132\,
            I => \N__34094\
        );

    \I__6557\ : Span4Mux_v
    port map (
            O => \N__34121\,
            I => \N__34094\
        );

    \I__6556\ : Span4Mux_h
    port map (
            O => \N__34118\,
            I => \N__34089\
        );

    \I__6555\ : Span4Mux_h
    port map (
            O => \N__34115\,
            I => \N__34089\
        );

    \I__6554\ : Odrv4
    port map (
            O => \N__34110\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__6553\ : Odrv4
    port map (
            O => \N__34107\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__6552\ : LocalMux
    port map (
            O => \N__34104\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__6551\ : Odrv12
    port map (
            O => \N__34099\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__6550\ : Odrv4
    port map (
            O => \N__34094\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__6549\ : Odrv4
    port map (
            O => \N__34089\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__6548\ : InMux
    port map (
            O => \N__34076\,
            I => \N__34070\
        );

    \I__6547\ : InMux
    port map (
            O => \N__34075\,
            I => \N__34070\
        );

    \I__6546\ : LocalMux
    port map (
            O => \N__34070\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_22\
        );

    \I__6545\ : IoInMux
    port map (
            O => \N__34067\,
            I => \N__34064\
        );

    \I__6544\ : LocalMux
    port map (
            O => \N__34064\,
            I => \N__34061\
        );

    \I__6543\ : Span4Mux_s0_v
    port map (
            O => \N__34061\,
            I => \N__34058\
        );

    \I__6542\ : Odrv4
    port map (
            O => \N__34058\,
            I => \pll_inst.red_c_i\
        );

    \I__6541\ : ClkMux
    port map (
            O => \N__34055\,
            I => \N__34049\
        );

    \I__6540\ : ClkMux
    port map (
            O => \N__34054\,
            I => \N__34049\
        );

    \I__6539\ : GlobalMux
    port map (
            O => \N__34049\,
            I => \N__34046\
        );

    \I__6538\ : gio2CtrlBuf
    port map (
            O => \N__34046\,
            I => delay_hc_input_c_g
        );

    \I__6537\ : InMux
    port map (
            O => \N__34043\,
            I => \N__34040\
        );

    \I__6536\ : LocalMux
    port map (
            O => \N__34040\,
            I => \N__34035\
        );

    \I__6535\ : InMux
    port map (
            O => \N__34039\,
            I => \N__34032\
        );

    \I__6534\ : InMux
    port map (
            O => \N__34038\,
            I => \N__34029\
        );

    \I__6533\ : Span4Mux_v
    port map (
            O => \N__34035\,
            I => \N__34026\
        );

    \I__6532\ : LocalMux
    port map (
            O => \N__34032\,
            I => \N__34023\
        );

    \I__6531\ : LocalMux
    port map (
            O => \N__34029\,
            I => \N__34020\
        );

    \I__6530\ : Span4Mux_v
    port map (
            O => \N__34026\,
            I => \N__34014\
        );

    \I__6529\ : Span4Mux_v
    port map (
            O => \N__34023\,
            I => \N__34014\
        );

    \I__6528\ : Span12Mux_v
    port map (
            O => \N__34020\,
            I => \N__34011\
        );

    \I__6527\ : InMux
    port map (
            O => \N__34019\,
            I => \N__34008\
        );

    \I__6526\ : Odrv4
    port map (
            O => \N__34014\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__6525\ : Odrv12
    port map (
            O => \N__34011\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__6524\ : LocalMux
    port map (
            O => \N__34008\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__6523\ : InMux
    port map (
            O => \N__34001\,
            I => \N__33998\
        );

    \I__6522\ : LocalMux
    port map (
            O => \N__33998\,
            I => \N__33993\
        );

    \I__6521\ : InMux
    port map (
            O => \N__33997\,
            I => \N__33990\
        );

    \I__6520\ : InMux
    port map (
            O => \N__33996\,
            I => \N__33987\
        );

    \I__6519\ : Span4Mux_h
    port map (
            O => \N__33993\,
            I => \N__33984\
        );

    \I__6518\ : LocalMux
    port map (
            O => \N__33990\,
            I => \N__33981\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__33987\,
            I => \N__33974\
        );

    \I__6516\ : Span4Mux_v
    port map (
            O => \N__33984\,
            I => \N__33974\
        );

    \I__6515\ : Span4Mux_v
    port map (
            O => \N__33981\,
            I => \N__33974\
        );

    \I__6514\ : Odrv4
    port map (
            O => \N__33974\,
            I => \elapsed_time_ns_1_RNIED91B_0_2\
        );

    \I__6513\ : CascadeMux
    port map (
            O => \N__33971\,
            I => \N__33968\
        );

    \I__6512\ : InMux
    port map (
            O => \N__33968\,
            I => \N__33965\
        );

    \I__6511\ : LocalMux
    port map (
            O => \N__33965\,
            I => \N__33962\
        );

    \I__6510\ : Span4Mux_h
    port map (
            O => \N__33962\,
            I => \N__33959\
        );

    \I__6509\ : Odrv4
    port map (
            O => \N__33959\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt24\
        );

    \I__6508\ : InMux
    port map (
            O => \N__33956\,
            I => \N__33951\
        );

    \I__6507\ : InMux
    port map (
            O => \N__33955\,
            I => \N__33946\
        );

    \I__6506\ : InMux
    port map (
            O => \N__33954\,
            I => \N__33946\
        );

    \I__6505\ : LocalMux
    port map (
            O => \N__33951\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__6504\ : LocalMux
    port map (
            O => \N__33946\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__6503\ : CascadeMux
    port map (
            O => \N__33941\,
            I => \N__33938\
        );

    \I__6502\ : InMux
    port map (
            O => \N__33938\,
            I => \N__33931\
        );

    \I__6501\ : InMux
    port map (
            O => \N__33937\,
            I => \N__33931\
        );

    \I__6500\ : InMux
    port map (
            O => \N__33936\,
            I => \N__33928\
        );

    \I__6499\ : LocalMux
    port map (
            O => \N__33931\,
            I => \N__33925\
        );

    \I__6498\ : LocalMux
    port map (
            O => \N__33928\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__6497\ : Odrv4
    port map (
            O => \N__33925\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__6496\ : InMux
    port map (
            O => \N__33920\,
            I => \N__33917\
        );

    \I__6495\ : LocalMux
    port map (
            O => \N__33917\,
            I => \N__33914\
        );

    \I__6494\ : Span4Mux_h
    port map (
            O => \N__33914\,
            I => \N__33911\
        );

    \I__6493\ : Odrv4
    port map (
            O => \N__33911\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24\
        );

    \I__6492\ : InMux
    port map (
            O => \N__33908\,
            I => \N__33905\
        );

    \I__6491\ : LocalMux
    port map (
            O => \N__33905\,
            I => \N__33902\
        );

    \I__6490\ : Span4Mux_v
    port map (
            O => \N__33902\,
            I => \N__33897\
        );

    \I__6489\ : InMux
    port map (
            O => \N__33901\,
            I => \N__33894\
        );

    \I__6488\ : InMux
    port map (
            O => \N__33900\,
            I => \N__33891\
        );

    \I__6487\ : Span4Mux_h
    port map (
            O => \N__33897\,
            I => \N__33888\
        );

    \I__6486\ : LocalMux
    port map (
            O => \N__33894\,
            I => \N__33885\
        );

    \I__6485\ : LocalMux
    port map (
            O => \N__33891\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25\
        );

    \I__6484\ : Odrv4
    port map (
            O => \N__33888\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25\
        );

    \I__6483\ : Odrv4
    port map (
            O => \N__33885\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25\
        );

    \I__6482\ : InMux
    port map (
            O => \N__33878\,
            I => \N__33875\
        );

    \I__6481\ : LocalMux
    port map (
            O => \N__33875\,
            I => \N__33871\
        );

    \I__6480\ : InMux
    port map (
            O => \N__33874\,
            I => \N__33867\
        );

    \I__6479\ : Span4Mux_h
    port map (
            O => \N__33871\,
            I => \N__33864\
        );

    \I__6478\ : InMux
    port map (
            O => \N__33870\,
            I => \N__33861\
        );

    \I__6477\ : LocalMux
    port map (
            O => \N__33867\,
            I => \N__33857\
        );

    \I__6476\ : Span4Mux_h
    port map (
            O => \N__33864\,
            I => \N__33852\
        );

    \I__6475\ : LocalMux
    port map (
            O => \N__33861\,
            I => \N__33852\
        );

    \I__6474\ : InMux
    port map (
            O => \N__33860\,
            I => \N__33849\
        );

    \I__6473\ : Odrv4
    port map (
            O => \N__33857\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__6472\ : Odrv4
    port map (
            O => \N__33852\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__33849\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__6470\ : CascadeMux
    port map (
            O => \N__33842\,
            I => \N__33839\
        );

    \I__6469\ : InMux
    port map (
            O => \N__33839\,
            I => \N__33833\
        );

    \I__6468\ : InMux
    port map (
            O => \N__33838\,
            I => \N__33833\
        );

    \I__6467\ : LocalMux
    port map (
            O => \N__33833\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_25\
        );

    \I__6466\ : InMux
    port map (
            O => \N__33830\,
            I => \N__33827\
        );

    \I__6465\ : LocalMux
    port map (
            O => \N__33827\,
            I => \N__33824\
        );

    \I__6464\ : Span4Mux_h
    port map (
            O => \N__33824\,
            I => \N__33820\
        );

    \I__6463\ : InMux
    port map (
            O => \N__33823\,
            I => \N__33817\
        );

    \I__6462\ : Odrv4
    port map (
            O => \N__33820\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24\
        );

    \I__6461\ : LocalMux
    port map (
            O => \N__33817\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24\
        );

    \I__6460\ : InMux
    port map (
            O => \N__33812\,
            I => \current_shift_inst.un38_control_input_cry_25_s0\
        );

    \I__6459\ : InMux
    port map (
            O => \N__33809\,
            I => \current_shift_inst.un38_control_input_cry_26_s0\
        );

    \I__6458\ : InMux
    port map (
            O => \N__33806\,
            I => \current_shift_inst.un38_control_input_cry_27_s0\
        );

    \I__6457\ : InMux
    port map (
            O => \N__33803\,
            I => \current_shift_inst.un38_control_input_cry_28_s0\
        );

    \I__6456\ : InMux
    port map (
            O => \N__33800\,
            I => \N__33797\
        );

    \I__6455\ : LocalMux
    port map (
            O => \N__33797\,
            I => \current_shift_inst.un38_control_input_0_s0_30\
        );

    \I__6454\ : InMux
    port map (
            O => \N__33794\,
            I => \current_shift_inst.un38_control_input_cry_29_s0\
        );

    \I__6453\ : InMux
    port map (
            O => \N__33791\,
            I => \current_shift_inst.un38_control_input_cry_30_s0\
        );

    \I__6452\ : InMux
    port map (
            O => \N__33788\,
            I => \N__33785\
        );

    \I__6451\ : LocalMux
    port map (
            O => \N__33785\,
            I => \current_shift_inst.control_input_axb_28\
        );

    \I__6450\ : InMux
    port map (
            O => \N__33782\,
            I => \N__33779\
        );

    \I__6449\ : LocalMux
    port map (
            O => \N__33779\,
            I => \N__33776\
        );

    \I__6448\ : Odrv4
    port map (
            O => \N__33776\,
            I => \current_shift_inst.control_input_axb_29\
        );

    \I__6447\ : InMux
    port map (
            O => \N__33773\,
            I => \current_shift_inst.un38_control_input_cry_16_s0\
        );

    \I__6446\ : InMux
    port map (
            O => \N__33770\,
            I => \current_shift_inst.un38_control_input_cry_17_s0\
        );

    \I__6445\ : InMux
    port map (
            O => \N__33767\,
            I => \current_shift_inst.un38_control_input_cry_18_s0\
        );

    \I__6444\ : InMux
    port map (
            O => \N__33764\,
            I => \N__33761\
        );

    \I__6443\ : LocalMux
    port map (
            O => \N__33761\,
            I => \current_shift_inst.un38_control_input_0_s0_20\
        );

    \I__6442\ : InMux
    port map (
            O => \N__33758\,
            I => \current_shift_inst.un38_control_input_cry_19_s0\
        );

    \I__6441\ : InMux
    port map (
            O => \N__33755\,
            I => \N__33752\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__33752\,
            I => \current_shift_inst.un38_control_input_0_s0_21\
        );

    \I__6439\ : InMux
    port map (
            O => \N__33749\,
            I => \current_shift_inst.un38_control_input_cry_20_s0\
        );

    \I__6438\ : InMux
    port map (
            O => \N__33746\,
            I => \N__33743\
        );

    \I__6437\ : LocalMux
    port map (
            O => \N__33743\,
            I => \N__33740\
        );

    \I__6436\ : Span4Mux_h
    port map (
            O => \N__33740\,
            I => \N__33737\
        );

    \I__6435\ : Odrv4
    port map (
            O => \N__33737\,
            I => \current_shift_inst.un38_control_input_0_s0_22\
        );

    \I__6434\ : InMux
    port map (
            O => \N__33734\,
            I => \current_shift_inst.un38_control_input_cry_21_s0\
        );

    \I__6433\ : InMux
    port map (
            O => \N__33731\,
            I => \current_shift_inst.un38_control_input_cry_22_s0\
        );

    \I__6432\ : InMux
    port map (
            O => \N__33728\,
            I => \bfn_12_19_0_\
        );

    \I__6431\ : InMux
    port map (
            O => \N__33725\,
            I => \current_shift_inst.un38_control_input_cry_24_s0\
        );

    \I__6430\ : InMux
    port map (
            O => \N__33722\,
            I => \N__33719\
        );

    \I__6429\ : LocalMux
    port map (
            O => \N__33719\,
            I => \N__33716\
        );

    \I__6428\ : Odrv4
    port map (
            O => \N__33716\,
            I => \current_shift_inst.un38_control_input_0_s0_9\
        );

    \I__6427\ : InMux
    port map (
            O => \N__33713\,
            I => \current_shift_inst.un38_control_input_cry_8_s0\
        );

    \I__6426\ : InMux
    port map (
            O => \N__33710\,
            I => \current_shift_inst.un38_control_input_cry_9_s0\
        );

    \I__6425\ : InMux
    port map (
            O => \N__33707\,
            I => \N__33704\
        );

    \I__6424\ : LocalMux
    port map (
            O => \N__33704\,
            I => \N__33701\
        );

    \I__6423\ : Span4Mux_v
    port map (
            O => \N__33701\,
            I => \N__33698\
        );

    \I__6422\ : Odrv4
    port map (
            O => \N__33698\,
            I => \current_shift_inst.un38_control_input_0_s0_11\
        );

    \I__6421\ : InMux
    port map (
            O => \N__33695\,
            I => \current_shift_inst.un38_control_input_cry_10_s0\
        );

    \I__6420\ : InMux
    port map (
            O => \N__33692\,
            I => \N__33689\
        );

    \I__6419\ : LocalMux
    port map (
            O => \N__33689\,
            I => \N__33686\
        );

    \I__6418\ : Span4Mux_h
    port map (
            O => \N__33686\,
            I => \N__33683\
        );

    \I__6417\ : Odrv4
    port map (
            O => \N__33683\,
            I => \current_shift_inst.un38_control_input_0_s0_12\
        );

    \I__6416\ : InMux
    port map (
            O => \N__33680\,
            I => \current_shift_inst.un38_control_input_cry_11_s0\
        );

    \I__6415\ : InMux
    port map (
            O => \N__33677\,
            I => \N__33674\
        );

    \I__6414\ : LocalMux
    port map (
            O => \N__33674\,
            I => \N__33671\
        );

    \I__6413\ : Span4Mux_h
    port map (
            O => \N__33671\,
            I => \N__33668\
        );

    \I__6412\ : Odrv4
    port map (
            O => \N__33668\,
            I => \current_shift_inst.un38_control_input_0_s0_13\
        );

    \I__6411\ : InMux
    port map (
            O => \N__33665\,
            I => \current_shift_inst.un38_control_input_cry_12_s0\
        );

    \I__6410\ : InMux
    port map (
            O => \N__33662\,
            I => \current_shift_inst.un38_control_input_cry_13_s0\
        );

    \I__6409\ : InMux
    port map (
            O => \N__33659\,
            I => \current_shift_inst.un38_control_input_cry_14_s0\
        );

    \I__6408\ : InMux
    port map (
            O => \N__33656\,
            I => \bfn_12_18_0_\
        );

    \I__6407\ : InMux
    port map (
            O => \N__33653\,
            I => \N__33650\
        );

    \I__6406\ : LocalMux
    port map (
            O => \N__33650\,
            I => \N__33647\
        );

    \I__6405\ : Span4Mux_h
    port map (
            O => \N__33647\,
            I => \N__33644\
        );

    \I__6404\ : Odrv4
    port map (
            O => \N__33644\,
            I => \current_shift_inst.un38_control_input_0_s0_3\
        );

    \I__6403\ : InMux
    port map (
            O => \N__33641\,
            I => \current_shift_inst.un38_control_input_cry_2_s0\
        );

    \I__6402\ : CascadeMux
    port map (
            O => \N__33638\,
            I => \N__33635\
        );

    \I__6401\ : InMux
    port map (
            O => \N__33635\,
            I => \N__33632\
        );

    \I__6400\ : LocalMux
    port map (
            O => \N__33632\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5\
        );

    \I__6399\ : InMux
    port map (
            O => \N__33629\,
            I => \N__33626\
        );

    \I__6398\ : LocalMux
    port map (
            O => \N__33626\,
            I => \current_shift_inst.un38_control_input_0_s0_4\
        );

    \I__6397\ : InMux
    port map (
            O => \N__33623\,
            I => \current_shift_inst.un38_control_input_cry_3_s0\
        );

    \I__6396\ : InMux
    port map (
            O => \N__33620\,
            I => \N__33617\
        );

    \I__6395\ : LocalMux
    port map (
            O => \N__33617\,
            I => \current_shift_inst.un38_control_input_0_s0_5\
        );

    \I__6394\ : InMux
    port map (
            O => \N__33614\,
            I => \current_shift_inst.un38_control_input_cry_4_s0\
        );

    \I__6393\ : InMux
    port map (
            O => \N__33611\,
            I => \N__33608\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__33608\,
            I => \current_shift_inst.un38_control_input_0_s0_6\
        );

    \I__6391\ : InMux
    port map (
            O => \N__33605\,
            I => \current_shift_inst.un38_control_input_cry_5_s0\
        );

    \I__6390\ : InMux
    port map (
            O => \N__33602\,
            I => \N__33599\
        );

    \I__6389\ : LocalMux
    port map (
            O => \N__33599\,
            I => \current_shift_inst.un38_control_input_0_s0_7\
        );

    \I__6388\ : InMux
    port map (
            O => \N__33596\,
            I => \current_shift_inst.un38_control_input_cry_6_s0\
        );

    \I__6387\ : InMux
    port map (
            O => \N__33593\,
            I => \N__33590\
        );

    \I__6386\ : LocalMux
    port map (
            O => \N__33590\,
            I => \N__33587\
        );

    \I__6385\ : Odrv4
    port map (
            O => \N__33587\,
            I => \current_shift_inst.un38_control_input_0_s0_8\
        );

    \I__6384\ : InMux
    port map (
            O => \N__33584\,
            I => \bfn_12_17_0_\
        );

    \I__6383\ : InMux
    port map (
            O => \N__33581\,
            I => \N__33578\
        );

    \I__6382\ : LocalMux
    port map (
            O => \N__33578\,
            I => \N__33575\
        );

    \I__6381\ : Span4Mux_h
    port map (
            O => \N__33575\,
            I => \N__33572\
        );

    \I__6380\ : Span4Mux_h
    port map (
            O => \N__33572\,
            I => \N__33568\
        );

    \I__6379\ : InMux
    port map (
            O => \N__33571\,
            I => \N__33565\
        );

    \I__6378\ : Odrv4
    port map (
            O => \N__33568\,
            I => state_ns_i_a3_1
        );

    \I__6377\ : LocalMux
    port map (
            O => \N__33565\,
            I => state_ns_i_a3_1
        );

    \I__6376\ : InMux
    port map (
            O => \N__33560\,
            I => \N__33557\
        );

    \I__6375\ : LocalMux
    port map (
            O => \N__33557\,
            I => \N__33554\
        );

    \I__6374\ : Span4Mux_h
    port map (
            O => \N__33554\,
            I => \N__33550\
        );

    \I__6373\ : InMux
    port map (
            O => \N__33553\,
            I => \N__33547\
        );

    \I__6372\ : Span4Mux_v
    port map (
            O => \N__33550\,
            I => \N__33540\
        );

    \I__6371\ : LocalMux
    port map (
            O => \N__33547\,
            I => \N__33540\
        );

    \I__6370\ : InMux
    port map (
            O => \N__33546\,
            I => \N__33535\
        );

    \I__6369\ : InMux
    port map (
            O => \N__33545\,
            I => \N__33535\
        );

    \I__6368\ : Sp12to4
    port map (
            O => \N__33540\,
            I => \N__33532\
        );

    \I__6367\ : LocalMux
    port map (
            O => \N__33535\,
            I => \N__33529\
        );

    \I__6366\ : Span12Mux_v
    port map (
            O => \N__33532\,
            I => \N__33526\
        );

    \I__6365\ : Span4Mux_v
    port map (
            O => \N__33529\,
            I => \N__33523\
        );

    \I__6364\ : Span12Mux_v
    port map (
            O => \N__33526\,
            I => \N__33520\
        );

    \I__6363\ : Sp12to4
    port map (
            O => \N__33523\,
            I => \N__33517\
        );

    \I__6362\ : Span12Mux_h
    port map (
            O => \N__33520\,
            I => \N__33514\
        );

    \I__6361\ : Span12Mux_h
    port map (
            O => \N__33517\,
            I => \N__33511\
        );

    \I__6360\ : Odrv12
    port map (
            O => \N__33514\,
            I => start_stop_c
        );

    \I__6359\ : Odrv12
    port map (
            O => \N__33511\,
            I => start_stop_c
        );

    \I__6358\ : InMux
    port map (
            O => \N__33506\,
            I => \N__33503\
        );

    \I__6357\ : LocalMux
    port map (
            O => \N__33503\,
            I => \current_shift_inst.control_input_axb_1\
        );

    \I__6356\ : InMux
    port map (
            O => \N__33500\,
            I => \N__33497\
        );

    \I__6355\ : LocalMux
    port map (
            O => \N__33497\,
            I => \current_shift_inst.control_input_axb_2\
        );

    \I__6354\ : InMux
    port map (
            O => \N__33494\,
            I => \N__33491\
        );

    \I__6353\ : LocalMux
    port map (
            O => \N__33491\,
            I => \current_shift_inst.control_input_axb_3\
        );

    \I__6352\ : InMux
    port map (
            O => \N__33488\,
            I => \N__33485\
        );

    \I__6351\ : LocalMux
    port map (
            O => \N__33485\,
            I => \current_shift_inst.control_input_axb_4\
        );

    \I__6350\ : InMux
    port map (
            O => \N__33482\,
            I => \N__33479\
        );

    \I__6349\ : LocalMux
    port map (
            O => \N__33479\,
            I => \current_shift_inst.control_input_axb_5\
        );

    \I__6348\ : InMux
    port map (
            O => \N__33476\,
            I => \N__33473\
        );

    \I__6347\ : LocalMux
    port map (
            O => \N__33473\,
            I => \current_shift_inst.control_input_axb_6\
        );

    \I__6346\ : InMux
    port map (
            O => \N__33470\,
            I => \N__33461\
        );

    \I__6345\ : InMux
    port map (
            O => \N__33469\,
            I => \N__33461\
        );

    \I__6344\ : InMux
    port map (
            O => \N__33468\,
            I => \N__33461\
        );

    \I__6343\ : LocalMux
    port map (
            O => \N__33461\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__6342\ : CascadeMux
    port map (
            O => \N__33458\,
            I => \N__33454\
        );

    \I__6341\ : InMux
    port map (
            O => \N__33457\,
            I => \N__33450\
        );

    \I__6340\ : InMux
    port map (
            O => \N__33454\,
            I => \N__33447\
        );

    \I__6339\ : InMux
    port map (
            O => \N__33453\,
            I => \N__33444\
        );

    \I__6338\ : LocalMux
    port map (
            O => \N__33450\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__6337\ : LocalMux
    port map (
            O => \N__33447\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__6336\ : LocalMux
    port map (
            O => \N__33444\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__6335\ : CascadeMux
    port map (
            O => \N__33437\,
            I => \phase_controller_inst1.state_RNI7NN7Z0Z_0_cascade_\
        );

    \I__6334\ : InMux
    port map (
            O => \N__33434\,
            I => \N__33431\
        );

    \I__6333\ : LocalMux
    port map (
            O => \N__33431\,
            I => \N__33428\
        );

    \I__6332\ : Span4Mux_h
    port map (
            O => \N__33428\,
            I => \N__33424\
        );

    \I__6331\ : InMux
    port map (
            O => \N__33427\,
            I => \N__33421\
        );

    \I__6330\ : Odrv4
    port map (
            O => \N__33424\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17\
        );

    \I__6329\ : LocalMux
    port map (
            O => \N__33421\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17\
        );

    \I__6328\ : CascadeMux
    port map (
            O => \N__33416\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17_cascade_\
        );

    \I__6327\ : CascadeMux
    port map (
            O => \N__33413\,
            I => \N__33408\
        );

    \I__6326\ : InMux
    port map (
            O => \N__33412\,
            I => \N__33405\
        );

    \I__6325\ : InMux
    port map (
            O => \N__33411\,
            I => \N__33400\
        );

    \I__6324\ : InMux
    port map (
            O => \N__33408\,
            I => \N__33400\
        );

    \I__6323\ : LocalMux
    port map (
            O => \N__33405\,
            I => \N__33396\
        );

    \I__6322\ : LocalMux
    port map (
            O => \N__33400\,
            I => \N__33393\
        );

    \I__6321\ : CascadeMux
    port map (
            O => \N__33399\,
            I => \N__33390\
        );

    \I__6320\ : Span12Mux_v
    port map (
            O => \N__33396\,
            I => \N__33387\
        );

    \I__6319\ : Span4Mux_h
    port map (
            O => \N__33393\,
            I => \N__33384\
        );

    \I__6318\ : InMux
    port map (
            O => \N__33390\,
            I => \N__33381\
        );

    \I__6317\ : Odrv12
    port map (
            O => \N__33387\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__6316\ : Odrv4
    port map (
            O => \N__33384\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__6315\ : LocalMux
    port map (
            O => \N__33381\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__6314\ : CascadeMux
    port map (
            O => \N__33374\,
            I => \N__33371\
        );

    \I__6313\ : InMux
    port map (
            O => \N__33371\,
            I => \N__33368\
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__33368\,
            I => \N__33365\
        );

    \I__6311\ : Span4Mux_h
    port map (
            O => \N__33365\,
            I => \N__33362\
        );

    \I__6310\ : Odrv4
    port map (
            O => \N__33362\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\
        );

    \I__6309\ : CascadeMux
    port map (
            O => \N__33359\,
            I => \N__33356\
        );

    \I__6308\ : InMux
    port map (
            O => \N__33356\,
            I => \N__33349\
        );

    \I__6307\ : InMux
    port map (
            O => \N__33355\,
            I => \N__33349\
        );

    \I__6306\ : InMux
    port map (
            O => \N__33354\,
            I => \N__33346\
        );

    \I__6305\ : LocalMux
    port map (
            O => \N__33349\,
            I => \N__33343\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__33346\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__6303\ : Odrv4
    port map (
            O => \N__33343\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__6302\ : CascadeMux
    port map (
            O => \N__33338\,
            I => \N__33335\
        );

    \I__6301\ : InMux
    port map (
            O => \N__33335\,
            I => \N__33329\
        );

    \I__6300\ : InMux
    port map (
            O => \N__33334\,
            I => \N__33329\
        );

    \I__6299\ : LocalMux
    port map (
            O => \N__33329\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\
        );

    \I__6298\ : InMux
    port map (
            O => \N__33326\,
            I => \N__33319\
        );

    \I__6297\ : InMux
    port map (
            O => \N__33325\,
            I => \N__33319\
        );

    \I__6296\ : InMux
    port map (
            O => \N__33324\,
            I => \N__33316\
        );

    \I__6295\ : LocalMux
    port map (
            O => \N__33319\,
            I => \N__33313\
        );

    \I__6294\ : LocalMux
    port map (
            O => \N__33316\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__6293\ : Odrv12
    port map (
            O => \N__33313\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__6292\ : InMux
    port map (
            O => \N__33308\,
            I => \N__33305\
        );

    \I__6291\ : LocalMux
    port map (
            O => \N__33305\,
            I => \N__33302\
        );

    \I__6290\ : Odrv4
    port map (
            O => \N__33302\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt16\
        );

    \I__6289\ : InMux
    port map (
            O => \N__33299\,
            I => \N__33296\
        );

    \I__6288\ : LocalMux
    port map (
            O => \N__33296\,
            I => \N__33293\
        );

    \I__6287\ : Span4Mux_h
    port map (
            O => \N__33293\,
            I => \N__33289\
        );

    \I__6286\ : InMux
    port map (
            O => \N__33292\,
            I => \N__33286\
        );

    \I__6285\ : Odrv4
    port map (
            O => \N__33289\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16\
        );

    \I__6284\ : LocalMux
    port map (
            O => \N__33286\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16\
        );

    \I__6283\ : InMux
    port map (
            O => \N__33281\,
            I => \N__33278\
        );

    \I__6282\ : LocalMux
    port map (
            O => \N__33278\,
            I => \N__33273\
        );

    \I__6281\ : InMux
    port map (
            O => \N__33277\,
            I => \N__33268\
        );

    \I__6280\ : InMux
    port map (
            O => \N__33276\,
            I => \N__33268\
        );

    \I__6279\ : Span4Mux_v
    port map (
            O => \N__33273\,
            I => \N__33264\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__33268\,
            I => \N__33261\
        );

    \I__6277\ : CascadeMux
    port map (
            O => \N__33267\,
            I => \N__33258\
        );

    \I__6276\ : Span4Mux_v
    port map (
            O => \N__33264\,
            I => \N__33255\
        );

    \I__6275\ : Span4Mux_v
    port map (
            O => \N__33261\,
            I => \N__33252\
        );

    \I__6274\ : InMux
    port map (
            O => \N__33258\,
            I => \N__33249\
        );

    \I__6273\ : Odrv4
    port map (
            O => \N__33255\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__6272\ : Odrv4
    port map (
            O => \N__33252\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__6271\ : LocalMux
    port map (
            O => \N__33249\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__6270\ : CascadeMux
    port map (
            O => \N__33242\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16_cascade_\
        );

    \I__6269\ : InMux
    port map (
            O => \N__33239\,
            I => \N__33233\
        );

    \I__6268\ : InMux
    port map (
            O => \N__33238\,
            I => \N__33233\
        );

    \I__6267\ : LocalMux
    port map (
            O => \N__33233\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\
        );

    \I__6266\ : InMux
    port map (
            O => \N__33230\,
            I => \N__33227\
        );

    \I__6265\ : LocalMux
    port map (
            O => \N__33227\,
            I => \N__33223\
        );

    \I__6264\ : InMux
    port map (
            O => \N__33226\,
            I => \N__33220\
        );

    \I__6263\ : Span4Mux_v
    port map (
            O => \N__33223\,
            I => \N__33217\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__33220\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\
        );

    \I__6261\ : Odrv4
    port map (
            O => \N__33217\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\
        );

    \I__6260\ : CascadeMux
    port map (
            O => \N__33212\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\
        );

    \I__6259\ : InMux
    port map (
            O => \N__33209\,
            I => \N__33206\
        );

    \I__6258\ : LocalMux
    port map (
            O => \N__33206\,
            I => \N__33203\
        );

    \I__6257\ : Span4Mux_v
    port map (
            O => \N__33203\,
            I => \N__33200\
        );

    \I__6256\ : Odrv4
    port map (
            O => \N__33200\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1Z0Z_30\
        );

    \I__6255\ : CascadeMux
    port map (
            O => \N__33197\,
            I => \N__33192\
        );

    \I__6254\ : InMux
    port map (
            O => \N__33196\,
            I => \N__33189\
        );

    \I__6253\ : InMux
    port map (
            O => \N__33195\,
            I => \N__33184\
        );

    \I__6252\ : InMux
    port map (
            O => \N__33192\,
            I => \N__33184\
        );

    \I__6251\ : LocalMux
    port map (
            O => \N__33189\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__33184\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__6249\ : InMux
    port map (
            O => \N__33179\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\
        );

    \I__6248\ : CascadeMux
    port map (
            O => \N__33176\,
            I => \N__33171\
        );

    \I__6247\ : InMux
    port map (
            O => \N__33175\,
            I => \N__33168\
        );

    \I__6246\ : InMux
    port map (
            O => \N__33174\,
            I => \N__33163\
        );

    \I__6245\ : InMux
    port map (
            O => \N__33171\,
            I => \N__33163\
        );

    \I__6244\ : LocalMux
    port map (
            O => \N__33168\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__6243\ : LocalMux
    port map (
            O => \N__33163\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__6242\ : InMux
    port map (
            O => \N__33158\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\
        );

    \I__6241\ : InMux
    port map (
            O => \N__33155\,
            I => \N__33148\
        );

    \I__6240\ : InMux
    port map (
            O => \N__33154\,
            I => \N__33148\
        );

    \I__6239\ : InMux
    port map (
            O => \N__33153\,
            I => \N__33145\
        );

    \I__6238\ : LocalMux
    port map (
            O => \N__33148\,
            I => \N__33142\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__33145\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__6236\ : Odrv4
    port map (
            O => \N__33142\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__6235\ : InMux
    port map (
            O => \N__33137\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\
        );

    \I__6234\ : InMux
    port map (
            O => \N__33134\,
            I => \N__33127\
        );

    \I__6233\ : InMux
    port map (
            O => \N__33133\,
            I => \N__33127\
        );

    \I__6232\ : InMux
    port map (
            O => \N__33132\,
            I => \N__33124\
        );

    \I__6231\ : LocalMux
    port map (
            O => \N__33127\,
            I => \N__33121\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__33124\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__6229\ : Odrv4
    port map (
            O => \N__33121\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__6228\ : InMux
    port map (
            O => \N__33116\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\
        );

    \I__6227\ : CascadeMux
    port map (
            O => \N__33113\,
            I => \N__33108\
        );

    \I__6226\ : InMux
    port map (
            O => \N__33112\,
            I => \N__33105\
        );

    \I__6225\ : InMux
    port map (
            O => \N__33111\,
            I => \N__33102\
        );

    \I__6224\ : InMux
    port map (
            O => \N__33108\,
            I => \N__33099\
        );

    \I__6223\ : LocalMux
    port map (
            O => \N__33105\,
            I => \N__33096\
        );

    \I__6222\ : LocalMux
    port map (
            O => \N__33102\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__6221\ : LocalMux
    port map (
            O => \N__33099\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__6220\ : Odrv4
    port map (
            O => \N__33096\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__6219\ : InMux
    port map (
            O => \N__33089\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\
        );

    \I__6218\ : InMux
    port map (
            O => \N__33086\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\
        );

    \I__6217\ : CascadeMux
    port map (
            O => \N__33083\,
            I => \N__33080\
        );

    \I__6216\ : InMux
    port map (
            O => \N__33080\,
            I => \N__33075\
        );

    \I__6215\ : InMux
    port map (
            O => \N__33079\,
            I => \N__33072\
        );

    \I__6214\ : InMux
    port map (
            O => \N__33078\,
            I => \N__33069\
        );

    \I__6213\ : LocalMux
    port map (
            O => \N__33075\,
            I => \N__33066\
        );

    \I__6212\ : LocalMux
    port map (
            O => \N__33072\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__6211\ : LocalMux
    port map (
            O => \N__33069\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__6210\ : Odrv4
    port map (
            O => \N__33066\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__6209\ : InMux
    port map (
            O => \N__33059\,
            I => \N__33056\
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__33056\,
            I => \N__33052\
        );

    \I__6207\ : InMux
    port map (
            O => \N__33055\,
            I => \N__33049\
        );

    \I__6206\ : Span4Mux_h
    port map (
            O => \N__33052\,
            I => \N__33046\
        );

    \I__6205\ : LocalMux
    port map (
            O => \N__33049\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13\
        );

    \I__6204\ : Odrv4
    port map (
            O => \N__33046\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13\
        );

    \I__6203\ : InMux
    port map (
            O => \N__33041\,
            I => \N__33038\
        );

    \I__6202\ : LocalMux
    port map (
            O => \N__33038\,
            I => \N__33033\
        );

    \I__6201\ : InMux
    port map (
            O => \N__33037\,
            I => \N__33028\
        );

    \I__6200\ : InMux
    port map (
            O => \N__33036\,
            I => \N__33028\
        );

    \I__6199\ : Span4Mux_h
    port map (
            O => \N__33033\,
            I => \N__33023\
        );

    \I__6198\ : LocalMux
    port map (
            O => \N__33028\,
            I => \N__33023\
        );

    \I__6197\ : Span4Mux_v
    port map (
            O => \N__33023\,
            I => \N__33019\
        );

    \I__6196\ : InMux
    port map (
            O => \N__33022\,
            I => \N__33016\
        );

    \I__6195\ : Odrv4
    port map (
            O => \N__33019\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__6194\ : LocalMux
    port map (
            O => \N__33016\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__6193\ : CascadeMux
    port map (
            O => \N__33011\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13_cascade_\
        );

    \I__6192\ : CascadeMux
    port map (
            O => \N__33008\,
            I => \N__33005\
        );

    \I__6191\ : InMux
    port map (
            O => \N__33005\,
            I => \N__33002\
        );

    \I__6190\ : LocalMux
    port map (
            O => \N__33002\,
            I => \N__32999\
        );

    \I__6189\ : Odrv4
    port map (
            O => \N__32999\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\
        );

    \I__6188\ : InMux
    port map (
            O => \N__32996\,
            I => \bfn_12_9_0_\
        );

    \I__6187\ : CascadeMux
    port map (
            O => \N__32993\,
            I => \N__32989\
        );

    \I__6186\ : CascadeMux
    port map (
            O => \N__32992\,
            I => \N__32986\
        );

    \I__6185\ : InMux
    port map (
            O => \N__32989\,
            I => \N__32980\
        );

    \I__6184\ : InMux
    port map (
            O => \N__32986\,
            I => \N__32980\
        );

    \I__6183\ : InMux
    port map (
            O => \N__32985\,
            I => \N__32977\
        );

    \I__6182\ : LocalMux
    port map (
            O => \N__32980\,
            I => \N__32974\
        );

    \I__6181\ : LocalMux
    port map (
            O => \N__32977\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__6180\ : Odrv12
    port map (
            O => \N__32974\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__6179\ : InMux
    port map (
            O => \N__32969\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\
        );

    \I__6178\ : InMux
    port map (
            O => \N__32966\,
            I => \N__32959\
        );

    \I__6177\ : InMux
    port map (
            O => \N__32965\,
            I => \N__32959\
        );

    \I__6176\ : InMux
    port map (
            O => \N__32964\,
            I => \N__32956\
        );

    \I__6175\ : LocalMux
    port map (
            O => \N__32959\,
            I => \N__32953\
        );

    \I__6174\ : LocalMux
    port map (
            O => \N__32956\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__6173\ : Odrv4
    port map (
            O => \N__32953\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__6172\ : InMux
    port map (
            O => \N__32948\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\
        );

    \I__6171\ : CascadeMux
    port map (
            O => \N__32945\,
            I => \N__32941\
        );

    \I__6170\ : InMux
    port map (
            O => \N__32944\,
            I => \N__32935\
        );

    \I__6169\ : InMux
    port map (
            O => \N__32941\,
            I => \N__32935\
        );

    \I__6168\ : InMux
    port map (
            O => \N__32940\,
            I => \N__32932\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__32935\,
            I => \N__32929\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__32932\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__6165\ : Odrv12
    port map (
            O => \N__32929\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__6164\ : InMux
    port map (
            O => \N__32924\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\
        );

    \I__6163\ : InMux
    port map (
            O => \N__32921\,
            I => \N__32914\
        );

    \I__6162\ : InMux
    port map (
            O => \N__32920\,
            I => \N__32914\
        );

    \I__6161\ : InMux
    port map (
            O => \N__32919\,
            I => \N__32911\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__32914\,
            I => \N__32908\
        );

    \I__6159\ : LocalMux
    port map (
            O => \N__32911\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__6158\ : Odrv4
    port map (
            O => \N__32908\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__6157\ : InMux
    port map (
            O => \N__32903\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__6156\ : InMux
    port map (
            O => \N__32900\,
            I => \N__32893\
        );

    \I__6155\ : InMux
    port map (
            O => \N__32899\,
            I => \N__32893\
        );

    \I__6154\ : InMux
    port map (
            O => \N__32898\,
            I => \N__32890\
        );

    \I__6153\ : LocalMux
    port map (
            O => \N__32893\,
            I => \N__32887\
        );

    \I__6152\ : LocalMux
    port map (
            O => \N__32890\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__6151\ : Odrv4
    port map (
            O => \N__32887\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__6150\ : InMux
    port map (
            O => \N__32882\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\
        );

    \I__6149\ : InMux
    port map (
            O => \N__32879\,
            I => \N__32872\
        );

    \I__6148\ : InMux
    port map (
            O => \N__32878\,
            I => \N__32872\
        );

    \I__6147\ : InMux
    port map (
            O => \N__32877\,
            I => \N__32869\
        );

    \I__6146\ : LocalMux
    port map (
            O => \N__32872\,
            I => \N__32866\
        );

    \I__6145\ : LocalMux
    port map (
            O => \N__32869\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__6144\ : Odrv4
    port map (
            O => \N__32866\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__6143\ : InMux
    port map (
            O => \N__32861\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\
        );

    \I__6142\ : InMux
    port map (
            O => \N__32858\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\
        );

    \I__6141\ : InMux
    port map (
            O => \N__32855\,
            I => \bfn_12_10_0_\
        );

    \I__6140\ : InMux
    port map (
            O => \N__32852\,
            I => \N__32848\
        );

    \I__6139\ : InMux
    port map (
            O => \N__32851\,
            I => \N__32845\
        );

    \I__6138\ : LocalMux
    port map (
            O => \N__32848\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__6137\ : LocalMux
    port map (
            O => \N__32845\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__6136\ : InMux
    port map (
            O => \N__32840\,
            I => \bfn_12_8_0_\
        );

    \I__6135\ : InMux
    port map (
            O => \N__32837\,
            I => \N__32833\
        );

    \I__6134\ : InMux
    port map (
            O => \N__32836\,
            I => \N__32830\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__32833\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__32830\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__6131\ : InMux
    port map (
            O => \N__32825\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\
        );

    \I__6130\ : InMux
    port map (
            O => \N__32822\,
            I => \N__32818\
        );

    \I__6129\ : InMux
    port map (
            O => \N__32821\,
            I => \N__32815\
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__32818\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__6127\ : LocalMux
    port map (
            O => \N__32815\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__6126\ : InMux
    port map (
            O => \N__32810\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\
        );

    \I__6125\ : InMux
    port map (
            O => \N__32807\,
            I => \N__32803\
        );

    \I__6124\ : InMux
    port map (
            O => \N__32806\,
            I => \N__32800\
        );

    \I__6123\ : LocalMux
    port map (
            O => \N__32803\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__32800\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__6121\ : InMux
    port map (
            O => \N__32795\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\
        );

    \I__6120\ : InMux
    port map (
            O => \N__32792\,
            I => \N__32788\
        );

    \I__6119\ : InMux
    port map (
            O => \N__32791\,
            I => \N__32785\
        );

    \I__6118\ : LocalMux
    port map (
            O => \N__32788\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__32785\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__6116\ : InMux
    port map (
            O => \N__32780\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\
        );

    \I__6115\ : InMux
    port map (
            O => \N__32777\,
            I => \N__32773\
        );

    \I__6114\ : InMux
    port map (
            O => \N__32776\,
            I => \N__32770\
        );

    \I__6113\ : LocalMux
    port map (
            O => \N__32773\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__6112\ : LocalMux
    port map (
            O => \N__32770\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__6111\ : InMux
    port map (
            O => \N__32765\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\
        );

    \I__6110\ : InMux
    port map (
            O => \N__32762\,
            I => \N__32758\
        );

    \I__6109\ : InMux
    port map (
            O => \N__32761\,
            I => \N__32755\
        );

    \I__6108\ : LocalMux
    port map (
            O => \N__32758\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__32755\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__6106\ : InMux
    port map (
            O => \N__32750\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\
        );

    \I__6105\ : InMux
    port map (
            O => \N__32747\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\
        );

    \I__6104\ : InMux
    port map (
            O => \N__32744\,
            I => \N__32741\
        );

    \I__6103\ : LocalMux
    port map (
            O => \N__32741\,
            I => \N__32738\
        );

    \I__6102\ : Span4Mux_h
    port map (
            O => \N__32738\,
            I => \N__32734\
        );

    \I__6101\ : InMux
    port map (
            O => \N__32737\,
            I => \N__32730\
        );

    \I__6100\ : Span4Mux_v
    port map (
            O => \N__32734\,
            I => \N__32727\
        );

    \I__6099\ : InMux
    port map (
            O => \N__32733\,
            I => \N__32724\
        );

    \I__6098\ : LocalMux
    port map (
            O => \N__32730\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__6097\ : Odrv4
    port map (
            O => \N__32727\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__6096\ : LocalMux
    port map (
            O => \N__32724\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__6095\ : InMux
    port map (
            O => \N__32717\,
            I => \N__32714\
        );

    \I__6094\ : LocalMux
    port map (
            O => \N__32714\,
            I => \N__32709\
        );

    \I__6093\ : InMux
    port map (
            O => \N__32713\,
            I => \N__32706\
        );

    \I__6092\ : InMux
    port map (
            O => \N__32712\,
            I => \N__32703\
        );

    \I__6091\ : Span4Mux_v
    port map (
            O => \N__32709\,
            I => \N__32700\
        );

    \I__6090\ : LocalMux
    port map (
            O => \N__32706\,
            I => \N__32697\
        );

    \I__6089\ : LocalMux
    port map (
            O => \N__32703\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__6088\ : Odrv4
    port map (
            O => \N__32700\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__6087\ : Odrv12
    port map (
            O => \N__32697\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__6086\ : CascadeMux
    port map (
            O => \N__32690\,
            I => \N__32687\
        );

    \I__6085\ : InMux
    port map (
            O => \N__32687\,
            I => \N__32684\
        );

    \I__6084\ : LocalMux
    port map (
            O => \N__32684\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\
        );

    \I__6083\ : InMux
    port map (
            O => \N__32681\,
            I => \N__32677\
        );

    \I__6082\ : InMux
    port map (
            O => \N__32680\,
            I => \N__32674\
        );

    \I__6081\ : LocalMux
    port map (
            O => \N__32677\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__6080\ : LocalMux
    port map (
            O => \N__32674\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__6079\ : InMux
    port map (
            O => \N__32669\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\
        );

    \I__6078\ : CascadeMux
    port map (
            O => \N__32666\,
            I => \N__32663\
        );

    \I__6077\ : InMux
    port map (
            O => \N__32663\,
            I => \N__32659\
        );

    \I__6076\ : InMux
    port map (
            O => \N__32662\,
            I => \N__32656\
        );

    \I__6075\ : LocalMux
    port map (
            O => \N__32659\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__6074\ : LocalMux
    port map (
            O => \N__32656\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__6073\ : InMux
    port map (
            O => \N__32651\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\
        );

    \I__6072\ : InMux
    port map (
            O => \N__32648\,
            I => \N__32644\
        );

    \I__6071\ : InMux
    port map (
            O => \N__32647\,
            I => \N__32641\
        );

    \I__6070\ : LocalMux
    port map (
            O => \N__32644\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__6069\ : LocalMux
    port map (
            O => \N__32641\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__6068\ : InMux
    port map (
            O => \N__32636\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\
        );

    \I__6067\ : InMux
    port map (
            O => \N__32633\,
            I => \N__32629\
        );

    \I__6066\ : InMux
    port map (
            O => \N__32632\,
            I => \N__32626\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__32629\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__6064\ : LocalMux
    port map (
            O => \N__32626\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__6063\ : InMux
    port map (
            O => \N__32621\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\
        );

    \I__6062\ : InMux
    port map (
            O => \N__32618\,
            I => \N__32614\
        );

    \I__6061\ : InMux
    port map (
            O => \N__32617\,
            I => \N__32611\
        );

    \I__6060\ : LocalMux
    port map (
            O => \N__32614\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__6059\ : LocalMux
    port map (
            O => \N__32611\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__6058\ : InMux
    port map (
            O => \N__32606\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\
        );

    \I__6057\ : InMux
    port map (
            O => \N__32603\,
            I => \N__32599\
        );

    \I__6056\ : InMux
    port map (
            O => \N__32602\,
            I => \N__32596\
        );

    \I__6055\ : LocalMux
    port map (
            O => \N__32599\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__6054\ : LocalMux
    port map (
            O => \N__32596\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__6053\ : InMux
    port map (
            O => \N__32591\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\
        );

    \I__6052\ : InMux
    port map (
            O => \N__32588\,
            I => \N__32584\
        );

    \I__6051\ : InMux
    port map (
            O => \N__32587\,
            I => \N__32581\
        );

    \I__6050\ : LocalMux
    port map (
            O => \N__32584\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__6049\ : LocalMux
    port map (
            O => \N__32581\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__6048\ : InMux
    port map (
            O => \N__32576\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\
        );

    \I__6047\ : InMux
    port map (
            O => \N__32573\,
            I => \N__32570\
        );

    \I__6046\ : LocalMux
    port map (
            O => \N__32570\,
            I => \N__32567\
        );

    \I__6045\ : Odrv4
    port map (
            O => \N__32567\,
            I => \current_shift_inst.control_input_axb_18\
        );

    \I__6044\ : InMux
    port map (
            O => \N__32564\,
            I => \N__32561\
        );

    \I__6043\ : LocalMux
    port map (
            O => \N__32561\,
            I => \N__32558\
        );

    \I__6042\ : Odrv4
    port map (
            O => \N__32558\,
            I => \current_shift_inst.control_input_axb_17\
        );

    \I__6041\ : InMux
    port map (
            O => \N__32555\,
            I => \N__32552\
        );

    \I__6040\ : LocalMux
    port map (
            O => \N__32552\,
            I => \N__32548\
        );

    \I__6039\ : InMux
    port map (
            O => \N__32551\,
            I => \N__32545\
        );

    \I__6038\ : Span4Mux_h
    port map (
            O => \N__32548\,
            I => \N__32542\
        );

    \I__6037\ : LocalMux
    port map (
            O => \N__32545\,
            I => \N__32539\
        );

    \I__6036\ : Sp12to4
    port map (
            O => \N__32542\,
            I => \N__32536\
        );

    \I__6035\ : Span12Mux_v
    port map (
            O => \N__32539\,
            I => \N__32533\
        );

    \I__6034\ : Span12Mux_s6_v
    port map (
            O => \N__32536\,
            I => \N__32530\
        );

    \I__6033\ : Span12Mux_h
    port map (
            O => \N__32533\,
            I => \N__32527\
        );

    \I__6032\ : Odrv12
    port map (
            O => \N__32530\,
            I => \pwm_generator_inst.un2_threshold_2_1_15\
        );

    \I__6031\ : Odrv12
    port map (
            O => \N__32527\,
            I => \pwm_generator_inst.un2_threshold_2_1_15\
        );

    \I__6030\ : InMux
    port map (
            O => \N__32522\,
            I => \N__32518\
        );

    \I__6029\ : InMux
    port map (
            O => \N__32521\,
            I => \N__32515\
        );

    \I__6028\ : LocalMux
    port map (
            O => \N__32518\,
            I => \N__32510\
        );

    \I__6027\ : LocalMux
    port map (
            O => \N__32515\,
            I => \N__32510\
        );

    \I__6026\ : Span4Mux_h
    port map (
            O => \N__32510\,
            I => \N__32507\
        );

    \I__6025\ : Span4Mux_v
    port map (
            O => \N__32507\,
            I => \N__32498\
        );

    \I__6024\ : InMux
    port map (
            O => \N__32506\,
            I => \N__32491\
        );

    \I__6023\ : InMux
    port map (
            O => \N__32505\,
            I => \N__32491\
        );

    \I__6022\ : InMux
    port map (
            O => \N__32504\,
            I => \N__32491\
        );

    \I__6021\ : InMux
    port map (
            O => \N__32503\,
            I => \N__32484\
        );

    \I__6020\ : InMux
    port map (
            O => \N__32502\,
            I => \N__32484\
        );

    \I__6019\ : InMux
    port map (
            O => \N__32501\,
            I => \N__32484\
        );

    \I__6018\ : Sp12to4
    port map (
            O => \N__32498\,
            I => \N__32477\
        );

    \I__6017\ : LocalMux
    port map (
            O => \N__32491\,
            I => \N__32477\
        );

    \I__6016\ : LocalMux
    port map (
            O => \N__32484\,
            I => \N__32477\
        );

    \I__6015\ : Span12Mux_h
    port map (
            O => \N__32477\,
            I => \N__32474\
        );

    \I__6014\ : Odrv12
    port map (
            O => \N__32474\,
            I => \pwm_generator_inst.un2_threshold_1_25\
        );

    \I__6013\ : InMux
    port map (
            O => \N__32471\,
            I => \N__32440\
        );

    \I__6012\ : InMux
    port map (
            O => \N__32470\,
            I => \N__32440\
        );

    \I__6011\ : InMux
    port map (
            O => \N__32469\,
            I => \N__32440\
        );

    \I__6010\ : InMux
    port map (
            O => \N__32468\,
            I => \N__32440\
        );

    \I__6009\ : InMux
    port map (
            O => \N__32467\,
            I => \N__32440\
        );

    \I__6008\ : InMux
    port map (
            O => \N__32466\,
            I => \N__32440\
        );

    \I__6007\ : InMux
    port map (
            O => \N__32465\,
            I => \N__32440\
        );

    \I__6006\ : InMux
    port map (
            O => \N__32464\,
            I => \N__32440\
        );

    \I__6005\ : InMux
    port map (
            O => \N__32463\,
            I => \N__32425\
        );

    \I__6004\ : InMux
    port map (
            O => \N__32462\,
            I => \N__32425\
        );

    \I__6003\ : InMux
    port map (
            O => \N__32461\,
            I => \N__32425\
        );

    \I__6002\ : InMux
    port map (
            O => \N__32460\,
            I => \N__32425\
        );

    \I__6001\ : InMux
    port map (
            O => \N__32459\,
            I => \N__32425\
        );

    \I__6000\ : InMux
    port map (
            O => \N__32458\,
            I => \N__32425\
        );

    \I__5999\ : InMux
    port map (
            O => \N__32457\,
            I => \N__32425\
        );

    \I__5998\ : LocalMux
    port map (
            O => \N__32440\,
            I => \N__32418\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__32425\,
            I => \N__32418\
        );

    \I__5996\ : InMux
    port map (
            O => \N__32424\,
            I => \N__32415\
        );

    \I__5995\ : InMux
    port map (
            O => \N__32423\,
            I => \N__32412\
        );

    \I__5994\ : Span4Mux_s3_h
    port map (
            O => \N__32418\,
            I => \N__32403\
        );

    \I__5993\ : LocalMux
    port map (
            O => \N__32415\,
            I => \N__32400\
        );

    \I__5992\ : LocalMux
    port map (
            O => \N__32412\,
            I => \N__32397\
        );

    \I__5991\ : CascadeMux
    port map (
            O => \N__32411\,
            I => \N__32386\
        );

    \I__5990\ : InMux
    port map (
            O => \N__32410\,
            I => \N__32381\
        );

    \I__5989\ : InMux
    port map (
            O => \N__32409\,
            I => \N__32381\
        );

    \I__5988\ : InMux
    port map (
            O => \N__32408\,
            I => \N__32374\
        );

    \I__5987\ : InMux
    port map (
            O => \N__32407\,
            I => \N__32374\
        );

    \I__5986\ : InMux
    port map (
            O => \N__32406\,
            I => \N__32374\
        );

    \I__5985\ : Span4Mux_h
    port map (
            O => \N__32403\,
            I => \N__32371\
        );

    \I__5984\ : Span4Mux_v
    port map (
            O => \N__32400\,
            I => \N__32368\
        );

    \I__5983\ : Span4Mux_v
    port map (
            O => \N__32397\,
            I => \N__32364\
        );

    \I__5982\ : InMux
    port map (
            O => \N__32396\,
            I => \N__32347\
        );

    \I__5981\ : InMux
    port map (
            O => \N__32395\,
            I => \N__32347\
        );

    \I__5980\ : InMux
    port map (
            O => \N__32394\,
            I => \N__32347\
        );

    \I__5979\ : InMux
    port map (
            O => \N__32393\,
            I => \N__32347\
        );

    \I__5978\ : InMux
    port map (
            O => \N__32392\,
            I => \N__32347\
        );

    \I__5977\ : InMux
    port map (
            O => \N__32391\,
            I => \N__32347\
        );

    \I__5976\ : InMux
    port map (
            O => \N__32390\,
            I => \N__32347\
        );

    \I__5975\ : InMux
    port map (
            O => \N__32389\,
            I => \N__32347\
        );

    \I__5974\ : InMux
    port map (
            O => \N__32386\,
            I => \N__32344\
        );

    \I__5973\ : LocalMux
    port map (
            O => \N__32381\,
            I => \N__32339\
        );

    \I__5972\ : LocalMux
    port map (
            O => \N__32374\,
            I => \N__32339\
        );

    \I__5971\ : Span4Mux_h
    port map (
            O => \N__32371\,
            I => \N__32336\
        );

    \I__5970\ : Span4Mux_h
    port map (
            O => \N__32368\,
            I => \N__32333\
        );

    \I__5969\ : InMux
    port map (
            O => \N__32367\,
            I => \N__32330\
        );

    \I__5968\ : Sp12to4
    port map (
            O => \N__32364\,
            I => \N__32321\
        );

    \I__5967\ : LocalMux
    port map (
            O => \N__32347\,
            I => \N__32321\
        );

    \I__5966\ : LocalMux
    port map (
            O => \N__32344\,
            I => \N__32321\
        );

    \I__5965\ : Span12Mux_s7_v
    port map (
            O => \N__32339\,
            I => \N__32321\
        );

    \I__5964\ : Span4Mux_h
    port map (
            O => \N__32336\,
            I => \N__32318\
        );

    \I__5963\ : Odrv4
    port map (
            O => \N__32333\,
            I => \N_19_1\
        );

    \I__5962\ : LocalMux
    port map (
            O => \N__32330\,
            I => \N_19_1\
        );

    \I__5961\ : Odrv12
    port map (
            O => \N__32321\,
            I => \N_19_1\
        );

    \I__5960\ : Odrv4
    port map (
            O => \N__32318\,
            I => \N_19_1\
        );

    \I__5959\ : InMux
    port map (
            O => \N__32309\,
            I => \N__32306\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__32306\,
            I => \N__32303\
        );

    \I__5957\ : Span4Mux_v
    port map (
            O => \N__32303\,
            I => \N__32300\
        );

    \I__5956\ : Sp12to4
    port map (
            O => \N__32300\,
            I => \N__32297\
        );

    \I__5955\ : Span12Mux_h
    port map (
            O => \N__32297\,
            I => \N__32294\
        );

    \I__5954\ : Odrv12
    port map (
            O => \N__32294\,
            I => \pwm_generator_inst.un2_threshold_2_1_16\
        );

    \I__5953\ : InMux
    port map (
            O => \N__32291\,
            I => \N__32288\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__32288\,
            I => \N__32285\
        );

    \I__5951\ : Span4Mux_v
    port map (
            O => \N__32285\,
            I => \N__32282\
        );

    \I__5950\ : Odrv4
    port map (
            O => \N__32282\,
            I => \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\
        );

    \I__5949\ : InMux
    port map (
            O => \N__32279\,
            I => \N__32276\
        );

    \I__5948\ : LocalMux
    port map (
            O => \N__32276\,
            I => \N__32273\
        );

    \I__5947\ : Span4Mux_v
    port map (
            O => \N__32273\,
            I => \N__32270\
        );

    \I__5946\ : Span4Mux_h
    port map (
            O => \N__32270\,
            I => \N__32267\
        );

    \I__5945\ : Odrv4
    port map (
            O => \N__32267\,
            I => il_max_comp1_c
        );

    \I__5944\ : InMux
    port map (
            O => \N__32264\,
            I => \N__32261\
        );

    \I__5943\ : LocalMux
    port map (
            O => \N__32261\,
            I => \il_max_comp1_D1\
        );

    \I__5942\ : InMux
    port map (
            O => \N__32258\,
            I => \N__32254\
        );

    \I__5941\ : InMux
    port map (
            O => \N__32257\,
            I => \N__32250\
        );

    \I__5940\ : LocalMux
    port map (
            O => \N__32254\,
            I => \N__32247\
        );

    \I__5939\ : InMux
    port map (
            O => \N__32253\,
            I => \N__32244\
        );

    \I__5938\ : LocalMux
    port map (
            O => \N__32250\,
            I => \N__32240\
        );

    \I__5937\ : Span4Mux_h
    port map (
            O => \N__32247\,
            I => \N__32235\
        );

    \I__5936\ : LocalMux
    port map (
            O => \N__32244\,
            I => \N__32235\
        );

    \I__5935\ : InMux
    port map (
            O => \N__32243\,
            I => \N__32232\
        );

    \I__5934\ : Span4Mux_v
    port map (
            O => \N__32240\,
            I => \N__32229\
        );

    \I__5933\ : Span4Mux_v
    port map (
            O => \N__32235\,
            I => \N__32226\
        );

    \I__5932\ : LocalMux
    port map (
            O => \N__32232\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__5931\ : Odrv4
    port map (
            O => \N__32229\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__5930\ : Odrv4
    port map (
            O => \N__32226\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__5929\ : InMux
    port map (
            O => \N__32219\,
            I => \N__32216\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__32216\,
            I => \N__32212\
        );

    \I__5927\ : InMux
    port map (
            O => \N__32215\,
            I => \N__32209\
        );

    \I__5926\ : Span4Mux_v
    port map (
            O => \N__32212\,
            I => \N__32205\
        );

    \I__5925\ : LocalMux
    port map (
            O => \N__32209\,
            I => \N__32202\
        );

    \I__5924\ : InMux
    port map (
            O => \N__32208\,
            I => \N__32199\
        );

    \I__5923\ : Span4Mux_h
    port map (
            O => \N__32205\,
            I => \N__32196\
        );

    \I__5922\ : Span4Mux_v
    port map (
            O => \N__32202\,
            I => \N__32193\
        );

    \I__5921\ : LocalMux
    port map (
            O => \N__32199\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__5920\ : Odrv4
    port map (
            O => \N__32196\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__5919\ : Odrv4
    port map (
            O => \N__32193\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__5918\ : InMux
    port map (
            O => \N__32186\,
            I => \N__32183\
        );

    \I__5917\ : LocalMux
    port map (
            O => \N__32183\,
            I => \N__32180\
        );

    \I__5916\ : Span4Mux_v
    port map (
            O => \N__32180\,
            I => \N__32175\
        );

    \I__5915\ : InMux
    port map (
            O => \N__32179\,
            I => \N__32172\
        );

    \I__5914\ : InMux
    port map (
            O => \N__32178\,
            I => \N__32169\
        );

    \I__5913\ : Span4Mux_v
    port map (
            O => \N__32175\,
            I => \N__32165\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__32172\,
            I => \N__32160\
        );

    \I__5911\ : LocalMux
    port map (
            O => \N__32169\,
            I => \N__32160\
        );

    \I__5910\ : InMux
    port map (
            O => \N__32168\,
            I => \N__32157\
        );

    \I__5909\ : Odrv4
    port map (
            O => \N__32165\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__5908\ : Odrv12
    port map (
            O => \N__32160\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__5907\ : LocalMux
    port map (
            O => \N__32157\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__5906\ : InMux
    port map (
            O => \N__32150\,
            I => \N__32147\
        );

    \I__5905\ : LocalMux
    port map (
            O => \N__32147\,
            I => \N__32144\
        );

    \I__5904\ : Odrv4
    port map (
            O => \N__32144\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24\
        );

    \I__5903\ : InMux
    port map (
            O => \N__32141\,
            I => \bfn_11_18_0_\
        );

    \I__5902\ : CascadeMux
    port map (
            O => \N__32138\,
            I => \N__32135\
        );

    \I__5901\ : InMux
    port map (
            O => \N__32135\,
            I => \N__32132\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__32132\,
            I => \N__32129\
        );

    \I__5899\ : Odrv4
    port map (
            O => \N__32129\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25\
        );

    \I__5898\ : InMux
    port map (
            O => \N__32126\,
            I => \current_shift_inst.control_input_cry_24\
        );

    \I__5897\ : InMux
    port map (
            O => \N__32123\,
            I => \N__32120\
        );

    \I__5896\ : LocalMux
    port map (
            O => \N__32120\,
            I => \N__32117\
        );

    \I__5895\ : Odrv4
    port map (
            O => \N__32117\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26\
        );

    \I__5894\ : InMux
    port map (
            O => \N__32114\,
            I => \current_shift_inst.control_input_cry_25\
        );

    \I__5893\ : InMux
    port map (
            O => \N__32111\,
            I => \N__32108\
        );

    \I__5892\ : LocalMux
    port map (
            O => \N__32108\,
            I => \N__32105\
        );

    \I__5891\ : Odrv4
    port map (
            O => \N__32105\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27\
        );

    \I__5890\ : InMux
    port map (
            O => \N__32102\,
            I => \current_shift_inst.control_input_cry_26\
        );

    \I__5889\ : CascadeMux
    port map (
            O => \N__32099\,
            I => \N__32096\
        );

    \I__5888\ : InMux
    port map (
            O => \N__32096\,
            I => \N__32093\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__32093\,
            I => \N__32090\
        );

    \I__5886\ : Odrv4
    port map (
            O => \N__32090\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28\
        );

    \I__5885\ : InMux
    port map (
            O => \N__32087\,
            I => \current_shift_inst.control_input_cry_27\
        );

    \I__5884\ : InMux
    port map (
            O => \N__32084\,
            I => \N__32081\
        );

    \I__5883\ : LocalMux
    port map (
            O => \N__32081\,
            I => \N__32078\
        );

    \I__5882\ : Odrv4
    port map (
            O => \N__32078\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29\
        );

    \I__5881\ : InMux
    port map (
            O => \N__32075\,
            I => \current_shift_inst.control_input_cry_28\
        );

    \I__5880\ : InMux
    port map (
            O => \N__32072\,
            I => \current_shift_inst.control_input_cry_29\
        );

    \I__5879\ : InMux
    port map (
            O => \N__32069\,
            I => \N__32066\
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__32066\,
            I => \N__32062\
        );

    \I__5877\ : InMux
    port map (
            O => \N__32065\,
            I => \N__32059\
        );

    \I__5876\ : Odrv4
    port map (
            O => \N__32062\,
            I => \current_shift_inst.control_input_31\
        );

    \I__5875\ : LocalMux
    port map (
            O => \N__32059\,
            I => \current_shift_inst.control_input_31\
        );

    \I__5874\ : InMux
    port map (
            O => \N__32054\,
            I => \N__32051\
        );

    \I__5873\ : LocalMux
    port map (
            O => \N__32051\,
            I => \current_shift_inst.control_input_axb_27\
        );

    \I__5872\ : CascadeMux
    port map (
            O => \N__32048\,
            I => \N__32045\
        );

    \I__5871\ : InMux
    port map (
            O => \N__32045\,
            I => \N__32042\
        );

    \I__5870\ : LocalMux
    port map (
            O => \N__32042\,
            I => \N__32039\
        );

    \I__5869\ : Odrv12
    port map (
            O => \N__32039\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16\
        );

    \I__5868\ : InMux
    port map (
            O => \N__32036\,
            I => \bfn_11_17_0_\
        );

    \I__5867\ : CascadeMux
    port map (
            O => \N__32033\,
            I => \N__32030\
        );

    \I__5866\ : InMux
    port map (
            O => \N__32030\,
            I => \N__32027\
        );

    \I__5865\ : LocalMux
    port map (
            O => \N__32027\,
            I => \N__32024\
        );

    \I__5864\ : Odrv4
    port map (
            O => \N__32024\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17\
        );

    \I__5863\ : InMux
    port map (
            O => \N__32021\,
            I => \current_shift_inst.control_input_cry_16\
        );

    \I__5862\ : InMux
    port map (
            O => \N__32018\,
            I => \N__32015\
        );

    \I__5861\ : LocalMux
    port map (
            O => \N__32015\,
            I => \N__32012\
        );

    \I__5860\ : Span4Mux_h
    port map (
            O => \N__32012\,
            I => \N__32009\
        );

    \I__5859\ : Odrv4
    port map (
            O => \N__32009\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18\
        );

    \I__5858\ : InMux
    port map (
            O => \N__32006\,
            I => \current_shift_inst.control_input_cry_17\
        );

    \I__5857\ : InMux
    port map (
            O => \N__32003\,
            I => \N__32000\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__32000\,
            I => \current_shift_inst.control_input_axb_19\
        );

    \I__5855\ : InMux
    port map (
            O => \N__31997\,
            I => \N__31994\
        );

    \I__5854\ : LocalMux
    port map (
            O => \N__31994\,
            I => \N__31991\
        );

    \I__5853\ : Odrv4
    port map (
            O => \N__31991\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19\
        );

    \I__5852\ : InMux
    port map (
            O => \N__31988\,
            I => \current_shift_inst.control_input_cry_18\
        );

    \I__5851\ : InMux
    port map (
            O => \N__31985\,
            I => \N__31982\
        );

    \I__5850\ : LocalMux
    port map (
            O => \N__31982\,
            I => \N__31979\
        );

    \I__5849\ : Odrv4
    port map (
            O => \N__31979\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20\
        );

    \I__5848\ : InMux
    port map (
            O => \N__31976\,
            I => \current_shift_inst.control_input_cry_19\
        );

    \I__5847\ : InMux
    port map (
            O => \N__31973\,
            I => \N__31970\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__31970\,
            I => \N__31967\
        );

    \I__5845\ : Odrv4
    port map (
            O => \N__31967\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21\
        );

    \I__5844\ : InMux
    port map (
            O => \N__31964\,
            I => \current_shift_inst.control_input_cry_20\
        );

    \I__5843\ : InMux
    port map (
            O => \N__31961\,
            I => \N__31958\
        );

    \I__5842\ : LocalMux
    port map (
            O => \N__31958\,
            I => \N__31955\
        );

    \I__5841\ : Odrv4
    port map (
            O => \N__31955\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22\
        );

    \I__5840\ : InMux
    port map (
            O => \N__31952\,
            I => \current_shift_inst.control_input_cry_21\
        );

    \I__5839\ : CascadeMux
    port map (
            O => \N__31949\,
            I => \N__31946\
        );

    \I__5838\ : InMux
    port map (
            O => \N__31946\,
            I => \N__31943\
        );

    \I__5837\ : LocalMux
    port map (
            O => \N__31943\,
            I => \N__31940\
        );

    \I__5836\ : Odrv4
    port map (
            O => \N__31940\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23\
        );

    \I__5835\ : InMux
    port map (
            O => \N__31937\,
            I => \current_shift_inst.control_input_cry_22\
        );

    \I__5834\ : InMux
    port map (
            O => \N__31934\,
            I => \N__31931\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__31931\,
            I => \current_shift_inst.control_input_axb_8\
        );

    \I__5832\ : InMux
    port map (
            O => \N__31928\,
            I => \N__31925\
        );

    \I__5831\ : LocalMux
    port map (
            O => \N__31925\,
            I => \N__31922\
        );

    \I__5830\ : Odrv4
    port map (
            O => \N__31922\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\
        );

    \I__5829\ : InMux
    port map (
            O => \N__31919\,
            I => \bfn_11_16_0_\
        );

    \I__5828\ : InMux
    port map (
            O => \N__31916\,
            I => \N__31913\
        );

    \I__5827\ : LocalMux
    port map (
            O => \N__31913\,
            I => \current_shift_inst.control_input_axb_9\
        );

    \I__5826\ : InMux
    port map (
            O => \N__31910\,
            I => \N__31907\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__31907\,
            I => \N__31904\
        );

    \I__5824\ : Odrv4
    port map (
            O => \N__31904\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\
        );

    \I__5823\ : InMux
    port map (
            O => \N__31901\,
            I => \current_shift_inst.control_input_cry_8\
        );

    \I__5822\ : CascadeMux
    port map (
            O => \N__31898\,
            I => \N__31895\
        );

    \I__5821\ : InMux
    port map (
            O => \N__31895\,
            I => \N__31892\
        );

    \I__5820\ : LocalMux
    port map (
            O => \N__31892\,
            I => \current_shift_inst.control_input_axb_10\
        );

    \I__5819\ : InMux
    port map (
            O => \N__31889\,
            I => \N__31886\
        );

    \I__5818\ : LocalMux
    port map (
            O => \N__31886\,
            I => \N__31883\
        );

    \I__5817\ : Span4Mux_h
    port map (
            O => \N__31883\,
            I => \N__31880\
        );

    \I__5816\ : Odrv4
    port map (
            O => \N__31880\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\
        );

    \I__5815\ : InMux
    port map (
            O => \N__31877\,
            I => \current_shift_inst.control_input_cry_9\
        );

    \I__5814\ : InMux
    port map (
            O => \N__31874\,
            I => \N__31871\
        );

    \I__5813\ : LocalMux
    port map (
            O => \N__31871\,
            I => \N__31868\
        );

    \I__5812\ : Odrv4
    port map (
            O => \N__31868\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\
        );

    \I__5811\ : InMux
    port map (
            O => \N__31865\,
            I => \current_shift_inst.control_input_cry_10\
        );

    \I__5810\ : CascadeMux
    port map (
            O => \N__31862\,
            I => \N__31859\
        );

    \I__5809\ : InMux
    port map (
            O => \N__31859\,
            I => \N__31856\
        );

    \I__5808\ : LocalMux
    port map (
            O => \N__31856\,
            I => \N__31853\
        );

    \I__5807\ : Odrv4
    port map (
            O => \N__31853\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\
        );

    \I__5806\ : InMux
    port map (
            O => \N__31850\,
            I => \current_shift_inst.control_input_cry_11\
        );

    \I__5805\ : CascadeMux
    port map (
            O => \N__31847\,
            I => \N__31844\
        );

    \I__5804\ : InMux
    port map (
            O => \N__31844\,
            I => \N__31841\
        );

    \I__5803\ : LocalMux
    port map (
            O => \N__31841\,
            I => \N__31838\
        );

    \I__5802\ : Odrv4
    port map (
            O => \N__31838\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\
        );

    \I__5801\ : InMux
    port map (
            O => \N__31835\,
            I => \current_shift_inst.control_input_cry_12\
        );

    \I__5800\ : CascadeMux
    port map (
            O => \N__31832\,
            I => \N__31829\
        );

    \I__5799\ : InMux
    port map (
            O => \N__31829\,
            I => \N__31826\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__31826\,
            I => \N__31823\
        );

    \I__5797\ : Odrv4
    port map (
            O => \N__31823\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14\
        );

    \I__5796\ : InMux
    port map (
            O => \N__31820\,
            I => \current_shift_inst.control_input_cry_13\
        );

    \I__5795\ : CascadeMux
    port map (
            O => \N__31817\,
            I => \N__31814\
        );

    \I__5794\ : InMux
    port map (
            O => \N__31814\,
            I => \N__31811\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__31811\,
            I => \N__31808\
        );

    \I__5792\ : Odrv4
    port map (
            O => \N__31808\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15\
        );

    \I__5791\ : InMux
    port map (
            O => \N__31805\,
            I => \current_shift_inst.control_input_cry_14\
        );

    \I__5790\ : IoInMux
    port map (
            O => \N__31802\,
            I => \N__31799\
        );

    \I__5789\ : LocalMux
    port map (
            O => \N__31799\,
            I => \N__31796\
        );

    \I__5788\ : Span4Mux_s3_v
    port map (
            O => \N__31796\,
            I => \N__31793\
        );

    \I__5787\ : Span4Mux_h
    port map (
            O => \N__31793\,
            I => \N__31790\
        );

    \I__5786\ : Sp12to4
    port map (
            O => \N__31790\,
            I => \N__31787\
        );

    \I__5785\ : Span12Mux_v
    port map (
            O => \N__31787\,
            I => \N__31783\
        );

    \I__5784\ : InMux
    port map (
            O => \N__31786\,
            I => \N__31780\
        );

    \I__5783\ : Odrv12
    port map (
            O => \N__31783\,
            I => \T45_c\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__31780\,
            I => \T45_c\
        );

    \I__5781\ : InMux
    port map (
            O => \N__31775\,
            I => \N__31772\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__31772\,
            I => \current_shift_inst.control_input_axb_0\
        );

    \I__5779\ : CascadeMux
    port map (
            O => \N__31769\,
            I => \N__31764\
        );

    \I__5778\ : InMux
    port map (
            O => \N__31768\,
            I => \N__31761\
        );

    \I__5777\ : InMux
    port map (
            O => \N__31767\,
            I => \N__31758\
        );

    \I__5776\ : InMux
    port map (
            O => \N__31764\,
            I => \N__31755\
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__31761\,
            I => \current_shift_inst.N_1269_i\
        );

    \I__5774\ : LocalMux
    port map (
            O => \N__31758\,
            I => \current_shift_inst.N_1269_i\
        );

    \I__5773\ : LocalMux
    port map (
            O => \N__31755\,
            I => \current_shift_inst.N_1269_i\
        );

    \I__5772\ : InMux
    port map (
            O => \N__31748\,
            I => \N__31745\
        );

    \I__5771\ : LocalMux
    port map (
            O => \N__31745\,
            I => \N__31742\
        );

    \I__5770\ : Odrv4
    port map (
            O => \N__31742\,
            I => \current_shift_inst.control_input_1\
        );

    \I__5769\ : InMux
    port map (
            O => \N__31739\,
            I => \N__31736\
        );

    \I__5768\ : LocalMux
    port map (
            O => \N__31736\,
            I => \N__31733\
        );

    \I__5767\ : Odrv4
    port map (
            O => \N__31733\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\
        );

    \I__5766\ : InMux
    port map (
            O => \N__31730\,
            I => \current_shift_inst.control_input_cry_0\
        );

    \I__5765\ : InMux
    port map (
            O => \N__31727\,
            I => \N__31724\
        );

    \I__5764\ : LocalMux
    port map (
            O => \N__31724\,
            I => \N__31721\
        );

    \I__5763\ : Odrv4
    port map (
            O => \N__31721\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\
        );

    \I__5762\ : InMux
    port map (
            O => \N__31718\,
            I => \current_shift_inst.control_input_cry_1\
        );

    \I__5761\ : InMux
    port map (
            O => \N__31715\,
            I => \N__31712\
        );

    \I__5760\ : LocalMux
    port map (
            O => \N__31712\,
            I => \N__31709\
        );

    \I__5759\ : Odrv4
    port map (
            O => \N__31709\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\
        );

    \I__5758\ : InMux
    port map (
            O => \N__31706\,
            I => \current_shift_inst.control_input_cry_2\
        );

    \I__5757\ : InMux
    port map (
            O => \N__31703\,
            I => \N__31700\
        );

    \I__5756\ : LocalMux
    port map (
            O => \N__31700\,
            I => \N__31697\
        );

    \I__5755\ : Odrv4
    port map (
            O => \N__31697\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\
        );

    \I__5754\ : InMux
    port map (
            O => \N__31694\,
            I => \current_shift_inst.control_input_cry_3\
        );

    \I__5753\ : CascadeMux
    port map (
            O => \N__31691\,
            I => \N__31688\
        );

    \I__5752\ : InMux
    port map (
            O => \N__31688\,
            I => \N__31685\
        );

    \I__5751\ : LocalMux
    port map (
            O => \N__31685\,
            I => \N__31682\
        );

    \I__5750\ : Odrv4
    port map (
            O => \N__31682\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\
        );

    \I__5749\ : InMux
    port map (
            O => \N__31679\,
            I => \current_shift_inst.control_input_cry_4\
        );

    \I__5748\ : CascadeMux
    port map (
            O => \N__31676\,
            I => \N__31673\
        );

    \I__5747\ : InMux
    port map (
            O => \N__31673\,
            I => \N__31670\
        );

    \I__5746\ : LocalMux
    port map (
            O => \N__31670\,
            I => \N__31667\
        );

    \I__5745\ : Odrv4
    port map (
            O => \N__31667\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\
        );

    \I__5744\ : InMux
    port map (
            O => \N__31664\,
            I => \current_shift_inst.control_input_cry_5\
        );

    \I__5743\ : CascadeMux
    port map (
            O => \N__31661\,
            I => \N__31658\
        );

    \I__5742\ : InMux
    port map (
            O => \N__31658\,
            I => \N__31655\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__31655\,
            I => \N__31652\
        );

    \I__5740\ : Odrv4
    port map (
            O => \N__31652\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\
        );

    \I__5739\ : InMux
    port map (
            O => \N__31649\,
            I => \current_shift_inst.control_input_cry_6\
        );

    \I__5738\ : InMux
    port map (
            O => \N__31646\,
            I => \N__31642\
        );

    \I__5737\ : InMux
    port map (
            O => \N__31645\,
            I => \N__31639\
        );

    \I__5736\ : LocalMux
    port map (
            O => \N__31642\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\
        );

    \I__5735\ : LocalMux
    port map (
            O => \N__31639\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\
        );

    \I__5734\ : InMux
    port map (
            O => \N__31634\,
            I => \N__31630\
        );

    \I__5733\ : InMux
    port map (
            O => \N__31633\,
            I => \N__31627\
        );

    \I__5732\ : LocalMux
    port map (
            O => \N__31630\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\
        );

    \I__5731\ : LocalMux
    port map (
            O => \N__31627\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\
        );

    \I__5730\ : InMux
    port map (
            O => \N__31622\,
            I => \N__31619\
        );

    \I__5729\ : LocalMux
    port map (
            O => \N__31619\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30\
        );

    \I__5728\ : CascadeMux
    port map (
            O => \N__31616\,
            I => \N__31611\
        );

    \I__5727\ : CascadeMux
    port map (
            O => \N__31615\,
            I => \N__31608\
        );

    \I__5726\ : InMux
    port map (
            O => \N__31614\,
            I => \N__31605\
        );

    \I__5725\ : InMux
    port map (
            O => \N__31611\,
            I => \N__31599\
        );

    \I__5724\ : InMux
    port map (
            O => \N__31608\,
            I => \N__31599\
        );

    \I__5723\ : LocalMux
    port map (
            O => \N__31605\,
            I => \N__31596\
        );

    \I__5722\ : InMux
    port map (
            O => \N__31604\,
            I => \N__31592\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__31599\,
            I => \N__31587\
        );

    \I__5720\ : Span4Mux_h
    port map (
            O => \N__31596\,
            I => \N__31587\
        );

    \I__5719\ : InMux
    port map (
            O => \N__31595\,
            I => \N__31584\
        );

    \I__5718\ : LocalMux
    port map (
            O => \N__31592\,
            I => \N__31581\
        );

    \I__5717\ : Odrv4
    port map (
            O => \N__31587\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__31584\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__5715\ : Odrv4
    port map (
            O => \N__31581\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__5714\ : InMux
    port map (
            O => \N__31574\,
            I => \N__31570\
        );

    \I__5713\ : CascadeMux
    port map (
            O => \N__31573\,
            I => \N__31566\
        );

    \I__5712\ : LocalMux
    port map (
            O => \N__31570\,
            I => \N__31562\
        );

    \I__5711\ : InMux
    port map (
            O => \N__31569\,
            I => \N__31559\
        );

    \I__5710\ : InMux
    port map (
            O => \N__31566\,
            I => \N__31554\
        );

    \I__5709\ : InMux
    port map (
            O => \N__31565\,
            I => \N__31554\
        );

    \I__5708\ : Span4Mux_v
    port map (
            O => \N__31562\,
            I => \N__31551\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__31559\,
            I => \N__31548\
        );

    \I__5706\ : LocalMux
    port map (
            O => \N__31554\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__5705\ : Odrv4
    port map (
            O => \N__31551\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__5704\ : Odrv4
    port map (
            O => \N__31548\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__5703\ : IoInMux
    port map (
            O => \N__31541\,
            I => \N__31516\
        );

    \I__5702\ : InMux
    port map (
            O => \N__31540\,
            I => \N__31499\
        );

    \I__5701\ : InMux
    port map (
            O => \N__31539\,
            I => \N__31499\
        );

    \I__5700\ : InMux
    port map (
            O => \N__31538\,
            I => \N__31499\
        );

    \I__5699\ : InMux
    port map (
            O => \N__31537\,
            I => \N__31499\
        );

    \I__5698\ : InMux
    port map (
            O => \N__31536\,
            I => \N__31492\
        );

    \I__5697\ : InMux
    port map (
            O => \N__31535\,
            I => \N__31492\
        );

    \I__5696\ : InMux
    port map (
            O => \N__31534\,
            I => \N__31492\
        );

    \I__5695\ : InMux
    port map (
            O => \N__31533\,
            I => \N__31483\
        );

    \I__5694\ : InMux
    port map (
            O => \N__31532\,
            I => \N__31483\
        );

    \I__5693\ : InMux
    port map (
            O => \N__31531\,
            I => \N__31483\
        );

    \I__5692\ : InMux
    port map (
            O => \N__31530\,
            I => \N__31483\
        );

    \I__5691\ : InMux
    port map (
            O => \N__31529\,
            I => \N__31476\
        );

    \I__5690\ : InMux
    port map (
            O => \N__31528\,
            I => \N__31476\
        );

    \I__5689\ : InMux
    port map (
            O => \N__31527\,
            I => \N__31476\
        );

    \I__5688\ : InMux
    port map (
            O => \N__31526\,
            I => \N__31467\
        );

    \I__5687\ : InMux
    port map (
            O => \N__31525\,
            I => \N__31467\
        );

    \I__5686\ : InMux
    port map (
            O => \N__31524\,
            I => \N__31467\
        );

    \I__5685\ : InMux
    port map (
            O => \N__31523\,
            I => \N__31467\
        );

    \I__5684\ : InMux
    port map (
            O => \N__31522\,
            I => \N__31458\
        );

    \I__5683\ : InMux
    port map (
            O => \N__31521\,
            I => \N__31458\
        );

    \I__5682\ : InMux
    port map (
            O => \N__31520\,
            I => \N__31458\
        );

    \I__5681\ : InMux
    port map (
            O => \N__31519\,
            I => \N__31458\
        );

    \I__5680\ : LocalMux
    port map (
            O => \N__31516\,
            I => \N__31455\
        );

    \I__5679\ : InMux
    port map (
            O => \N__31515\,
            I => \N__31446\
        );

    \I__5678\ : InMux
    port map (
            O => \N__31514\,
            I => \N__31446\
        );

    \I__5677\ : InMux
    port map (
            O => \N__31513\,
            I => \N__31446\
        );

    \I__5676\ : InMux
    port map (
            O => \N__31512\,
            I => \N__31446\
        );

    \I__5675\ : InMux
    port map (
            O => \N__31511\,
            I => \N__31437\
        );

    \I__5674\ : InMux
    port map (
            O => \N__31510\,
            I => \N__31437\
        );

    \I__5673\ : InMux
    port map (
            O => \N__31509\,
            I => \N__31437\
        );

    \I__5672\ : InMux
    port map (
            O => \N__31508\,
            I => \N__31437\
        );

    \I__5671\ : LocalMux
    port map (
            O => \N__31499\,
            I => \N__31430\
        );

    \I__5670\ : LocalMux
    port map (
            O => \N__31492\,
            I => \N__31430\
        );

    \I__5669\ : LocalMux
    port map (
            O => \N__31483\,
            I => \N__31430\
        );

    \I__5668\ : LocalMux
    port map (
            O => \N__31476\,
            I => \N__31427\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__31467\,
            I => \N__31424\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__31458\,
            I => \N__31421\
        );

    \I__5665\ : Span4Mux_s3_v
    port map (
            O => \N__31455\,
            I => \N__31418\
        );

    \I__5664\ : LocalMux
    port map (
            O => \N__31446\,
            I => \N__31411\
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__31437\,
            I => \N__31411\
        );

    \I__5662\ : Span4Mux_v
    port map (
            O => \N__31430\,
            I => \N__31411\
        );

    \I__5661\ : Span4Mux_h
    port map (
            O => \N__31427\,
            I => \N__31406\
        );

    \I__5660\ : Span4Mux_h
    port map (
            O => \N__31424\,
            I => \N__31406\
        );

    \I__5659\ : Span4Mux_h
    port map (
            O => \N__31421\,
            I => \N__31403\
        );

    \I__5658\ : Span4Mux_v
    port map (
            O => \N__31418\,
            I => \N__31400\
        );

    \I__5657\ : Odrv4
    port map (
            O => \N__31411\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__5656\ : Odrv4
    port map (
            O => \N__31406\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__5655\ : Odrv4
    port map (
            O => \N__31403\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__5654\ : Odrv4
    port map (
            O => \N__31400\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__5653\ : InMux
    port map (
            O => \N__31391\,
            I => \N__31386\
        );

    \I__5652\ : InMux
    port map (
            O => \N__31390\,
            I => \N__31381\
        );

    \I__5651\ : InMux
    port map (
            O => \N__31389\,
            I => \N__31381\
        );

    \I__5650\ : LocalMux
    port map (
            O => \N__31386\,
            I => \N__31376\
        );

    \I__5649\ : LocalMux
    port map (
            O => \N__31381\,
            I => \N__31373\
        );

    \I__5648\ : InMux
    port map (
            O => \N__31380\,
            I => \N__31368\
        );

    \I__5647\ : InMux
    port map (
            O => \N__31379\,
            I => \N__31368\
        );

    \I__5646\ : Span4Mux_v
    port map (
            O => \N__31376\,
            I => \N__31365\
        );

    \I__5645\ : Span4Mux_v
    port map (
            O => \N__31373\,
            I => \N__31362\
        );

    \I__5644\ : LocalMux
    port map (
            O => \N__31368\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__5643\ : Odrv4
    port map (
            O => \N__31365\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__5642\ : Odrv4
    port map (
            O => \N__31362\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__5641\ : InMux
    port map (
            O => \N__31355\,
            I => \N__31352\
        );

    \I__5640\ : LocalMux
    port map (
            O => \N__31352\,
            I => \N__31347\
        );

    \I__5639\ : InMux
    port map (
            O => \N__31351\,
            I => \N__31344\
        );

    \I__5638\ : InMux
    port map (
            O => \N__31350\,
            I => \N__31341\
        );

    \I__5637\ : Odrv12
    port map (
            O => \N__31347\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__31344\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\
        );

    \I__5635\ : LocalMux
    port map (
            O => \N__31341\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\
        );

    \I__5634\ : CascadeMux
    port map (
            O => \N__31334\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0_cascade_\
        );

    \I__5633\ : InMux
    port map (
            O => \N__31331\,
            I => \N__31328\
        );

    \I__5632\ : LocalMux
    port map (
            O => \N__31328\,
            I => \N__31323\
        );

    \I__5631\ : InMux
    port map (
            O => \N__31327\,
            I => \N__31320\
        );

    \I__5630\ : InMux
    port map (
            O => \N__31326\,
            I => \N__31317\
        );

    \I__5629\ : Span4Mux_v
    port map (
            O => \N__31323\,
            I => \N__31312\
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__31320\,
            I => \N__31312\
        );

    \I__5627\ : LocalMux
    port map (
            O => \N__31317\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__5626\ : Odrv4
    port map (
            O => \N__31312\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__5625\ : CascadeMux
    port map (
            O => \N__31307\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0_cascade_\
        );

    \I__5624\ : InMux
    port map (
            O => \N__31304\,
            I => \N__31298\
        );

    \I__5623\ : InMux
    port map (
            O => \N__31303\,
            I => \N__31298\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__31298\,
            I => \phase_controller_inst2.stoper_hc.runningZ0\
        );

    \I__5621\ : InMux
    port map (
            O => \N__31295\,
            I => \N__31291\
        );

    \I__5620\ : InMux
    port map (
            O => \N__31294\,
            I => \N__31287\
        );

    \I__5619\ : LocalMux
    port map (
            O => \N__31291\,
            I => \N__31284\
        );

    \I__5618\ : InMux
    port map (
            O => \N__31290\,
            I => \N__31281\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__31287\,
            I => \N__31277\
        );

    \I__5616\ : Span4Mux_v
    port map (
            O => \N__31284\,
            I => \N__31272\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__31281\,
            I => \N__31272\
        );

    \I__5614\ : InMux
    port map (
            O => \N__31280\,
            I => \N__31269\
        );

    \I__5613\ : Span4Mux_v
    port map (
            O => \N__31277\,
            I => \N__31264\
        );

    \I__5612\ : Span4Mux_h
    port map (
            O => \N__31272\,
            I => \N__31264\
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__31269\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__5610\ : Odrv4
    port map (
            O => \N__31264\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__5609\ : CascadeMux
    port map (
            O => \N__31259\,
            I => \N__31256\
        );

    \I__5608\ : InMux
    port map (
            O => \N__31256\,
            I => \N__31252\
        );

    \I__5607\ : InMux
    port map (
            O => \N__31255\,
            I => \N__31249\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__31252\,
            I => \N__31244\
        );

    \I__5605\ : LocalMux
    port map (
            O => \N__31249\,
            I => \N__31244\
        );

    \I__5604\ : Span4Mux_v
    port map (
            O => \N__31244\,
            I => \N__31238\
        );

    \I__5603\ : InMux
    port map (
            O => \N__31243\,
            I => \N__31231\
        );

    \I__5602\ : InMux
    port map (
            O => \N__31242\,
            I => \N__31231\
        );

    \I__5601\ : InMux
    port map (
            O => \N__31241\,
            I => \N__31231\
        );

    \I__5600\ : Odrv4
    port map (
            O => \N__31238\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__31231\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__5598\ : CascadeMux
    port map (
            O => \N__31226\,
            I => \N__31223\
        );

    \I__5597\ : InMux
    port map (
            O => \N__31223\,
            I => \N__31220\
        );

    \I__5596\ : LocalMux
    port map (
            O => \N__31220\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt30\
        );

    \I__5595\ : InMux
    port map (
            O => \N__31217\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_30\
        );

    \I__5594\ : CascadeMux
    port map (
            O => \N__31214\,
            I => \N__31211\
        );

    \I__5593\ : InMux
    port map (
            O => \N__31211\,
            I => \N__31208\
        );

    \I__5592\ : LocalMux
    port map (
            O => \N__31208\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt26\
        );

    \I__5591\ : InMux
    port map (
            O => \N__31205\,
            I => \N__31202\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__31202\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26\
        );

    \I__5589\ : InMux
    port map (
            O => \N__31199\,
            I => \N__31196\
        );

    \I__5588\ : LocalMux
    port map (
            O => \N__31196\,
            I => \N__31193\
        );

    \I__5587\ : Span4Mux_h
    port map (
            O => \N__31193\,
            I => \N__31189\
        );

    \I__5586\ : InMux
    port map (
            O => \N__31192\,
            I => \N__31186\
        );

    \I__5585\ : Odrv4
    port map (
            O => \N__31189\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__31186\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27\
        );

    \I__5583\ : CascadeMux
    port map (
            O => \N__31181\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27_cascade_\
        );

    \I__5582\ : InMux
    port map (
            O => \N__31178\,
            I => \N__31175\
        );

    \I__5581\ : LocalMux
    port map (
            O => \N__31175\,
            I => \N__31170\
        );

    \I__5580\ : InMux
    port map (
            O => \N__31174\,
            I => \N__31165\
        );

    \I__5579\ : InMux
    port map (
            O => \N__31173\,
            I => \N__31165\
        );

    \I__5578\ : Span4Mux_v
    port map (
            O => \N__31170\,
            I => \N__31159\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__31165\,
            I => \N__31159\
        );

    \I__5576\ : InMux
    port map (
            O => \N__31164\,
            I => \N__31156\
        );

    \I__5575\ : Span4Mux_h
    port map (
            O => \N__31159\,
            I => \N__31153\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__31156\,
            I => \N__31150\
        );

    \I__5573\ : Odrv4
    port map (
            O => \N__31153\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__5572\ : Odrv4
    port map (
            O => \N__31150\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__5571\ : InMux
    port map (
            O => \N__31145\,
            I => \N__31139\
        );

    \I__5570\ : InMux
    port map (
            O => \N__31144\,
            I => \N__31139\
        );

    \I__5569\ : LocalMux
    port map (
            O => \N__31139\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\
        );

    \I__5568\ : InMux
    port map (
            O => \N__31136\,
            I => \N__31132\
        );

    \I__5567\ : InMux
    port map (
            O => \N__31135\,
            I => \N__31129\
        );

    \I__5566\ : LocalMux
    port map (
            O => \N__31132\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26\
        );

    \I__5565\ : LocalMux
    port map (
            O => \N__31129\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26\
        );

    \I__5564\ : CascadeMux
    port map (
            O => \N__31124\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26_cascade_\
        );

    \I__5563\ : InMux
    port map (
            O => \N__31121\,
            I => \N__31116\
        );

    \I__5562\ : InMux
    port map (
            O => \N__31120\,
            I => \N__31111\
        );

    \I__5561\ : InMux
    port map (
            O => \N__31119\,
            I => \N__31111\
        );

    \I__5560\ : LocalMux
    port map (
            O => \N__31116\,
            I => \N__31108\
        );

    \I__5559\ : LocalMux
    port map (
            O => \N__31111\,
            I => \N__31105\
        );

    \I__5558\ : Span4Mux_h
    port map (
            O => \N__31108\,
            I => \N__31101\
        );

    \I__5557\ : Span4Mux_h
    port map (
            O => \N__31105\,
            I => \N__31098\
        );

    \I__5556\ : InMux
    port map (
            O => \N__31104\,
            I => \N__31095\
        );

    \I__5555\ : Odrv4
    port map (
            O => \N__31101\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__5554\ : Odrv4
    port map (
            O => \N__31098\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__5553\ : LocalMux
    port map (
            O => \N__31095\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__5552\ : InMux
    port map (
            O => \N__31088\,
            I => \N__31082\
        );

    \I__5551\ : InMux
    port map (
            O => \N__31087\,
            I => \N__31082\
        );

    \I__5550\ : LocalMux
    port map (
            O => \N__31082\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\
        );

    \I__5549\ : CascadeMux
    port map (
            O => \N__31079\,
            I => \N__31076\
        );

    \I__5548\ : InMux
    port map (
            O => \N__31076\,
            I => \N__31073\
        );

    \I__5547\ : LocalMux
    port map (
            O => \N__31073\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\
        );

    \I__5546\ : InMux
    port map (
            O => \N__31070\,
            I => \N__31067\
        );

    \I__5545\ : LocalMux
    port map (
            O => \N__31067\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\
        );

    \I__5544\ : InMux
    port map (
            O => \N__31064\,
            I => \N__31061\
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__31061\,
            I => \N__31058\
        );

    \I__5542\ : Span4Mux_h
    port map (
            O => \N__31058\,
            I => \N__31055\
        );

    \I__5541\ : Odrv4
    port map (
            O => \N__31055\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt18\
        );

    \I__5540\ : CascadeMux
    port map (
            O => \N__31052\,
            I => \N__31049\
        );

    \I__5539\ : InMux
    port map (
            O => \N__31049\,
            I => \N__31046\
        );

    \I__5538\ : LocalMux
    port map (
            O => \N__31046\,
            I => \N__31043\
        );

    \I__5537\ : Span4Mux_v
    port map (
            O => \N__31043\,
            I => \N__31040\
        );

    \I__5536\ : Span4Mux_h
    port map (
            O => \N__31040\,
            I => \N__31037\
        );

    \I__5535\ : Odrv4
    port map (
            O => \N__31037\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\
        );

    \I__5534\ : InMux
    port map (
            O => \N__31034\,
            I => \N__31031\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__31031\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20\
        );

    \I__5532\ : CascadeMux
    port map (
            O => \N__31028\,
            I => \N__31025\
        );

    \I__5531\ : InMux
    port map (
            O => \N__31025\,
            I => \N__31022\
        );

    \I__5530\ : LocalMux
    port map (
            O => \N__31022\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt20\
        );

    \I__5529\ : InMux
    port map (
            O => \N__31019\,
            I => \N__31016\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__31016\,
            I => \N__31013\
        );

    \I__5527\ : Odrv4
    port map (
            O => \N__31013\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22\
        );

    \I__5526\ : CascadeMux
    port map (
            O => \N__31010\,
            I => \N__31007\
        );

    \I__5525\ : InMux
    port map (
            O => \N__31007\,
            I => \N__31004\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__31004\,
            I => \N__31001\
        );

    \I__5523\ : Odrv12
    port map (
            O => \N__31001\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt22\
        );

    \I__5522\ : InMux
    port map (
            O => \N__30998\,
            I => \N__30995\
        );

    \I__5521\ : LocalMux
    port map (
            O => \N__30995\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28\
        );

    \I__5520\ : CascadeMux
    port map (
            O => \N__30992\,
            I => \N__30989\
        );

    \I__5519\ : InMux
    port map (
            O => \N__30989\,
            I => \N__30986\
        );

    \I__5518\ : LocalMux
    port map (
            O => \N__30986\,
            I => \N__30983\
        );

    \I__5517\ : Odrv12
    port map (
            O => \N__30983\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt28\
        );

    \I__5516\ : CascadeMux
    port map (
            O => \N__30980\,
            I => \N__30977\
        );

    \I__5515\ : InMux
    port map (
            O => \N__30977\,
            I => \N__30974\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__30974\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\
        );

    \I__5513\ : CascadeMux
    port map (
            O => \N__30971\,
            I => \N__30968\
        );

    \I__5512\ : InMux
    port map (
            O => \N__30968\,
            I => \N__30965\
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__30965\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\
        );

    \I__5510\ : InMux
    port map (
            O => \N__30962\,
            I => \N__30959\
        );

    \I__5509\ : LocalMux
    port map (
            O => \N__30959\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\
        );

    \I__5508\ : CascadeMux
    port map (
            O => \N__30956\,
            I => \N__30953\
        );

    \I__5507\ : InMux
    port map (
            O => \N__30953\,
            I => \N__30950\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__30950\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\
        );

    \I__5505\ : InMux
    port map (
            O => \N__30947\,
            I => \N__30944\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__30944\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\
        );

    \I__5503\ : CascadeMux
    port map (
            O => \N__30941\,
            I => \N__30938\
        );

    \I__5502\ : InMux
    port map (
            O => \N__30938\,
            I => \N__30935\
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__30935\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\
        );

    \I__5500\ : InMux
    port map (
            O => \N__30932\,
            I => \N__30929\
        );

    \I__5499\ : LocalMux
    port map (
            O => \N__30929\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\
        );

    \I__5498\ : CascadeMux
    port map (
            O => \N__30926\,
            I => \N__30923\
        );

    \I__5497\ : InMux
    port map (
            O => \N__30923\,
            I => \N__30920\
        );

    \I__5496\ : LocalMux
    port map (
            O => \N__30920\,
            I => \N__30917\
        );

    \I__5495\ : Odrv4
    port map (
            O => \N__30917\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\
        );

    \I__5494\ : InMux
    port map (
            O => \N__30914\,
            I => \N__30911\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__30911\,
            I => \N__30908\
        );

    \I__5492\ : Odrv4
    port map (
            O => \N__30908\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\
        );

    \I__5491\ : CascadeMux
    port map (
            O => \N__30905\,
            I => \N__30902\
        );

    \I__5490\ : InMux
    port map (
            O => \N__30902\,
            I => \N__30899\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__30899\,
            I => \N__30896\
        );

    \I__5488\ : Odrv4
    port map (
            O => \N__30896\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\
        );

    \I__5487\ : InMux
    port map (
            O => \N__30893\,
            I => \N__30890\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__30890\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\
        );

    \I__5485\ : InMux
    port map (
            O => \N__30887\,
            I => \N__30884\
        );

    \I__5484\ : LocalMux
    port map (
            O => \N__30884\,
            I => \N__30881\
        );

    \I__5483\ : Odrv4
    port map (
            O => \N__30881\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\
        );

    \I__5482\ : CascadeMux
    port map (
            O => \N__30878\,
            I => \N__30875\
        );

    \I__5481\ : InMux
    port map (
            O => \N__30875\,
            I => \N__30872\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__30872\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\
        );

    \I__5479\ : CascadeMux
    port map (
            O => \N__30869\,
            I => \N__30865\
        );

    \I__5478\ : CascadeMux
    port map (
            O => \N__30868\,
            I => \N__30862\
        );

    \I__5477\ : InMux
    port map (
            O => \N__30865\,
            I => \N__30857\
        );

    \I__5476\ : InMux
    port map (
            O => \N__30862\,
            I => \N__30857\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__30857\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_22\
        );

    \I__5474\ : InMux
    port map (
            O => \N__30854\,
            I => \N__30848\
        );

    \I__5473\ : InMux
    port map (
            O => \N__30853\,
            I => \N__30848\
        );

    \I__5472\ : LocalMux
    port map (
            O => \N__30848\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_23\
        );

    \I__5471\ : InMux
    port map (
            O => \N__30845\,
            I => \N__30842\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__30842\,
            I => \N__30839\
        );

    \I__5469\ : Span4Mux_h
    port map (
            O => \N__30839\,
            I => \N__30835\
        );

    \I__5468\ : InMux
    port map (
            O => \N__30838\,
            I => \N__30832\
        );

    \I__5467\ : Span4Mux_v
    port map (
            O => \N__30835\,
            I => \N__30826\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__30832\,
            I => \N__30826\
        );

    \I__5465\ : InMux
    port map (
            O => \N__30831\,
            I => \N__30823\
        );

    \I__5464\ : Span4Mux_h
    port map (
            O => \N__30826\,
            I => \N__30820\
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__30823\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4\
        );

    \I__5462\ : Odrv4
    port map (
            O => \N__30820\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4\
        );

    \I__5461\ : InMux
    port map (
            O => \N__30815\,
            I => \N__30811\
        );

    \I__5460\ : InMux
    port map (
            O => \N__30814\,
            I => \N__30808\
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__30811\,
            I => \N__30804\
        );

    \I__5458\ : LocalMux
    port map (
            O => \N__30808\,
            I => \N__30801\
        );

    \I__5457\ : CascadeMux
    port map (
            O => \N__30807\,
            I => \N__30797\
        );

    \I__5456\ : Span4Mux_h
    port map (
            O => \N__30804\,
            I => \N__30792\
        );

    \I__5455\ : Span4Mux_v
    port map (
            O => \N__30801\,
            I => \N__30792\
        );

    \I__5454\ : InMux
    port map (
            O => \N__30800\,
            I => \N__30787\
        );

    \I__5453\ : InMux
    port map (
            O => \N__30797\,
            I => \N__30787\
        );

    \I__5452\ : Odrv4
    port map (
            O => \N__30792\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__5451\ : LocalMux
    port map (
            O => \N__30787\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__5450\ : CascadeMux
    port map (
            O => \N__30782\,
            I => \N__30779\
        );

    \I__5449\ : InMux
    port map (
            O => \N__30779\,
            I => \N__30776\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__30776\,
            I => \N__30773\
        );

    \I__5447\ : Odrv4
    port map (
            O => \N__30773\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\
        );

    \I__5446\ : InMux
    port map (
            O => \N__30770\,
            I => \N__30767\
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__30767\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\
        );

    \I__5444\ : InMux
    port map (
            O => \N__30764\,
            I => \N__30761\
        );

    \I__5443\ : LocalMux
    port map (
            O => \N__30761\,
            I => \N__30758\
        );

    \I__5442\ : Odrv12
    port map (
            O => \N__30758\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\
        );

    \I__5441\ : CascadeMux
    port map (
            O => \N__30755\,
            I => \N__30752\
        );

    \I__5440\ : InMux
    port map (
            O => \N__30752\,
            I => \N__30749\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__30749\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\
        );

    \I__5438\ : InMux
    port map (
            O => \N__30746\,
            I => \N__30743\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__30743\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\
        );

    \I__5436\ : CascadeMux
    port map (
            O => \N__30740\,
            I => \N__30737\
        );

    \I__5435\ : InMux
    port map (
            O => \N__30737\,
            I => \N__30734\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__30734\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\
        );

    \I__5433\ : CascadeMux
    port map (
            O => \N__30731\,
            I => \N__30728\
        );

    \I__5432\ : InMux
    port map (
            O => \N__30728\,
            I => \N__30725\
        );

    \I__5431\ : LocalMux
    port map (
            O => \N__30725\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\
        );

    \I__5430\ : InMux
    port map (
            O => \N__30722\,
            I => \N__30719\
        );

    \I__5429\ : LocalMux
    port map (
            O => \N__30719\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\
        );

    \I__5428\ : InMux
    port map (
            O => \N__30716\,
            I => \N__30713\
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__30713\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\
        );

    \I__5426\ : CascadeMux
    port map (
            O => \N__30710\,
            I => \N__30707\
        );

    \I__5425\ : InMux
    port map (
            O => \N__30707\,
            I => \N__30704\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__30704\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\
        );

    \I__5423\ : InMux
    port map (
            O => \N__30701\,
            I => \N__30698\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__30698\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\
        );

    \I__5421\ : CascadeMux
    port map (
            O => \N__30695\,
            I => \N__30692\
        );

    \I__5420\ : InMux
    port map (
            O => \N__30692\,
            I => \N__30689\
        );

    \I__5419\ : LocalMux
    port map (
            O => \N__30689\,
            I => \N__30686\
        );

    \I__5418\ : Odrv4
    port map (
            O => \N__30686\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\
        );

    \I__5417\ : CascadeMux
    port map (
            O => \N__30683\,
            I => \N__30680\
        );

    \I__5416\ : InMux
    port map (
            O => \N__30680\,
            I => \N__30677\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__30677\,
            I => \N__30674\
        );

    \I__5414\ : Span4Mux_h
    port map (
            O => \N__30674\,
            I => \N__30671\
        );

    \I__5413\ : Span4Mux_h
    port map (
            O => \N__30671\,
            I => \N__30668\
        );

    \I__5412\ : Span4Mux_h
    port map (
            O => \N__30668\,
            I => \N__30665\
        );

    \I__5411\ : Span4Mux_h
    port map (
            O => \N__30665\,
            I => \N__30662\
        );

    \I__5410\ : Odrv4
    port map (
            O => \N__30662\,
            I => \pwm_generator_inst.un2_threshold_2_11\
        );

    \I__5409\ : InMux
    port map (
            O => \N__30659\,
            I => \N__30656\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__30656\,
            I => \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0\
        );

    \I__5407\ : InMux
    port map (
            O => \N__30653\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_10\
        );

    \I__5406\ : CascadeMux
    port map (
            O => \N__30650\,
            I => \N__30647\
        );

    \I__5405\ : InMux
    port map (
            O => \N__30647\,
            I => \N__30644\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__30644\,
            I => \N__30641\
        );

    \I__5403\ : Span4Mux_v
    port map (
            O => \N__30641\,
            I => \N__30638\
        );

    \I__5402\ : Sp12to4
    port map (
            O => \N__30638\,
            I => \N__30635\
        );

    \I__5401\ : Span12Mux_h
    port map (
            O => \N__30635\,
            I => \N__30632\
        );

    \I__5400\ : Odrv12
    port map (
            O => \N__30632\,
            I => \pwm_generator_inst.un2_threshold_2_12\
        );

    \I__5399\ : InMux
    port map (
            O => \N__30629\,
            I => \N__30626\
        );

    \I__5398\ : LocalMux
    port map (
            O => \N__30626\,
            I => \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0\
        );

    \I__5397\ : InMux
    port map (
            O => \N__30623\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_11\
        );

    \I__5396\ : CascadeMux
    port map (
            O => \N__30620\,
            I => \N__30617\
        );

    \I__5395\ : InMux
    port map (
            O => \N__30617\,
            I => \N__30614\
        );

    \I__5394\ : LocalMux
    port map (
            O => \N__30614\,
            I => \N__30611\
        );

    \I__5393\ : Span4Mux_v
    port map (
            O => \N__30611\,
            I => \N__30608\
        );

    \I__5392\ : Sp12to4
    port map (
            O => \N__30608\,
            I => \N__30605\
        );

    \I__5391\ : Span12Mux_h
    port map (
            O => \N__30605\,
            I => \N__30602\
        );

    \I__5390\ : Odrv12
    port map (
            O => \N__30602\,
            I => \pwm_generator_inst.un2_threshold_2_13\
        );

    \I__5389\ : InMux
    port map (
            O => \N__30599\,
            I => \N__30596\
        );

    \I__5388\ : LocalMux
    port map (
            O => \N__30596\,
            I => \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0\
        );

    \I__5387\ : InMux
    port map (
            O => \N__30593\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_12\
        );

    \I__5386\ : CascadeMux
    port map (
            O => \N__30590\,
            I => \N__30587\
        );

    \I__5385\ : InMux
    port map (
            O => \N__30587\,
            I => \N__30584\
        );

    \I__5384\ : LocalMux
    port map (
            O => \N__30584\,
            I => \N__30581\
        );

    \I__5383\ : Span4Mux_v
    port map (
            O => \N__30581\,
            I => \N__30578\
        );

    \I__5382\ : Span4Mux_h
    port map (
            O => \N__30578\,
            I => \N__30575\
        );

    \I__5381\ : Sp12to4
    port map (
            O => \N__30575\,
            I => \N__30572\
        );

    \I__5380\ : Odrv12
    port map (
            O => \N__30572\,
            I => \pwm_generator_inst.un2_threshold_2_14\
        );

    \I__5379\ : InMux
    port map (
            O => \N__30569\,
            I => \N__30566\
        );

    \I__5378\ : LocalMux
    port map (
            O => \N__30566\,
            I => \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0\
        );

    \I__5377\ : InMux
    port map (
            O => \N__30563\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_13\
        );

    \I__5376\ : CascadeMux
    port map (
            O => \N__30560\,
            I => \N__30557\
        );

    \I__5375\ : InMux
    port map (
            O => \N__30557\,
            I => \N__30554\
        );

    \I__5374\ : LocalMux
    port map (
            O => \N__30554\,
            I => \N__30551\
        );

    \I__5373\ : Odrv12
    port map (
            O => \N__30551\,
            I => \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\
        );

    \I__5372\ : InMux
    port map (
            O => \N__30548\,
            I => \N__30545\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__30545\,
            I => \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0\
        );

    \I__5370\ : InMux
    port map (
            O => \N__30542\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_14\
        );

    \I__5369\ : InMux
    port map (
            O => \N__30539\,
            I => \N__30536\
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__30536\,
            I => \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\
        );

    \I__5367\ : InMux
    port map (
            O => \N__30533\,
            I => \bfn_10_28_0_\
        );

    \I__5366\ : CascadeMux
    port map (
            O => \N__30530\,
            I => \N__30526\
        );

    \I__5365\ : CascadeMux
    port map (
            O => \N__30529\,
            I => \N__30522\
        );

    \I__5364\ : InMux
    port map (
            O => \N__30526\,
            I => \N__30516\
        );

    \I__5363\ : InMux
    port map (
            O => \N__30525\,
            I => \N__30513\
        );

    \I__5362\ : InMux
    port map (
            O => \N__30522\,
            I => \N__30510\
        );

    \I__5361\ : CascadeMux
    port map (
            O => \N__30521\,
            I => \N__30507\
        );

    \I__5360\ : CascadeMux
    port map (
            O => \N__30520\,
            I => \N__30504\
        );

    \I__5359\ : InMux
    port map (
            O => \N__30519\,
            I => \N__30495\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__30516\,
            I => \N__30492\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__30513\,
            I => \N__30487\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__30510\,
            I => \N__30487\
        );

    \I__5355\ : InMux
    port map (
            O => \N__30507\,
            I => \N__30482\
        );

    \I__5354\ : InMux
    port map (
            O => \N__30504\,
            I => \N__30482\
        );

    \I__5353\ : InMux
    port map (
            O => \N__30503\,
            I => \N__30477\
        );

    \I__5352\ : InMux
    port map (
            O => \N__30502\,
            I => \N__30477\
        );

    \I__5351\ : InMux
    port map (
            O => \N__30501\,
            I => \N__30474\
        );

    \I__5350\ : InMux
    port map (
            O => \N__30500\,
            I => \N__30471\
        );

    \I__5349\ : InMux
    port map (
            O => \N__30499\,
            I => \N__30468\
        );

    \I__5348\ : InMux
    port map (
            O => \N__30498\,
            I => \N__30465\
        );

    \I__5347\ : LocalMux
    port map (
            O => \N__30495\,
            I => \N__30462\
        );

    \I__5346\ : Span4Mux_v
    port map (
            O => \N__30492\,
            I => \N__30457\
        );

    \I__5345\ : Span4Mux_v
    port map (
            O => \N__30487\,
            I => \N__30457\
        );

    \I__5344\ : LocalMux
    port map (
            O => \N__30482\,
            I => \N__30454\
        );

    \I__5343\ : LocalMux
    port map (
            O => \N__30477\,
            I => \N__30449\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__30474\,
            I => \N__30449\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__30471\,
            I => \N__30440\
        );

    \I__5340\ : LocalMux
    port map (
            O => \N__30468\,
            I => \N__30440\
        );

    \I__5339\ : LocalMux
    port map (
            O => \N__30465\,
            I => \N__30440\
        );

    \I__5338\ : Span4Mux_s2_h
    port map (
            O => \N__30462\,
            I => \N__30440\
        );

    \I__5337\ : Span4Mux_h
    port map (
            O => \N__30457\,
            I => \N__30437\
        );

    \I__5336\ : Span4Mux_h
    port map (
            O => \N__30454\,
            I => \N__30432\
        );

    \I__5335\ : Span4Mux_h
    port map (
            O => \N__30449\,
            I => \N__30432\
        );

    \I__5334\ : Span4Mux_h
    port map (
            O => \N__30440\,
            I => \N__30429\
        );

    \I__5333\ : Span4Mux_h
    port map (
            O => \N__30437\,
            I => \N__30426\
        );

    \I__5332\ : Span4Mux_h
    port map (
            O => \N__30432\,
            I => \N__30423\
        );

    \I__5331\ : Span4Mux_h
    port map (
            O => \N__30429\,
            I => \N__30420\
        );

    \I__5330\ : Odrv4
    port map (
            O => \N__30426\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__5329\ : Odrv4
    port map (
            O => \N__30423\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__5328\ : Odrv4
    port map (
            O => \N__30420\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__5327\ : InMux
    port map (
            O => \N__30413\,
            I => \N__30410\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__30410\,
            I => \N__30407\
        );

    \I__5325\ : Span4Mux_v
    port map (
            O => \N__30407\,
            I => \N__30404\
        );

    \I__5324\ : Sp12to4
    port map (
            O => \N__30404\,
            I => \N__30401\
        );

    \I__5323\ : Span12Mux_h
    port map (
            O => \N__30401\,
            I => \N__30398\
        );

    \I__5322\ : Odrv12
    port map (
            O => \N__30398\,
            I => \pwm_generator_inst.un2_threshold_2_4\
        );

    \I__5321\ : CascadeMux
    port map (
            O => \N__30395\,
            I => \N__30392\
        );

    \I__5320\ : InMux
    port map (
            O => \N__30392\,
            I => \N__30389\
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__30389\,
            I => \N__30386\
        );

    \I__5318\ : Span4Mux_h
    port map (
            O => \N__30386\,
            I => \N__30383\
        );

    \I__5317\ : Span4Mux_h
    port map (
            O => \N__30383\,
            I => \N__30380\
        );

    \I__5316\ : Span4Mux_h
    port map (
            O => \N__30380\,
            I => \N__30377\
        );

    \I__5315\ : Odrv4
    port map (
            O => \N__30377\,
            I => \pwm_generator_inst.un2_threshold_1_19\
        );

    \I__5314\ : InMux
    port map (
            O => \N__30374\,
            I => \N__30371\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__30371\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01\
        );

    \I__5312\ : InMux
    port map (
            O => \N__30368\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_3\
        );

    \I__5311\ : InMux
    port map (
            O => \N__30365\,
            I => \N__30362\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__30362\,
            I => \N__30359\
        );

    \I__5309\ : Span4Mux_v
    port map (
            O => \N__30359\,
            I => \N__30356\
        );

    \I__5308\ : Sp12to4
    port map (
            O => \N__30356\,
            I => \N__30353\
        );

    \I__5307\ : Span12Mux_h
    port map (
            O => \N__30353\,
            I => \N__30350\
        );

    \I__5306\ : Odrv12
    port map (
            O => \N__30350\,
            I => \pwm_generator_inst.un2_threshold_2_5\
        );

    \I__5305\ : CascadeMux
    port map (
            O => \N__30347\,
            I => \N__30344\
        );

    \I__5304\ : InMux
    port map (
            O => \N__30344\,
            I => \N__30341\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__30341\,
            I => \N__30338\
        );

    \I__5302\ : Span4Mux_v
    port map (
            O => \N__30338\,
            I => \N__30335\
        );

    \I__5301\ : Sp12to4
    port map (
            O => \N__30335\,
            I => \N__30332\
        );

    \I__5300\ : Odrv12
    port map (
            O => \N__30332\,
            I => \pwm_generator_inst.un2_threshold_1_20\
        );

    \I__5299\ : InMux
    port map (
            O => \N__30329\,
            I => \N__30326\
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__30326\,
            I => \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0\
        );

    \I__5297\ : InMux
    port map (
            O => \N__30323\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_4\
        );

    \I__5296\ : InMux
    port map (
            O => \N__30320\,
            I => \N__30317\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__30317\,
            I => \N__30314\
        );

    \I__5294\ : Span4Mux_v
    port map (
            O => \N__30314\,
            I => \N__30311\
        );

    \I__5293\ : Sp12to4
    port map (
            O => \N__30311\,
            I => \N__30308\
        );

    \I__5292\ : Span12Mux_h
    port map (
            O => \N__30308\,
            I => \N__30305\
        );

    \I__5291\ : Odrv12
    port map (
            O => \N__30305\,
            I => \pwm_generator_inst.un2_threshold_2_6\
        );

    \I__5290\ : CascadeMux
    port map (
            O => \N__30302\,
            I => \N__30299\
        );

    \I__5289\ : InMux
    port map (
            O => \N__30299\,
            I => \N__30296\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__30296\,
            I => \N__30293\
        );

    \I__5287\ : Sp12to4
    port map (
            O => \N__30293\,
            I => \N__30290\
        );

    \I__5286\ : Span12Mux_s5_v
    port map (
            O => \N__30290\,
            I => \N__30287\
        );

    \I__5285\ : Odrv12
    port map (
            O => \N__30287\,
            I => \pwm_generator_inst.un2_threshold_1_21\
        );

    \I__5284\ : InMux
    port map (
            O => \N__30284\,
            I => \N__30281\
        );

    \I__5283\ : LocalMux
    port map (
            O => \N__30281\,
            I => \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0\
        );

    \I__5282\ : InMux
    port map (
            O => \N__30278\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_5\
        );

    \I__5281\ : InMux
    port map (
            O => \N__30275\,
            I => \N__30272\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__30272\,
            I => \N__30269\
        );

    \I__5279\ : Span12Mux_s7_v
    port map (
            O => \N__30269\,
            I => \N__30266\
        );

    \I__5278\ : Span12Mux_h
    port map (
            O => \N__30266\,
            I => \N__30263\
        );

    \I__5277\ : Odrv12
    port map (
            O => \N__30263\,
            I => \pwm_generator_inst.un2_threshold_2_7\
        );

    \I__5276\ : CascadeMux
    port map (
            O => \N__30260\,
            I => \N__30257\
        );

    \I__5275\ : InMux
    port map (
            O => \N__30257\,
            I => \N__30254\
        );

    \I__5274\ : LocalMux
    port map (
            O => \N__30254\,
            I => \N__30251\
        );

    \I__5273\ : Sp12to4
    port map (
            O => \N__30251\,
            I => \N__30248\
        );

    \I__5272\ : Span12Mux_s5_v
    port map (
            O => \N__30248\,
            I => \N__30245\
        );

    \I__5271\ : Odrv12
    port map (
            O => \N__30245\,
            I => \pwm_generator_inst.un2_threshold_1_22\
        );

    \I__5270\ : InMux
    port map (
            O => \N__30242\,
            I => \N__30239\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__30239\,
            I => \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0\
        );

    \I__5268\ : InMux
    port map (
            O => \N__30236\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_6\
        );

    \I__5267\ : InMux
    port map (
            O => \N__30233\,
            I => \N__30230\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__30230\,
            I => \N__30227\
        );

    \I__5265\ : Span4Mux_v
    port map (
            O => \N__30227\,
            I => \N__30224\
        );

    \I__5264\ : Sp12to4
    port map (
            O => \N__30224\,
            I => \N__30221\
        );

    \I__5263\ : Odrv12
    port map (
            O => \N__30221\,
            I => \pwm_generator_inst.un2_threshold_1_23\
        );

    \I__5262\ : CascadeMux
    port map (
            O => \N__30218\,
            I => \N__30215\
        );

    \I__5261\ : InMux
    port map (
            O => \N__30215\,
            I => \N__30212\
        );

    \I__5260\ : LocalMux
    port map (
            O => \N__30212\,
            I => \N__30209\
        );

    \I__5259\ : Span4Mux_v
    port map (
            O => \N__30209\,
            I => \N__30206\
        );

    \I__5258\ : Sp12to4
    port map (
            O => \N__30206\,
            I => \N__30203\
        );

    \I__5257\ : Span12Mux_h
    port map (
            O => \N__30203\,
            I => \N__30200\
        );

    \I__5256\ : Odrv12
    port map (
            O => \N__30200\,
            I => \pwm_generator_inst.un2_threshold_2_8\
        );

    \I__5255\ : InMux
    port map (
            O => \N__30197\,
            I => \N__30194\
        );

    \I__5254\ : LocalMux
    port map (
            O => \N__30194\,
            I => \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0\
        );

    \I__5253\ : InMux
    port map (
            O => \N__30191\,
            I => \bfn_10_27_0_\
        );

    \I__5252\ : InMux
    port map (
            O => \N__30188\,
            I => \N__30185\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__30185\,
            I => \N__30182\
        );

    \I__5250\ : Span4Mux_h
    port map (
            O => \N__30182\,
            I => \N__30179\
        );

    \I__5249\ : Span4Mux_h
    port map (
            O => \N__30179\,
            I => \N__30176\
        );

    \I__5248\ : Span4Mux_h
    port map (
            O => \N__30176\,
            I => \N__30173\
        );

    \I__5247\ : Odrv4
    port map (
            O => \N__30173\,
            I => \pwm_generator_inst.un2_threshold_1_24\
        );

    \I__5246\ : CascadeMux
    port map (
            O => \N__30170\,
            I => \N__30167\
        );

    \I__5245\ : InMux
    port map (
            O => \N__30167\,
            I => \N__30164\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__30164\,
            I => \N__30161\
        );

    \I__5243\ : Span4Mux_v
    port map (
            O => \N__30161\,
            I => \N__30158\
        );

    \I__5242\ : Span4Mux_h
    port map (
            O => \N__30158\,
            I => \N__30155\
        );

    \I__5241\ : Span4Mux_h
    port map (
            O => \N__30155\,
            I => \N__30152\
        );

    \I__5240\ : Span4Mux_h
    port map (
            O => \N__30152\,
            I => \N__30149\
        );

    \I__5239\ : Odrv4
    port map (
            O => \N__30149\,
            I => \pwm_generator_inst.un2_threshold_2_9\
        );

    \I__5238\ : InMux
    port map (
            O => \N__30146\,
            I => \N__30143\
        );

    \I__5237\ : LocalMux
    port map (
            O => \N__30143\,
            I => \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0\
        );

    \I__5236\ : InMux
    port map (
            O => \N__30140\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_8\
        );

    \I__5235\ : CascadeMux
    port map (
            O => \N__30137\,
            I => \N__30134\
        );

    \I__5234\ : InMux
    port map (
            O => \N__30134\,
            I => \N__30131\
        );

    \I__5233\ : LocalMux
    port map (
            O => \N__30131\,
            I => \N__30128\
        );

    \I__5232\ : Span4Mux_v
    port map (
            O => \N__30128\,
            I => \N__30125\
        );

    \I__5231\ : Sp12to4
    port map (
            O => \N__30125\,
            I => \N__30122\
        );

    \I__5230\ : Span12Mux_h
    port map (
            O => \N__30122\,
            I => \N__30119\
        );

    \I__5229\ : Odrv12
    port map (
            O => \N__30119\,
            I => \pwm_generator_inst.un2_threshold_2_10\
        );

    \I__5228\ : InMux
    port map (
            O => \N__30116\,
            I => \N__30113\
        );

    \I__5227\ : LocalMux
    port map (
            O => \N__30113\,
            I => \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0\
        );

    \I__5226\ : InMux
    port map (
            O => \N__30110\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_9\
        );

    \I__5225\ : InMux
    port map (
            O => \N__30107\,
            I => \N__30104\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__30104\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30\
        );

    \I__5223\ : InMux
    port map (
            O => \N__30101\,
            I => \N__30098\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__30098\,
            I => \N__30095\
        );

    \I__5221\ : Span4Mux_v
    port map (
            O => \N__30095\,
            I => \N__30092\
        );

    \I__5220\ : Sp12to4
    port map (
            O => \N__30092\,
            I => \N__30089\
        );

    \I__5219\ : Span12Mux_h
    port map (
            O => \N__30089\,
            I => \N__30086\
        );

    \I__5218\ : Odrv12
    port map (
            O => \N__30086\,
            I => \pwm_generator_inst.un2_threshold_2_0\
        );

    \I__5217\ : CascadeMux
    port map (
            O => \N__30083\,
            I => \N__30080\
        );

    \I__5216\ : InMux
    port map (
            O => \N__30080\,
            I => \N__30077\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__30077\,
            I => \N__30074\
        );

    \I__5214\ : Span4Mux_h
    port map (
            O => \N__30074\,
            I => \N__30071\
        );

    \I__5213\ : Span4Mux_h
    port map (
            O => \N__30071\,
            I => \N__30068\
        );

    \I__5212\ : Span4Mux_h
    port map (
            O => \N__30068\,
            I => \N__30065\
        );

    \I__5211\ : Odrv4
    port map (
            O => \N__30065\,
            I => \pwm_generator_inst.un2_threshold_1_15\
        );

    \I__5210\ : InMux
    port map (
            O => \N__30062\,
            I => \N__30059\
        );

    \I__5209\ : LocalMux
    port map (
            O => \N__30059\,
            I => \pwm_generator_inst.un3_threshold_axbZ0Z_4\
        );

    \I__5208\ : InMux
    port map (
            O => \N__30056\,
            I => \N__30053\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__30053\,
            I => \N__30050\
        );

    \I__5206\ : Span4Mux_v
    port map (
            O => \N__30050\,
            I => \N__30047\
        );

    \I__5205\ : Sp12to4
    port map (
            O => \N__30047\,
            I => \N__30044\
        );

    \I__5204\ : Span12Mux_h
    port map (
            O => \N__30044\,
            I => \N__30041\
        );

    \I__5203\ : Odrv12
    port map (
            O => \N__30041\,
            I => \pwm_generator_inst.un2_threshold_2_1\
        );

    \I__5202\ : CascadeMux
    port map (
            O => \N__30038\,
            I => \N__30035\
        );

    \I__5201\ : InMux
    port map (
            O => \N__30035\,
            I => \N__30032\
        );

    \I__5200\ : LocalMux
    port map (
            O => \N__30032\,
            I => \N__30029\
        );

    \I__5199\ : Span4Mux_h
    port map (
            O => \N__30029\,
            I => \N__30026\
        );

    \I__5198\ : Span4Mux_h
    port map (
            O => \N__30026\,
            I => \N__30023\
        );

    \I__5197\ : Span4Mux_h
    port map (
            O => \N__30023\,
            I => \N__30020\
        );

    \I__5196\ : Odrv4
    port map (
            O => \N__30020\,
            I => \pwm_generator_inst.un2_threshold_1_16\
        );

    \I__5195\ : CascadeMux
    port map (
            O => \N__30017\,
            I => \N__30014\
        );

    \I__5194\ : InMux
    port map (
            O => \N__30014\,
            I => \N__30011\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__30011\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701\
        );

    \I__5192\ : InMux
    port map (
            O => \N__30008\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_0\
        );

    \I__5191\ : InMux
    port map (
            O => \N__30005\,
            I => \N__30002\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__30002\,
            I => \N__29999\
        );

    \I__5189\ : Span4Mux_v
    port map (
            O => \N__29999\,
            I => \N__29996\
        );

    \I__5188\ : Sp12to4
    port map (
            O => \N__29996\,
            I => \N__29993\
        );

    \I__5187\ : Span12Mux_h
    port map (
            O => \N__29993\,
            I => \N__29990\
        );

    \I__5186\ : Odrv12
    port map (
            O => \N__29990\,
            I => \pwm_generator_inst.un2_threshold_2_2\
        );

    \I__5185\ : CascadeMux
    port map (
            O => \N__29987\,
            I => \N__29984\
        );

    \I__5184\ : InMux
    port map (
            O => \N__29984\,
            I => \N__29981\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__29981\,
            I => \N__29978\
        );

    \I__5182\ : Span4Mux_h
    port map (
            O => \N__29978\,
            I => \N__29975\
        );

    \I__5181\ : Span4Mux_h
    port map (
            O => \N__29975\,
            I => \N__29972\
        );

    \I__5180\ : Span4Mux_h
    port map (
            O => \N__29972\,
            I => \N__29969\
        );

    \I__5179\ : Odrv4
    port map (
            O => \N__29969\,
            I => \pwm_generator_inst.un2_threshold_1_17\
        );

    \I__5178\ : InMux
    port map (
            O => \N__29966\,
            I => \N__29963\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__29963\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801\
        );

    \I__5176\ : InMux
    port map (
            O => \N__29960\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_1\
        );

    \I__5175\ : InMux
    port map (
            O => \N__29957\,
            I => \N__29954\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__29954\,
            I => \N__29951\
        );

    \I__5173\ : Span12Mux_h
    port map (
            O => \N__29951\,
            I => \N__29948\
        );

    \I__5172\ : Span12Mux_h
    port map (
            O => \N__29948\,
            I => \N__29945\
        );

    \I__5171\ : Odrv12
    port map (
            O => \N__29945\,
            I => \pwm_generator_inst.un2_threshold_2_3\
        );

    \I__5170\ : CascadeMux
    port map (
            O => \N__29942\,
            I => \N__29939\
        );

    \I__5169\ : InMux
    port map (
            O => \N__29939\,
            I => \N__29936\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__29936\,
            I => \N__29933\
        );

    \I__5167\ : Span4Mux_h
    port map (
            O => \N__29933\,
            I => \N__29930\
        );

    \I__5166\ : Span4Mux_h
    port map (
            O => \N__29930\,
            I => \N__29927\
        );

    \I__5165\ : Span4Mux_h
    port map (
            O => \N__29927\,
            I => \N__29924\
        );

    \I__5164\ : Odrv4
    port map (
            O => \N__29924\,
            I => \pwm_generator_inst.un2_threshold_1_18\
        );

    \I__5163\ : CascadeMux
    port map (
            O => \N__29921\,
            I => \N__29918\
        );

    \I__5162\ : InMux
    port map (
            O => \N__29918\,
            I => \N__29915\
        );

    \I__5161\ : LocalMux
    port map (
            O => \N__29915\,
            I => \N__29912\
        );

    \I__5160\ : Odrv4
    port map (
            O => \N__29912\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901\
        );

    \I__5159\ : InMux
    port map (
            O => \N__29909\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_2\
        );

    \I__5158\ : CascadeMux
    port map (
            O => \N__29906\,
            I => \N__29903\
        );

    \I__5157\ : InMux
    port map (
            O => \N__29903\,
            I => \N__29900\
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__29900\,
            I => \N__29897\
        );

    \I__5155\ : Odrv4
    port map (
            O => \N__29897\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt16\
        );

    \I__5154\ : InMux
    port map (
            O => \N__29894\,
            I => \N__29888\
        );

    \I__5153\ : InMux
    port map (
            O => \N__29893\,
            I => \N__29888\
        );

    \I__5152\ : LocalMux
    port map (
            O => \N__29888\,
            I => \N__29884\
        );

    \I__5151\ : InMux
    port map (
            O => \N__29887\,
            I => \N__29881\
        );

    \I__5150\ : Span4Mux_h
    port map (
            O => \N__29884\,
            I => \N__29878\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__29881\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__5148\ : Odrv4
    port map (
            O => \N__29878\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__5147\ : CascadeMux
    port map (
            O => \N__29873\,
            I => \N__29870\
        );

    \I__5146\ : InMux
    port map (
            O => \N__29870\,
            I => \N__29864\
        );

    \I__5145\ : InMux
    port map (
            O => \N__29869\,
            I => \N__29864\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__29864\,
            I => \N__29860\
        );

    \I__5143\ : InMux
    port map (
            O => \N__29863\,
            I => \N__29857\
        );

    \I__5142\ : Span4Mux_h
    port map (
            O => \N__29860\,
            I => \N__29854\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__29857\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__5140\ : Odrv4
    port map (
            O => \N__29854\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__5139\ : InMux
    port map (
            O => \N__29849\,
            I => \N__29846\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__29846\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\
        );

    \I__5137\ : InMux
    port map (
            O => \N__29843\,
            I => \N__29837\
        );

    \I__5136\ : InMux
    port map (
            O => \N__29842\,
            I => \N__29837\
        );

    \I__5135\ : LocalMux
    port map (
            O => \N__29837\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\
        );

    \I__5134\ : CascadeMux
    port map (
            O => \N__29834\,
            I => \N__29831\
        );

    \I__5133\ : InMux
    port map (
            O => \N__29831\,
            I => \N__29825\
        );

    \I__5132\ : InMux
    port map (
            O => \N__29830\,
            I => \N__29825\
        );

    \I__5131\ : LocalMux
    port map (
            O => \N__29825\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\
        );

    \I__5130\ : InMux
    port map (
            O => \N__29822\,
            I => \N__29819\
        );

    \I__5129\ : LocalMux
    port map (
            O => \N__29819\,
            I => \N__29814\
        );

    \I__5128\ : InMux
    port map (
            O => \N__29818\,
            I => \N__29809\
        );

    \I__5127\ : InMux
    port map (
            O => \N__29817\,
            I => \N__29809\
        );

    \I__5126\ : Span4Mux_v
    port map (
            O => \N__29814\,
            I => \N__29804\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__29809\,
            I => \N__29804\
        );

    \I__5124\ : Span4Mux_v
    port map (
            O => \N__29804\,
            I => \N__29800\
        );

    \I__5123\ : InMux
    port map (
            O => \N__29803\,
            I => \N__29797\
        );

    \I__5122\ : Odrv4
    port map (
            O => \N__29800\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\
        );

    \I__5121\ : LocalMux
    port map (
            O => \N__29797\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\
        );

    \I__5120\ : InMux
    port map (
            O => \N__29792\,
            I => \N__29789\
        );

    \I__5119\ : LocalMux
    port map (
            O => \N__29789\,
            I => \N__29785\
        );

    \I__5118\ : InMux
    port map (
            O => \N__29788\,
            I => \N__29782\
        );

    \I__5117\ : Odrv12
    port map (
            O => \N__29785\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__29782\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15\
        );

    \I__5115\ : CascadeMux
    port map (
            O => \N__29777\,
            I => \N__29774\
        );

    \I__5114\ : InMux
    port map (
            O => \N__29774\,
            I => \N__29771\
        );

    \I__5113\ : LocalMux
    port map (
            O => \N__29771\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\
        );

    \I__5112\ : CEMux
    port map (
            O => \N__29768\,
            I => \N__29735\
        );

    \I__5111\ : CEMux
    port map (
            O => \N__29767\,
            I => \N__29735\
        );

    \I__5110\ : CEMux
    port map (
            O => \N__29766\,
            I => \N__29735\
        );

    \I__5109\ : CEMux
    port map (
            O => \N__29765\,
            I => \N__29735\
        );

    \I__5108\ : CEMux
    port map (
            O => \N__29764\,
            I => \N__29735\
        );

    \I__5107\ : CEMux
    port map (
            O => \N__29763\,
            I => \N__29735\
        );

    \I__5106\ : CEMux
    port map (
            O => \N__29762\,
            I => \N__29735\
        );

    \I__5105\ : CEMux
    port map (
            O => \N__29761\,
            I => \N__29735\
        );

    \I__5104\ : CEMux
    port map (
            O => \N__29760\,
            I => \N__29735\
        );

    \I__5103\ : CEMux
    port map (
            O => \N__29759\,
            I => \N__29735\
        );

    \I__5102\ : CEMux
    port map (
            O => \N__29758\,
            I => \N__29735\
        );

    \I__5101\ : GlobalMux
    port map (
            O => \N__29735\,
            I => \N__29732\
        );

    \I__5100\ : gio2CtrlBuf
    port map (
            O => \N__29732\,
            I => \phase_controller_inst2.stoper_tr.un1_start_g\
        );

    \I__5099\ : CascadeMux
    port map (
            O => \N__29729\,
            I => \current_shift_inst.control_input_axb_0_cascade_\
        );

    \I__5098\ : InMux
    port map (
            O => \N__29726\,
            I => \N__29722\
        );

    \I__5097\ : InMux
    port map (
            O => \N__29725\,
            I => \N__29719\
        );

    \I__5096\ : LocalMux
    port map (
            O => \N__29722\,
            I => \N__29716\
        );

    \I__5095\ : LocalMux
    port map (
            O => \N__29719\,
            I => \N__29713\
        );

    \I__5094\ : Span4Mux_s2_h
    port map (
            O => \N__29716\,
            I => \N__29710\
        );

    \I__5093\ : Span4Mux_v
    port map (
            O => \N__29713\,
            I => \N__29707\
        );

    \I__5092\ : Span4Mux_h
    port map (
            O => \N__29710\,
            I => \N__29704\
        );

    \I__5091\ : Span4Mux_h
    port map (
            O => \N__29707\,
            I => \N__29701\
        );

    \I__5090\ : Span4Mux_h
    port map (
            O => \N__29704\,
            I => \N__29698\
        );

    \I__5089\ : Odrv4
    port map (
            O => \N__29701\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__5088\ : Odrv4
    port map (
            O => \N__29698\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__5087\ : InMux
    port map (
            O => \N__29693\,
            I => \N__29690\
        );

    \I__5086\ : LocalMux
    port map (
            O => \N__29690\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\
        );

    \I__5085\ : InMux
    port map (
            O => \N__29687\,
            I => \N__29684\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__29684\,
            I => \N__29681\
        );

    \I__5083\ : Span4Mux_h
    port map (
            O => \N__29681\,
            I => \N__29675\
        );

    \I__5082\ : InMux
    port map (
            O => \N__29680\,
            I => \N__29668\
        );

    \I__5081\ : InMux
    port map (
            O => \N__29679\,
            I => \N__29668\
        );

    \I__5080\ : InMux
    port map (
            O => \N__29678\,
            I => \N__29668\
        );

    \I__5079\ : Odrv4
    port map (
            O => \N__29675\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__29668\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__5077\ : InMux
    port map (
            O => \N__29663\,
            I => \N__29660\
        );

    \I__5076\ : LocalMux
    port map (
            O => \N__29660\,
            I => \N__29657\
        );

    \I__5075\ : Span4Mux_v
    port map (
            O => \N__29657\,
            I => \N__29653\
        );

    \I__5074\ : InMux
    port map (
            O => \N__29656\,
            I => \N__29650\
        );

    \I__5073\ : Odrv4
    port map (
            O => \N__29653\,
            I => \elapsed_time_ns_1_RNIV9PBB_0_21\
        );

    \I__5072\ : LocalMux
    port map (
            O => \N__29650\,
            I => \elapsed_time_ns_1_RNIV9PBB_0_21\
        );

    \I__5071\ : InMux
    port map (
            O => \N__29645\,
            I => \N__29642\
        );

    \I__5070\ : LocalMux
    port map (
            O => \N__29642\,
            I => \N__29637\
        );

    \I__5069\ : InMux
    port map (
            O => \N__29641\,
            I => \N__29632\
        );

    \I__5068\ : InMux
    port map (
            O => \N__29640\,
            I => \N__29632\
        );

    \I__5067\ : Span4Mux_v
    port map (
            O => \N__29637\,
            I => \N__29628\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__29632\,
            I => \N__29625\
        );

    \I__5065\ : InMux
    port map (
            O => \N__29631\,
            I => \N__29622\
        );

    \I__5064\ : Odrv4
    port map (
            O => \N__29628\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__5063\ : Odrv12
    port map (
            O => \N__29625\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__29622\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__5061\ : InMux
    port map (
            O => \N__29615\,
            I => \N__29612\
        );

    \I__5060\ : LocalMux
    port map (
            O => \N__29612\,
            I => \N__29608\
        );

    \I__5059\ : InMux
    port map (
            O => \N__29611\,
            I => \N__29605\
        );

    \I__5058\ : Odrv12
    port map (
            O => \N__29608\,
            I => \elapsed_time_ns_1_RNIU8PBB_0_20\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__29605\,
            I => \elapsed_time_ns_1_RNIU8PBB_0_20\
        );

    \I__5056\ : InMux
    port map (
            O => \N__29600\,
            I => \N__29597\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__29597\,
            I => \N__29594\
        );

    \I__5054\ : Span4Mux_h
    port map (
            O => \N__29594\,
            I => \N__29589\
        );

    \I__5053\ : InMux
    port map (
            O => \N__29593\,
            I => \N__29584\
        );

    \I__5052\ : InMux
    port map (
            O => \N__29592\,
            I => \N__29584\
        );

    \I__5051\ : Span4Mux_v
    port map (
            O => \N__29589\,
            I => \N__29579\
        );

    \I__5050\ : LocalMux
    port map (
            O => \N__29584\,
            I => \N__29579\
        );

    \I__5049\ : Span4Mux_h
    port map (
            O => \N__29579\,
            I => \N__29575\
        );

    \I__5048\ : InMux
    port map (
            O => \N__29578\,
            I => \N__29572\
        );

    \I__5047\ : Odrv4
    port map (
            O => \N__29575\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\
        );

    \I__5046\ : LocalMux
    port map (
            O => \N__29572\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\
        );

    \I__5045\ : InMux
    port map (
            O => \N__29567\,
            I => \N__29564\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__29564\,
            I => \N__29560\
        );

    \I__5043\ : InMux
    port map (
            O => \N__29563\,
            I => \N__29557\
        );

    \I__5042\ : Odrv12
    port map (
            O => \N__29560\,
            I => \elapsed_time_ns_1_RNILK91B_0_9\
        );

    \I__5041\ : LocalMux
    port map (
            O => \N__29557\,
            I => \elapsed_time_ns_1_RNILK91B_0_9\
        );

    \I__5040\ : CascadeMux
    port map (
            O => \N__29552\,
            I => \N__29549\
        );

    \I__5039\ : InMux
    port map (
            O => \N__29549\,
            I => \N__29546\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__29546\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\
        );

    \I__5037\ : InMux
    port map (
            O => \N__29543\,
            I => \N__29540\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__29540\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\
        );

    \I__5035\ : CascadeMux
    port map (
            O => \N__29537\,
            I => \N__29534\
        );

    \I__5034\ : InMux
    port map (
            O => \N__29534\,
            I => \N__29531\
        );

    \I__5033\ : LocalMux
    port map (
            O => \N__29531\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt20\
        );

    \I__5032\ : InMux
    port map (
            O => \N__29528\,
            I => \N__29522\
        );

    \I__5031\ : InMux
    port map (
            O => \N__29527\,
            I => \N__29522\
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__29522\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_20\
        );

    \I__5029\ : InMux
    port map (
            O => \N__29519\,
            I => \N__29512\
        );

    \I__5028\ : InMux
    port map (
            O => \N__29518\,
            I => \N__29512\
        );

    \I__5027\ : InMux
    port map (
            O => \N__29517\,
            I => \N__29509\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__29512\,
            I => \N__29506\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__29509\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__5024\ : Odrv4
    port map (
            O => \N__29506\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__5023\ : CascadeMux
    port map (
            O => \N__29501\,
            I => \N__29497\
        );

    \I__5022\ : InMux
    port map (
            O => \N__29500\,
            I => \N__29491\
        );

    \I__5021\ : InMux
    port map (
            O => \N__29497\,
            I => \N__29491\
        );

    \I__5020\ : InMux
    port map (
            O => \N__29496\,
            I => \N__29488\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__29491\,
            I => \N__29485\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__29488\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__5017\ : Odrv4
    port map (
            O => \N__29485\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__5016\ : CascadeMux
    port map (
            O => \N__29480\,
            I => \N__29476\
        );

    \I__5015\ : InMux
    port map (
            O => \N__29479\,
            I => \N__29471\
        );

    \I__5014\ : InMux
    port map (
            O => \N__29476\,
            I => \N__29471\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__29471\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_21\
        );

    \I__5012\ : InMux
    port map (
            O => \N__29468\,
            I => \N__29465\
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__29465\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20\
        );

    \I__5010\ : InMux
    port map (
            O => \N__29462\,
            I => \N__29459\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__29459\,
            I => \N__29455\
        );

    \I__5008\ : InMux
    port map (
            O => \N__29458\,
            I => \N__29451\
        );

    \I__5007\ : Span4Mux_v
    port map (
            O => \N__29455\,
            I => \N__29448\
        );

    \I__5006\ : InMux
    port map (
            O => \N__29454\,
            I => \N__29445\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__29451\,
            I => \N__29442\
        );

    \I__5004\ : Span4Mux_v
    port map (
            O => \N__29448\,
            I => \N__29436\
        );

    \I__5003\ : LocalMux
    port map (
            O => \N__29445\,
            I => \N__29436\
        );

    \I__5002\ : Span4Mux_h
    port map (
            O => \N__29442\,
            I => \N__29433\
        );

    \I__5001\ : InMux
    port map (
            O => \N__29441\,
            I => \N__29430\
        );

    \I__5000\ : Odrv4
    port map (
            O => \N__29436\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\
        );

    \I__4999\ : Odrv4
    port map (
            O => \N__29433\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__29430\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\
        );

    \I__4997\ : InMux
    port map (
            O => \N__29423\,
            I => \N__29420\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__29420\,
            I => \N__29416\
        );

    \I__4995\ : InMux
    port map (
            O => \N__29419\,
            I => \N__29412\
        );

    \I__4994\ : Span4Mux_v
    port map (
            O => \N__29416\,
            I => \N__29409\
        );

    \I__4993\ : InMux
    port map (
            O => \N__29415\,
            I => \N__29406\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__29412\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6\
        );

    \I__4991\ : Odrv4
    port map (
            O => \N__29409\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__29406\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6\
        );

    \I__4989\ : InMux
    port map (
            O => \N__29399\,
            I => \N__29396\
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__29396\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\
        );

    \I__4987\ : CascadeMux
    port map (
            O => \N__29393\,
            I => \N__29390\
        );

    \I__4986\ : InMux
    port map (
            O => \N__29390\,
            I => \N__29387\
        );

    \I__4985\ : LocalMux
    port map (
            O => \N__29387\,
            I => \N__29384\
        );

    \I__4984\ : Span4Mux_v
    port map (
            O => \N__29384\,
            I => \N__29381\
        );

    \I__4983\ : Odrv4
    port map (
            O => \N__29381\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt18\
        );

    \I__4982\ : InMux
    port map (
            O => \N__29378\,
            I => \N__29372\
        );

    \I__4981\ : InMux
    port map (
            O => \N__29377\,
            I => \N__29372\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__29372\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\
        );

    \I__4979\ : InMux
    port map (
            O => \N__29369\,
            I => \N__29363\
        );

    \I__4978\ : InMux
    port map (
            O => \N__29368\,
            I => \N__29363\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__29363\,
            I => \N__29359\
        );

    \I__4976\ : InMux
    port map (
            O => \N__29362\,
            I => \N__29356\
        );

    \I__4975\ : Span4Mux_h
    port map (
            O => \N__29359\,
            I => \N__29353\
        );

    \I__4974\ : LocalMux
    port map (
            O => \N__29356\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__4973\ : Odrv4
    port map (
            O => \N__29353\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__4972\ : CascadeMux
    port map (
            O => \N__29348\,
            I => \N__29344\
        );

    \I__4971\ : InMux
    port map (
            O => \N__29347\,
            I => \N__29339\
        );

    \I__4970\ : InMux
    port map (
            O => \N__29344\,
            I => \N__29339\
        );

    \I__4969\ : LocalMux
    port map (
            O => \N__29339\,
            I => \N__29335\
        );

    \I__4968\ : InMux
    port map (
            O => \N__29338\,
            I => \N__29332\
        );

    \I__4967\ : Span12Mux_h
    port map (
            O => \N__29335\,
            I => \N__29329\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__29332\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__4965\ : Odrv12
    port map (
            O => \N__29329\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__4964\ : InMux
    port map (
            O => \N__29324\,
            I => \N__29321\
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__29321\,
            I => \N__29318\
        );

    \I__4962\ : Span4Mux_v
    port map (
            O => \N__29318\,
            I => \N__29315\
        );

    \I__4961\ : Odrv4
    port map (
            O => \N__29315\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\
        );

    \I__4960\ : InMux
    port map (
            O => \N__29312\,
            I => \N__29309\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__29309\,
            I => \N__29304\
        );

    \I__4958\ : InMux
    port map (
            O => \N__29308\,
            I => \N__29301\
        );

    \I__4957\ : InMux
    port map (
            O => \N__29307\,
            I => \N__29298\
        );

    \I__4956\ : Span4Mux_v
    port map (
            O => \N__29304\,
            I => \N__29293\
        );

    \I__4955\ : LocalMux
    port map (
            O => \N__29301\,
            I => \N__29293\
        );

    \I__4954\ : LocalMux
    port map (
            O => \N__29298\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19\
        );

    \I__4953\ : Odrv4
    port map (
            O => \N__29293\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19\
        );

    \I__4952\ : InMux
    port map (
            O => \N__29288\,
            I => \N__29283\
        );

    \I__4951\ : InMux
    port map (
            O => \N__29287\,
            I => \N__29280\
        );

    \I__4950\ : CascadeMux
    port map (
            O => \N__29286\,
            I => \N__29277\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__29283\,
            I => \N__29274\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__29280\,
            I => \N__29271\
        );

    \I__4947\ : InMux
    port map (
            O => \N__29277\,
            I => \N__29267\
        );

    \I__4946\ : Span4Mux_h
    port map (
            O => \N__29274\,
            I => \N__29264\
        );

    \I__4945\ : Span4Mux_h
    port map (
            O => \N__29271\,
            I => \N__29261\
        );

    \I__4944\ : InMux
    port map (
            O => \N__29270\,
            I => \N__29258\
        );

    \I__4943\ : LocalMux
    port map (
            O => \N__29267\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__4942\ : Odrv4
    port map (
            O => \N__29264\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__4941\ : Odrv4
    port map (
            O => \N__29261\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__29258\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__4939\ : CascadeMux
    port map (
            O => \N__29249\,
            I => \N__29246\
        );

    \I__4938\ : InMux
    port map (
            O => \N__29246\,
            I => \N__29240\
        );

    \I__4937\ : InMux
    port map (
            O => \N__29245\,
            I => \N__29240\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__29240\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\
        );

    \I__4935\ : InMux
    port map (
            O => \N__29237\,
            I => \N__29234\
        );

    \I__4934\ : LocalMux
    port map (
            O => \N__29234\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\
        );

    \I__4933\ : InMux
    port map (
            O => \N__29231\,
            I => \N__29228\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__29228\,
            I => \N__29225\
        );

    \I__4931\ : Span4Mux_h
    port map (
            O => \N__29225\,
            I => \N__29221\
        );

    \I__4930\ : InMux
    port map (
            O => \N__29224\,
            I => \N__29218\
        );

    \I__4929\ : Span4Mux_v
    port map (
            O => \N__29221\,
            I => \N__29212\
        );

    \I__4928\ : LocalMux
    port map (
            O => \N__29218\,
            I => \N__29212\
        );

    \I__4927\ : InMux
    port map (
            O => \N__29217\,
            I => \N__29209\
        );

    \I__4926\ : Span4Mux_h
    port map (
            O => \N__29212\,
            I => \N__29206\
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__29209\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3\
        );

    \I__4924\ : Odrv4
    port map (
            O => \N__29206\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3\
        );

    \I__4923\ : InMux
    port map (
            O => \N__29201\,
            I => \N__29198\
        );

    \I__4922\ : LocalMux
    port map (
            O => \N__29198\,
            I => \N__29194\
        );

    \I__4921\ : InMux
    port map (
            O => \N__29197\,
            I => \N__29191\
        );

    \I__4920\ : Span4Mux_v
    port map (
            O => \N__29194\,
            I => \N__29184\
        );

    \I__4919\ : LocalMux
    port map (
            O => \N__29191\,
            I => \N__29184\
        );

    \I__4918\ : InMux
    port map (
            O => \N__29190\,
            I => \N__29179\
        );

    \I__4917\ : InMux
    port map (
            O => \N__29189\,
            I => \N__29179\
        );

    \I__4916\ : Odrv4
    port map (
            O => \N__29184\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__29179\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__4914\ : InMux
    port map (
            O => \N__29174\,
            I => \N__29171\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__29171\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\
        );

    \I__4912\ : InMux
    port map (
            O => \N__29168\,
            I => \N__29165\
        );

    \I__4911\ : LocalMux
    port map (
            O => \N__29165\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\
        );

    \I__4910\ : InMux
    port map (
            O => \N__29162\,
            I => \N__29156\
        );

    \I__4909\ : InMux
    port map (
            O => \N__29161\,
            I => \N__29156\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__29156\,
            I => \N__29153\
        );

    \I__4907\ : Span4Mux_h
    port map (
            O => \N__29153\,
            I => \N__29150\
        );

    \I__4906\ : Odrv4
    port map (
            O => \N__29150\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_26\
        );

    \I__4905\ : CascadeMux
    port map (
            O => \N__29147\,
            I => \N__29144\
        );

    \I__4904\ : InMux
    port map (
            O => \N__29144\,
            I => \N__29141\
        );

    \I__4903\ : LocalMux
    port map (
            O => \N__29141\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\
        );

    \I__4902\ : CascadeMux
    port map (
            O => \N__29138\,
            I => \elapsed_time_ns_1_RNIU8PBB_0_20_cascade_\
        );

    \I__4901\ : CascadeMux
    port map (
            O => \N__29135\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15_cascade_\
        );

    \I__4900\ : InMux
    port map (
            O => \N__29132\,
            I => \N__29126\
        );

    \I__4899\ : InMux
    port map (
            O => \N__29131\,
            I => \N__29126\
        );

    \I__4898\ : LocalMux
    port map (
            O => \N__29126\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_20\
        );

    \I__4897\ : CascadeMux
    port map (
            O => \N__29123\,
            I => \N__29119\
        );

    \I__4896\ : InMux
    port map (
            O => \N__29122\,
            I => \N__29114\
        );

    \I__4895\ : InMux
    port map (
            O => \N__29119\,
            I => \N__29114\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__29114\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_21\
        );

    \I__4893\ : InMux
    port map (
            O => \N__29111\,
            I => \N__29108\
        );

    \I__4892\ : LocalMux
    port map (
            O => \N__29108\,
            I => \N__29102\
        );

    \I__4891\ : InMux
    port map (
            O => \N__29107\,
            I => \N__29099\
        );

    \I__4890\ : InMux
    port map (
            O => \N__29106\,
            I => \N__29096\
        );

    \I__4889\ : InMux
    port map (
            O => \N__29105\,
            I => \N__29093\
        );

    \I__4888\ : Span4Mux_v
    port map (
            O => \N__29102\,
            I => \N__29090\
        );

    \I__4887\ : LocalMux
    port map (
            O => \N__29099\,
            I => \N__29085\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__29096\,
            I => \N__29085\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__29093\,
            I => \N__29082\
        );

    \I__4884\ : Odrv4
    port map (
            O => \N__29090\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__4883\ : Odrv12
    port map (
            O => \N__29085\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__4882\ : Odrv4
    port map (
            O => \N__29082\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__4881\ : InMux
    port map (
            O => \N__29075\,
            I => \N__29071\
        );

    \I__4880\ : InMux
    port map (
            O => \N__29074\,
            I => \N__29067\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__29071\,
            I => \N__29064\
        );

    \I__4878\ : InMux
    port map (
            O => \N__29070\,
            I => \N__29061\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__29067\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28\
        );

    \I__4876\ : Odrv12
    port map (
            O => \N__29064\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__29061\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28\
        );

    \I__4874\ : InMux
    port map (
            O => \N__29054\,
            I => \N__29048\
        );

    \I__4873\ : InMux
    port map (
            O => \N__29053\,
            I => \N__29048\
        );

    \I__4872\ : LocalMux
    port map (
            O => \N__29048\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_28\
        );

    \I__4871\ : CascadeMux
    port map (
            O => \N__29045\,
            I => \N__29041\
        );

    \I__4870\ : CascadeMux
    port map (
            O => \N__29044\,
            I => \N__29038\
        );

    \I__4869\ : InMux
    port map (
            O => \N__29041\,
            I => \N__29033\
        );

    \I__4868\ : InMux
    port map (
            O => \N__29038\,
            I => \N__29033\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__29033\,
            I => \N__29030\
        );

    \I__4866\ : Odrv4
    port map (
            O => \N__29030\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_29\
        );

    \I__4865\ : InMux
    port map (
            O => \N__29027\,
            I => \N__29022\
        );

    \I__4864\ : InMux
    port map (
            O => \N__29026\,
            I => \N__29019\
        );

    \I__4863\ : InMux
    port map (
            O => \N__29025\,
            I => \N__29016\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__29022\,
            I => \N__29011\
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__29019\,
            I => \N__29011\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__29016\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30\
        );

    \I__4859\ : Odrv4
    port map (
            O => \N__29011\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30\
        );

    \I__4858\ : CascadeMux
    port map (
            O => \N__29006\,
            I => \N__29002\
        );

    \I__4857\ : InMux
    port map (
            O => \N__29005\,
            I => \N__28998\
        );

    \I__4856\ : InMux
    port map (
            O => \N__29002\,
            I => \N__28995\
        );

    \I__4855\ : InMux
    port map (
            O => \N__29001\,
            I => \N__28991\
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__28998\,
            I => \N__28986\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__28995\,
            I => \N__28986\
        );

    \I__4852\ : InMux
    port map (
            O => \N__28994\,
            I => \N__28983\
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__28991\,
            I => \N__28980\
        );

    \I__4850\ : Span4Mux_v
    port map (
            O => \N__28986\,
            I => \N__28977\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__28983\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__4848\ : Odrv12
    port map (
            O => \N__28980\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__4847\ : Odrv4
    port map (
            O => \N__28977\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__4846\ : InMux
    port map (
            O => \N__28970\,
            I => \N__28967\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__28967\,
            I => \N__28963\
        );

    \I__4844\ : InMux
    port map (
            O => \N__28966\,
            I => \N__28959\
        );

    \I__4843\ : Span4Mux_v
    port map (
            O => \N__28963\,
            I => \N__28956\
        );

    \I__4842\ : InMux
    port map (
            O => \N__28962\,
            I => \N__28953\
        );

    \I__4841\ : LocalMux
    port map (
            O => \N__28959\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23\
        );

    \I__4840\ : Odrv4
    port map (
            O => \N__28956\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23\
        );

    \I__4839\ : LocalMux
    port map (
            O => \N__28953\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23\
        );

    \I__4838\ : InMux
    port map (
            O => \N__28946\,
            I => \N__28942\
        );

    \I__4837\ : InMux
    port map (
            O => \N__28945\,
            I => \N__28939\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__28942\,
            I => \N__28935\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__28939\,
            I => \N__28932\
        );

    \I__4834\ : InMux
    port map (
            O => \N__28938\,
            I => \N__28929\
        );

    \I__4833\ : Span4Mux_h
    port map (
            O => \N__28935\,
            I => \N__28925\
        );

    \I__4832\ : Span4Mux_h
    port map (
            O => \N__28932\,
            I => \N__28922\
        );

    \I__4831\ : LocalMux
    port map (
            O => \N__28929\,
            I => \N__28919\
        );

    \I__4830\ : InMux
    port map (
            O => \N__28928\,
            I => \N__28916\
        );

    \I__4829\ : Odrv4
    port map (
            O => \N__28925\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__4828\ : Odrv4
    port map (
            O => \N__28922\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__4827\ : Odrv12
    port map (
            O => \N__28919\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__28916\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__4825\ : InMux
    port map (
            O => \N__28907\,
            I => \N__28903\
        );

    \I__4824\ : InMux
    port map (
            O => \N__28906\,
            I => \N__28899\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__28903\,
            I => \N__28896\
        );

    \I__4822\ : InMux
    port map (
            O => \N__28902\,
            I => \N__28893\
        );

    \I__4821\ : LocalMux
    port map (
            O => \N__28899\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29\
        );

    \I__4820\ : Odrv4
    port map (
            O => \N__28896\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29\
        );

    \I__4819\ : LocalMux
    port map (
            O => \N__28893\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29\
        );

    \I__4818\ : InMux
    port map (
            O => \N__28886\,
            I => \N__28881\
        );

    \I__4817\ : InMux
    port map (
            O => \N__28885\,
            I => \N__28878\
        );

    \I__4816\ : InMux
    port map (
            O => \N__28884\,
            I => \N__28874\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__28881\,
            I => \N__28871\
        );

    \I__4814\ : LocalMux
    port map (
            O => \N__28878\,
            I => \N__28868\
        );

    \I__4813\ : InMux
    port map (
            O => \N__28877\,
            I => \N__28865\
        );

    \I__4812\ : LocalMux
    port map (
            O => \N__28874\,
            I => \N__28862\
        );

    \I__4811\ : Span4Mux_h
    port map (
            O => \N__28871\,
            I => \N__28855\
        );

    \I__4810\ : Span4Mux_h
    port map (
            O => \N__28868\,
            I => \N__28855\
        );

    \I__4809\ : LocalMux
    port map (
            O => \N__28865\,
            I => \N__28855\
        );

    \I__4808\ : Span4Mux_h
    port map (
            O => \N__28862\,
            I => \N__28852\
        );

    \I__4807\ : Span4Mux_v
    port map (
            O => \N__28855\,
            I => \N__28849\
        );

    \I__4806\ : Odrv4
    port map (
            O => \N__28852\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__4805\ : Odrv4
    port map (
            O => \N__28849\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__4804\ : InMux
    port map (
            O => \N__28844\,
            I => \N__28841\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__28841\,
            I => \N__28837\
        );

    \I__4802\ : InMux
    port map (
            O => \N__28840\,
            I => \N__28834\
        );

    \I__4801\ : Odrv4
    port map (
            O => \N__28837\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__28834\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11\
        );

    \I__4799\ : InMux
    port map (
            O => \N__28829\,
            I => \N__28824\
        );

    \I__4798\ : InMux
    port map (
            O => \N__28828\,
            I => \N__28819\
        );

    \I__4797\ : InMux
    port map (
            O => \N__28827\,
            I => \N__28819\
        );

    \I__4796\ : LocalMux
    port map (
            O => \N__28824\,
            I => \N__28815\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__28819\,
            I => \N__28812\
        );

    \I__4794\ : InMux
    port map (
            O => \N__28818\,
            I => \N__28809\
        );

    \I__4793\ : Odrv4
    port map (
            O => \N__28815\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__4792\ : Odrv4
    port map (
            O => \N__28812\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__28809\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__4790\ : CascadeMux
    port map (
            O => \N__28802\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11_cascade_\
        );

    \I__4789\ : InMux
    port map (
            O => \N__28799\,
            I => \N__28796\
        );

    \I__4788\ : LocalMux
    port map (
            O => \N__28796\,
            I => \N__28792\
        );

    \I__4787\ : InMux
    port map (
            O => \N__28795\,
            I => \N__28789\
        );

    \I__4786\ : Odrv4
    port map (
            O => \N__28792\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10\
        );

    \I__4785\ : LocalMux
    port map (
            O => \N__28789\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10\
        );

    \I__4784\ : InMux
    port map (
            O => \N__28784\,
            I => \N__28777\
        );

    \I__4783\ : InMux
    port map (
            O => \N__28783\,
            I => \N__28777\
        );

    \I__4782\ : InMux
    port map (
            O => \N__28782\,
            I => \N__28774\
        );

    \I__4781\ : LocalMux
    port map (
            O => \N__28777\,
            I => \N__28771\
        );

    \I__4780\ : LocalMux
    port map (
            O => \N__28774\,
            I => \N__28767\
        );

    \I__4779\ : Span4Mux_h
    port map (
            O => \N__28771\,
            I => \N__28764\
        );

    \I__4778\ : InMux
    port map (
            O => \N__28770\,
            I => \N__28761\
        );

    \I__4777\ : Odrv4
    port map (
            O => \N__28767\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__4776\ : Odrv4
    port map (
            O => \N__28764\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__28761\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__4774\ : CascadeMux
    port map (
            O => \N__28754\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10_cascade_\
        );

    \I__4773\ : CascadeMux
    port map (
            O => \N__28751\,
            I => \elapsed_time_ns_1_RNILK91B_0_9_cascade_\
        );

    \I__4772\ : InMux
    port map (
            O => \N__28748\,
            I => \N__28744\
        );

    \I__4771\ : InMux
    port map (
            O => \N__28747\,
            I => \N__28741\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__28744\,
            I => \N__28736\
        );

    \I__4769\ : LocalMux
    port map (
            O => \N__28741\,
            I => \N__28733\
        );

    \I__4768\ : InMux
    port map (
            O => \N__28740\,
            I => \N__28728\
        );

    \I__4767\ : InMux
    port map (
            O => \N__28739\,
            I => \N__28728\
        );

    \I__4766\ : Odrv4
    port map (
            O => \N__28736\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__4765\ : Odrv4
    port map (
            O => \N__28733\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__4764\ : LocalMux
    port map (
            O => \N__28728\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__4763\ : InMux
    port map (
            O => \N__28721\,
            I => \N__28716\
        );

    \I__4762\ : InMux
    port map (
            O => \N__28720\,
            I => \N__28713\
        );

    \I__4761\ : InMux
    port map (
            O => \N__28719\,
            I => \N__28710\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__28716\,
            I => \N__28705\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__28713\,
            I => \N__28705\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__28710\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5\
        );

    \I__4757\ : Odrv12
    port map (
            O => \N__28705\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5\
        );

    \I__4756\ : InMux
    port map (
            O => \N__28700\,
            I => \N__28695\
        );

    \I__4755\ : InMux
    port map (
            O => \N__28699\,
            I => \N__28692\
        );

    \I__4754\ : InMux
    port map (
            O => \N__28698\,
            I => \N__28689\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__28695\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__28692\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12\
        );

    \I__4751\ : LocalMux
    port map (
            O => \N__28689\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12\
        );

    \I__4750\ : InMux
    port map (
            O => \N__28682\,
            I => \N__28676\
        );

    \I__4749\ : InMux
    port map (
            O => \N__28681\,
            I => \N__28673\
        );

    \I__4748\ : InMux
    port map (
            O => \N__28680\,
            I => \N__28670\
        );

    \I__4747\ : CascadeMux
    port map (
            O => \N__28679\,
            I => \N__28667\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__28676\,
            I => \N__28664\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__28673\,
            I => \N__28659\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__28670\,
            I => \N__28659\
        );

    \I__4743\ : InMux
    port map (
            O => \N__28667\,
            I => \N__28656\
        );

    \I__4742\ : Span4Mux_v
    port map (
            O => \N__28664\,
            I => \N__28653\
        );

    \I__4741\ : Span4Mux_h
    port map (
            O => \N__28659\,
            I => \N__28650\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__28656\,
            I => \N__28647\
        );

    \I__4739\ : Odrv4
    port map (
            O => \N__28653\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__4738\ : Odrv4
    port map (
            O => \N__28650\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__4737\ : Odrv4
    port map (
            O => \N__28647\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__4736\ : InMux
    port map (
            O => \N__28640\,
            I => \N__28635\
        );

    \I__4735\ : InMux
    port map (
            O => \N__28639\,
            I => \N__28632\
        );

    \I__4734\ : InMux
    port map (
            O => \N__28638\,
            I => \N__28629\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__28635\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22\
        );

    \I__4732\ : LocalMux
    port map (
            O => \N__28632\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22\
        );

    \I__4731\ : LocalMux
    port map (
            O => \N__28629\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22\
        );

    \I__4730\ : CascadeMux
    port map (
            O => \N__28622\,
            I => \N__28619\
        );

    \I__4729\ : InMux
    port map (
            O => \N__28619\,
            I => \N__28614\
        );

    \I__4728\ : InMux
    port map (
            O => \N__28618\,
            I => \N__28611\
        );

    \I__4727\ : InMux
    port map (
            O => \N__28617\,
            I => \N__28608\
        );

    \I__4726\ : LocalMux
    port map (
            O => \N__28614\,
            I => \N__28604\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__28611\,
            I => \N__28599\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__28608\,
            I => \N__28599\
        );

    \I__4723\ : CascadeMux
    port map (
            O => \N__28607\,
            I => \N__28596\
        );

    \I__4722\ : Span4Mux_v
    port map (
            O => \N__28604\,
            I => \N__28593\
        );

    \I__4721\ : Span4Mux_h
    port map (
            O => \N__28599\,
            I => \N__28590\
        );

    \I__4720\ : InMux
    port map (
            O => \N__28596\,
            I => \N__28587\
        );

    \I__4719\ : Odrv4
    port map (
            O => \N__28593\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__4718\ : Odrv4
    port map (
            O => \N__28590\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__4717\ : LocalMux
    port map (
            O => \N__28587\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__4716\ : InMux
    port map (
            O => \N__28580\,
            I => \pwm_generator_inst.un3_threshold_cry_19\
        );

    \I__4715\ : InMux
    port map (
            O => \N__28577\,
            I => \N__28574\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__28574\,
            I => \N__28571\
        );

    \I__4713\ : Span4Mux_h
    port map (
            O => \N__28571\,
            I => \N__28568\
        );

    \I__4712\ : Odrv4
    port map (
            O => \N__28568\,
            I => il_min_comp1_c
        );

    \I__4711\ : InMux
    port map (
            O => \N__28565\,
            I => \N__28562\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__28562\,
            I => \il_min_comp1_D1\
        );

    \I__4709\ : InMux
    port map (
            O => \N__28559\,
            I => \N__28556\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__28556\,
            I => \N__28553\
        );

    \I__4707\ : Span4Mux_v
    port map (
            O => \N__28553\,
            I => \N__28549\
        );

    \I__4706\ : InMux
    port map (
            O => \N__28552\,
            I => \N__28546\
        );

    \I__4705\ : Sp12to4
    port map (
            O => \N__28549\,
            I => \N__28541\
        );

    \I__4704\ : LocalMux
    port map (
            O => \N__28546\,
            I => \N__28541\
        );

    \I__4703\ : Odrv12
    port map (
            O => \N__28541\,
            I => \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\
        );

    \I__4702\ : InMux
    port map (
            O => \N__28538\,
            I => \pwm_generator_inst.un3_threshold_cry_5\
        );

    \I__4701\ : CascadeMux
    port map (
            O => \N__28535\,
            I => \N__28532\
        );

    \I__4700\ : InMux
    port map (
            O => \N__28532\,
            I => \N__28529\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__28529\,
            I => \N__28526\
        );

    \I__4698\ : Span4Mux_v
    port map (
            O => \N__28526\,
            I => \N__28522\
        );

    \I__4697\ : InMux
    port map (
            O => \N__28525\,
            I => \N__28519\
        );

    \I__4696\ : Sp12to4
    port map (
            O => \N__28522\,
            I => \N__28514\
        );

    \I__4695\ : LocalMux
    port map (
            O => \N__28519\,
            I => \N__28514\
        );

    \I__4694\ : Odrv12
    port map (
            O => \N__28514\,
            I => \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\
        );

    \I__4693\ : InMux
    port map (
            O => \N__28511\,
            I => \pwm_generator_inst.un3_threshold_cry_6\
        );

    \I__4692\ : InMux
    port map (
            O => \N__28508\,
            I => \N__28505\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__28505\,
            I => \N__28502\
        );

    \I__4690\ : Span4Mux_h
    port map (
            O => \N__28502\,
            I => \N__28499\
        );

    \I__4689\ : Span4Mux_h
    port map (
            O => \N__28499\,
            I => \N__28496\
        );

    \I__4688\ : Odrv4
    port map (
            O => \N__28496\,
            I => \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11\
        );

    \I__4687\ : InMux
    port map (
            O => \N__28493\,
            I => \bfn_9_27_0_\
        );

    \I__4686\ : InMux
    port map (
            O => \N__28490\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_30\
        );

    \I__4685\ : InMux
    port map (
            O => \N__28487\,
            I => \N__28484\
        );

    \I__4684\ : LocalMux
    port map (
            O => \N__28484\,
            I => \N__28481\
        );

    \I__4683\ : Odrv4
    port map (
            O => \N__28481\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_31\
        );

    \I__4682\ : InMux
    port map (
            O => \N__28478\,
            I => \N__28475\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__28475\,
            I => \N__28472\
        );

    \I__4680\ : Odrv12
    port map (
            O => \N__28472\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_31\
        );

    \I__4679\ : InMux
    port map (
            O => \N__28469\,
            I => \N__28457\
        );

    \I__4678\ : InMux
    port map (
            O => \N__28468\,
            I => \N__28457\
        );

    \I__4677\ : InMux
    port map (
            O => \N__28467\,
            I => \N__28457\
        );

    \I__4676\ : InMux
    port map (
            O => \N__28466\,
            I => \N__28454\
        );

    \I__4675\ : InMux
    port map (
            O => \N__28465\,
            I => \N__28445\
        );

    \I__4674\ : InMux
    port map (
            O => \N__28464\,
            I => \N__28445\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__28457\,
            I => \N__28442\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__28454\,
            I => \N__28439\
        );

    \I__4671\ : InMux
    port map (
            O => \N__28453\,
            I => \N__28430\
        );

    \I__4670\ : InMux
    port map (
            O => \N__28452\,
            I => \N__28430\
        );

    \I__4669\ : InMux
    port map (
            O => \N__28451\,
            I => \N__28430\
        );

    \I__4668\ : InMux
    port map (
            O => \N__28450\,
            I => \N__28430\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__28445\,
            I => \N__28427\
        );

    \I__4666\ : Span4Mux_h
    port map (
            O => \N__28442\,
            I => \N__28422\
        );

    \I__4665\ : Span4Mux_h
    port map (
            O => \N__28439\,
            I => \N__28422\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__28430\,
            I => \N__28419\
        );

    \I__4663\ : Span4Mux_h
    port map (
            O => \N__28427\,
            I => \N__28416\
        );

    \I__4662\ : Span4Mux_h
    port map (
            O => \N__28422\,
            I => \N__28413\
        );

    \I__4661\ : Span4Mux_h
    port map (
            O => \N__28419\,
            I => \N__28410\
        );

    \I__4660\ : Odrv4
    port map (
            O => \N__28416\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__4659\ : Odrv4
    port map (
            O => \N__28413\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__4658\ : Odrv4
    port map (
            O => \N__28410\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__4657\ : InMux
    port map (
            O => \N__28403\,
            I => \N__28400\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__28400\,
            I => \N__28397\
        );

    \I__4655\ : Span4Mux_v
    port map (
            O => \N__28397\,
            I => \N__28394\
        );

    \I__4654\ : Span4Mux_h
    port map (
            O => \N__28394\,
            I => \N__28390\
        );

    \I__4653\ : InMux
    port map (
            O => \N__28393\,
            I => \N__28387\
        );

    \I__4652\ : Span4Mux_h
    port map (
            O => \N__28390\,
            I => \N__28384\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__28387\,
            I => \pwm_generator_inst.un3_threshold\
        );

    \I__4650\ : Odrv4
    port map (
            O => \N__28384\,
            I => \pwm_generator_inst.un3_threshold\
        );

    \I__4649\ : InMux
    port map (
            O => \N__28379\,
            I => \N__28376\
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__28376\,
            I => \N__28373\
        );

    \I__4647\ : Span4Mux_v
    port map (
            O => \N__28373\,
            I => \N__28370\
        );

    \I__4646\ : Sp12to4
    port map (
            O => \N__28370\,
            I => \N__28367\
        );

    \I__4645\ : Odrv12
    port map (
            O => \N__28367\,
            I => \pwm_generator_inst.O_12\
        );

    \I__4644\ : CascadeMux
    port map (
            O => \N__28364\,
            I => \N__28361\
        );

    \I__4643\ : InMux
    port map (
            O => \N__28361\,
            I => \N__28358\
        );

    \I__4642\ : LocalMux
    port map (
            O => \N__28358\,
            I => \N__28354\
        );

    \I__4641\ : InMux
    port map (
            O => \N__28357\,
            I => \N__28351\
        );

    \I__4640\ : Sp12to4
    port map (
            O => \N__28354\,
            I => \N__28348\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__28351\,
            I => \N__28345\
        );

    \I__4638\ : Span12Mux_v
    port map (
            O => \N__28348\,
            I => \N__28340\
        );

    \I__4637\ : Span12Mux_s4_h
    port map (
            O => \N__28345\,
            I => \N__28340\
        );

    \I__4636\ : Odrv12
    port map (
            O => \N__28340\,
            I => \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\
        );

    \I__4635\ : InMux
    port map (
            O => \N__28337\,
            I => \pwm_generator_inst.un3_threshold_cry_0\
        );

    \I__4634\ : InMux
    port map (
            O => \N__28334\,
            I => \N__28331\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__28331\,
            I => \N__28328\
        );

    \I__4632\ : Span4Mux_v
    port map (
            O => \N__28328\,
            I => \N__28325\
        );

    \I__4631\ : Sp12to4
    port map (
            O => \N__28325\,
            I => \N__28322\
        );

    \I__4630\ : Odrv12
    port map (
            O => \N__28322\,
            I => \pwm_generator_inst.O_13\
        );

    \I__4629\ : InMux
    port map (
            O => \N__28319\,
            I => \N__28315\
        );

    \I__4628\ : InMux
    port map (
            O => \N__28318\,
            I => \N__28312\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__28315\,
            I => \N__28309\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__28312\,
            I => \N__28306\
        );

    \I__4625\ : Span12Mux_v
    port map (
            O => \N__28309\,
            I => \N__28301\
        );

    \I__4624\ : Span12Mux_s3_h
    port map (
            O => \N__28306\,
            I => \N__28301\
        );

    \I__4623\ : Odrv12
    port map (
            O => \N__28301\,
            I => \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\
        );

    \I__4622\ : InMux
    port map (
            O => \N__28298\,
            I => \pwm_generator_inst.un3_threshold_cry_1\
        );

    \I__4621\ : InMux
    port map (
            O => \N__28295\,
            I => \N__28292\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__28292\,
            I => \N__28289\
        );

    \I__4619\ : Span4Mux_v
    port map (
            O => \N__28289\,
            I => \N__28286\
        );

    \I__4618\ : Sp12to4
    port map (
            O => \N__28286\,
            I => \N__28283\
        );

    \I__4617\ : Odrv12
    port map (
            O => \N__28283\,
            I => \pwm_generator_inst.O_14\
        );

    \I__4616\ : InMux
    port map (
            O => \N__28280\,
            I => \N__28277\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__28277\,
            I => \N__28274\
        );

    \I__4614\ : Span4Mux_v
    port map (
            O => \N__28274\,
            I => \N__28270\
        );

    \I__4613\ : InMux
    port map (
            O => \N__28273\,
            I => \N__28267\
        );

    \I__4612\ : Sp12to4
    port map (
            O => \N__28270\,
            I => \N__28262\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__28267\,
            I => \N__28262\
        );

    \I__4610\ : Odrv12
    port map (
            O => \N__28262\,
            I => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\
        );

    \I__4609\ : InMux
    port map (
            O => \N__28259\,
            I => \pwm_generator_inst.un3_threshold_cry_2\
        );

    \I__4608\ : InMux
    port map (
            O => \N__28256\,
            I => \N__28252\
        );

    \I__4607\ : InMux
    port map (
            O => \N__28255\,
            I => \N__28249\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__28252\,
            I => \N__28244\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__28249\,
            I => \N__28244\
        );

    \I__4604\ : Span4Mux_h
    port map (
            O => \N__28244\,
            I => \N__28241\
        );

    \I__4603\ : Span4Mux_h
    port map (
            O => \N__28241\,
            I => \N__28238\
        );

    \I__4602\ : Odrv4
    port map (
            O => \N__28238\,
            I => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\
        );

    \I__4601\ : InMux
    port map (
            O => \N__28235\,
            I => \pwm_generator_inst.un3_threshold_cry_3\
        );

    \I__4600\ : InMux
    port map (
            O => \N__28232\,
            I => \N__28229\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__28229\,
            I => \N__28226\
        );

    \I__4598\ : Span4Mux_v
    port map (
            O => \N__28226\,
            I => \N__28222\
        );

    \I__4597\ : InMux
    port map (
            O => \N__28225\,
            I => \N__28219\
        );

    \I__4596\ : Sp12to4
    port map (
            O => \N__28222\,
            I => \N__28214\
        );

    \I__4595\ : LocalMux
    port map (
            O => \N__28219\,
            I => \N__28214\
        );

    \I__4594\ : Odrv12
    port map (
            O => \N__28214\,
            I => \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\
        );

    \I__4593\ : InMux
    port map (
            O => \N__28211\,
            I => \pwm_generator_inst.un3_threshold_cry_4\
        );

    \I__4592\ : InMux
    port map (
            O => \N__28208\,
            I => \N__28205\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__28205\,
            I => \N__28202\
        );

    \I__4590\ : Span4Mux_v
    port map (
            O => \N__28202\,
            I => \N__28198\
        );

    \I__4589\ : InMux
    port map (
            O => \N__28201\,
            I => \N__28195\
        );

    \I__4588\ : Span4Mux_h
    port map (
            O => \N__28198\,
            I => \N__28192\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__28195\,
            I => \N__28189\
        );

    \I__4586\ : Span4Mux_v
    port map (
            O => \N__28192\,
            I => \N__28186\
        );

    \I__4585\ : Span4Mux_h
    port map (
            O => \N__28189\,
            I => \N__28181\
        );

    \I__4584\ : Span4Mux_h
    port map (
            O => \N__28186\,
            I => \N__28181\
        );

    \I__4583\ : Odrv4
    port map (
            O => \N__28181\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_23\
        );

    \I__4582\ : InMux
    port map (
            O => \N__28178\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_22\
        );

    \I__4581\ : InMux
    port map (
            O => \N__28175\,
            I => \N__28172\
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__28172\,
            I => \N__28168\
        );

    \I__4579\ : InMux
    port map (
            O => \N__28171\,
            I => \N__28165\
        );

    \I__4578\ : Span4Mux_v
    port map (
            O => \N__28168\,
            I => \N__28162\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__28165\,
            I => \N__28159\
        );

    \I__4576\ : Sp12to4
    port map (
            O => \N__28162\,
            I => \N__28156\
        );

    \I__4575\ : Span4Mux_h
    port map (
            O => \N__28159\,
            I => \N__28153\
        );

    \I__4574\ : Span12Mux_s9_h
    port map (
            O => \N__28156\,
            I => \N__28150\
        );

    \I__4573\ : Odrv4
    port map (
            O => \N__28153\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_24\
        );

    \I__4572\ : Odrv12
    port map (
            O => \N__28150\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_24\
        );

    \I__4571\ : InMux
    port map (
            O => \N__28145\,
            I => \bfn_9_18_0_\
        );

    \I__4570\ : InMux
    port map (
            O => \N__28142\,
            I => \N__28138\
        );

    \I__4569\ : InMux
    port map (
            O => \N__28141\,
            I => \N__28135\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__28138\,
            I => \N__28132\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__28135\,
            I => \N__28129\
        );

    \I__4566\ : Span4Mux_h
    port map (
            O => \N__28132\,
            I => \N__28126\
        );

    \I__4565\ : Span12Mux_s9_h
    port map (
            O => \N__28129\,
            I => \N__28123\
        );

    \I__4564\ : Odrv4
    port map (
            O => \N__28126\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_25\
        );

    \I__4563\ : Odrv12
    port map (
            O => \N__28123\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_25\
        );

    \I__4562\ : InMux
    port map (
            O => \N__28118\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_24\
        );

    \I__4561\ : InMux
    port map (
            O => \N__28115\,
            I => \N__28112\
        );

    \I__4560\ : LocalMux
    port map (
            O => \N__28112\,
            I => \N__28108\
        );

    \I__4559\ : InMux
    port map (
            O => \N__28111\,
            I => \N__28105\
        );

    \I__4558\ : Span4Mux_v
    port map (
            O => \N__28108\,
            I => \N__28102\
        );

    \I__4557\ : LocalMux
    port map (
            O => \N__28105\,
            I => \N__28099\
        );

    \I__4556\ : Sp12to4
    port map (
            O => \N__28102\,
            I => \N__28096\
        );

    \I__4555\ : Span4Mux_v
    port map (
            O => \N__28099\,
            I => \N__28093\
        );

    \I__4554\ : Span12Mux_s9_h
    port map (
            O => \N__28096\,
            I => \N__28090\
        );

    \I__4553\ : Odrv4
    port map (
            O => \N__28093\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_26\
        );

    \I__4552\ : Odrv12
    port map (
            O => \N__28090\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_26\
        );

    \I__4551\ : InMux
    port map (
            O => \N__28085\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_25\
        );

    \I__4550\ : InMux
    port map (
            O => \N__28082\,
            I => \N__28079\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__28079\,
            I => \N__28076\
        );

    \I__4548\ : Span4Mux_s2_h
    port map (
            O => \N__28076\,
            I => \N__28072\
        );

    \I__4547\ : InMux
    port map (
            O => \N__28075\,
            I => \N__28069\
        );

    \I__4546\ : Sp12to4
    port map (
            O => \N__28072\,
            I => \N__28066\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__28069\,
            I => \N__28061\
        );

    \I__4544\ : Span12Mux_v
    port map (
            O => \N__28066\,
            I => \N__28061\
        );

    \I__4543\ : Odrv12
    port map (
            O => \N__28061\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_27\
        );

    \I__4542\ : InMux
    port map (
            O => \N__28058\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_26\
        );

    \I__4541\ : InMux
    port map (
            O => \N__28055\,
            I => \N__28052\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__28052\,
            I => \N__28049\
        );

    \I__4539\ : Span4Mux_v
    port map (
            O => \N__28049\,
            I => \N__28045\
        );

    \I__4538\ : InMux
    port map (
            O => \N__28048\,
            I => \N__28042\
        );

    \I__4537\ : Sp12to4
    port map (
            O => \N__28045\,
            I => \N__28039\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__28042\,
            I => \N__28036\
        );

    \I__4535\ : Span12Mux_s9_h
    port map (
            O => \N__28039\,
            I => \N__28033\
        );

    \I__4534\ : Odrv12
    port map (
            O => \N__28036\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_28\
        );

    \I__4533\ : Odrv12
    port map (
            O => \N__28033\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_28\
        );

    \I__4532\ : InMux
    port map (
            O => \N__28028\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_27\
        );

    \I__4531\ : InMux
    port map (
            O => \N__28025\,
            I => \N__28021\
        );

    \I__4530\ : InMux
    port map (
            O => \N__28024\,
            I => \N__28018\
        );

    \I__4529\ : LocalMux
    port map (
            O => \N__28021\,
            I => \N__28015\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__28018\,
            I => \N__28012\
        );

    \I__4527\ : Span4Mux_v
    port map (
            O => \N__28015\,
            I => \N__28009\
        );

    \I__4526\ : Span12Mux_v
    port map (
            O => \N__28012\,
            I => \N__28006\
        );

    \I__4525\ : Odrv4
    port map (
            O => \N__28009\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_29\
        );

    \I__4524\ : Odrv12
    port map (
            O => \N__28006\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_29\
        );

    \I__4523\ : InMux
    port map (
            O => \N__28001\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_28\
        );

    \I__4522\ : InMux
    port map (
            O => \N__27998\,
            I => \N__27995\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__27995\,
            I => \N__27992\
        );

    \I__4520\ : Span4Mux_v
    port map (
            O => \N__27992\,
            I => \N__27988\
        );

    \I__4519\ : InMux
    port map (
            O => \N__27991\,
            I => \N__27985\
        );

    \I__4518\ : Span4Mux_v
    port map (
            O => \N__27988\,
            I => \N__27982\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__27985\,
            I => \N__27979\
        );

    \I__4516\ : Span4Mux_v
    port map (
            O => \N__27982\,
            I => \N__27976\
        );

    \I__4515\ : Span4Mux_h
    port map (
            O => \N__27979\,
            I => \N__27973\
        );

    \I__4514\ : Sp12to4
    port map (
            O => \N__27976\,
            I => \N__27970\
        );

    \I__4513\ : Odrv4
    port map (
            O => \N__27973\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_30\
        );

    \I__4512\ : Odrv12
    port map (
            O => \N__27970\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_30\
        );

    \I__4511\ : InMux
    port map (
            O => \N__27965\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_29\
        );

    \I__4510\ : InMux
    port map (
            O => \N__27962\,
            I => \N__27959\
        );

    \I__4509\ : LocalMux
    port map (
            O => \N__27959\,
            I => \N__27956\
        );

    \I__4508\ : Span4Mux_v
    port map (
            O => \N__27956\,
            I => \N__27952\
        );

    \I__4507\ : InMux
    port map (
            O => \N__27955\,
            I => \N__27949\
        );

    \I__4506\ : Span4Mux_v
    port map (
            O => \N__27952\,
            I => \N__27946\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__27949\,
            I => \N__27943\
        );

    \I__4504\ : Span4Mux_h
    port map (
            O => \N__27946\,
            I => \N__27940\
        );

    \I__4503\ : Span4Mux_h
    port map (
            O => \N__27943\,
            I => \N__27935\
        );

    \I__4502\ : Span4Mux_h
    port map (
            O => \N__27940\,
            I => \N__27935\
        );

    \I__4501\ : Odrv4
    port map (
            O => \N__27935\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_15\
        );

    \I__4500\ : InMux
    port map (
            O => \N__27932\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_14\
        );

    \I__4499\ : InMux
    port map (
            O => \N__27929\,
            I => \N__27926\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__27926\,
            I => \N__27923\
        );

    \I__4497\ : Span4Mux_v
    port map (
            O => \N__27923\,
            I => \N__27919\
        );

    \I__4496\ : InMux
    port map (
            O => \N__27922\,
            I => \N__27916\
        );

    \I__4495\ : Sp12to4
    port map (
            O => \N__27919\,
            I => \N__27913\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__27916\,
            I => \N__27910\
        );

    \I__4493\ : Span12Mux_s9_h
    port map (
            O => \N__27913\,
            I => \N__27907\
        );

    \I__4492\ : Odrv12
    port map (
            O => \N__27910\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_16\
        );

    \I__4491\ : Odrv12
    port map (
            O => \N__27907\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_16\
        );

    \I__4490\ : InMux
    port map (
            O => \N__27902\,
            I => \bfn_9_17_0_\
        );

    \I__4489\ : InMux
    port map (
            O => \N__27899\,
            I => \N__27896\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__27896\,
            I => \N__27893\
        );

    \I__4487\ : Span4Mux_v
    port map (
            O => \N__27893\,
            I => \N__27889\
        );

    \I__4486\ : InMux
    port map (
            O => \N__27892\,
            I => \N__27886\
        );

    \I__4485\ : Span4Mux_v
    port map (
            O => \N__27889\,
            I => \N__27883\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__27886\,
            I => \N__27880\
        );

    \I__4483\ : Span4Mux_h
    port map (
            O => \N__27883\,
            I => \N__27877\
        );

    \I__4482\ : Span4Mux_h
    port map (
            O => \N__27880\,
            I => \N__27874\
        );

    \I__4481\ : Span4Mux_h
    port map (
            O => \N__27877\,
            I => \N__27871\
        );

    \I__4480\ : Odrv4
    port map (
            O => \N__27874\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_17\
        );

    \I__4479\ : Odrv4
    port map (
            O => \N__27871\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_17\
        );

    \I__4478\ : InMux
    port map (
            O => \N__27866\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_16\
        );

    \I__4477\ : InMux
    port map (
            O => \N__27863\,
            I => \N__27860\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__27860\,
            I => \N__27856\
        );

    \I__4475\ : InMux
    port map (
            O => \N__27859\,
            I => \N__27853\
        );

    \I__4474\ : Span4Mux_h
    port map (
            O => \N__27856\,
            I => \N__27850\
        );

    \I__4473\ : LocalMux
    port map (
            O => \N__27853\,
            I => \N__27847\
        );

    \I__4472\ : Span4Mux_h
    port map (
            O => \N__27850\,
            I => \N__27844\
        );

    \I__4471\ : Span12Mux_s9_h
    port map (
            O => \N__27847\,
            I => \N__27841\
        );

    \I__4470\ : Odrv4
    port map (
            O => \N__27844\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_18\
        );

    \I__4469\ : Odrv12
    port map (
            O => \N__27841\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_18\
        );

    \I__4468\ : InMux
    port map (
            O => \N__27836\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_17\
        );

    \I__4467\ : InMux
    port map (
            O => \N__27833\,
            I => \N__27830\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__27830\,
            I => \N__27827\
        );

    \I__4465\ : Span4Mux_v
    port map (
            O => \N__27827\,
            I => \N__27823\
        );

    \I__4464\ : InMux
    port map (
            O => \N__27826\,
            I => \N__27820\
        );

    \I__4463\ : Span4Mux_h
    port map (
            O => \N__27823\,
            I => \N__27817\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__27820\,
            I => \N__27814\
        );

    \I__4461\ : Span4Mux_v
    port map (
            O => \N__27817\,
            I => \N__27811\
        );

    \I__4460\ : Span4Mux_h
    port map (
            O => \N__27814\,
            I => \N__27806\
        );

    \I__4459\ : Span4Mux_h
    port map (
            O => \N__27811\,
            I => \N__27806\
        );

    \I__4458\ : Odrv4
    port map (
            O => \N__27806\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_19\
        );

    \I__4457\ : InMux
    port map (
            O => \N__27803\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_18\
        );

    \I__4456\ : InMux
    port map (
            O => \N__27800\,
            I => \N__27796\
        );

    \I__4455\ : InMux
    port map (
            O => \N__27799\,
            I => \N__27793\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__27796\,
            I => \N__27790\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__27793\,
            I => \N__27787\
        );

    \I__4452\ : Span4Mux_v
    port map (
            O => \N__27790\,
            I => \N__27784\
        );

    \I__4451\ : Span4Mux_h
    port map (
            O => \N__27787\,
            I => \N__27781\
        );

    \I__4450\ : Sp12to4
    port map (
            O => \N__27784\,
            I => \N__27778\
        );

    \I__4449\ : Span4Mux_h
    port map (
            O => \N__27781\,
            I => \N__27775\
        );

    \I__4448\ : Span12Mux_s9_h
    port map (
            O => \N__27778\,
            I => \N__27772\
        );

    \I__4447\ : Odrv4
    port map (
            O => \N__27775\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_20\
        );

    \I__4446\ : Odrv12
    port map (
            O => \N__27772\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_20\
        );

    \I__4445\ : InMux
    port map (
            O => \N__27767\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_19\
        );

    \I__4444\ : InMux
    port map (
            O => \N__27764\,
            I => \N__27760\
        );

    \I__4443\ : InMux
    port map (
            O => \N__27763\,
            I => \N__27757\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__27760\,
            I => \N__27754\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__27757\,
            I => \N__27751\
        );

    \I__4440\ : Span4Mux_v
    port map (
            O => \N__27754\,
            I => \N__27748\
        );

    \I__4439\ : Span12Mux_v
    port map (
            O => \N__27751\,
            I => \N__27745\
        );

    \I__4438\ : Odrv4
    port map (
            O => \N__27748\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_21\
        );

    \I__4437\ : Odrv12
    port map (
            O => \N__27745\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_21\
        );

    \I__4436\ : InMux
    port map (
            O => \N__27740\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_20\
        );

    \I__4435\ : InMux
    port map (
            O => \N__27737\,
            I => \N__27734\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__27734\,
            I => \N__27730\
        );

    \I__4433\ : InMux
    port map (
            O => \N__27733\,
            I => \N__27727\
        );

    \I__4432\ : Span4Mux_v
    port map (
            O => \N__27730\,
            I => \N__27724\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__27727\,
            I => \N__27721\
        );

    \I__4430\ : Span4Mux_v
    port map (
            O => \N__27724\,
            I => \N__27718\
        );

    \I__4429\ : Span4Mux_v
    port map (
            O => \N__27721\,
            I => \N__27713\
        );

    \I__4428\ : Span4Mux_h
    port map (
            O => \N__27718\,
            I => \N__27713\
        );

    \I__4427\ : Span4Mux_h
    port map (
            O => \N__27713\,
            I => \N__27710\
        );

    \I__4426\ : Odrv4
    port map (
            O => \N__27710\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_22\
        );

    \I__4425\ : InMux
    port map (
            O => \N__27707\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_21\
        );

    \I__4424\ : InMux
    port map (
            O => \N__27704\,
            I => \N__27701\
        );

    \I__4423\ : LocalMux
    port map (
            O => \N__27701\,
            I => \N__27697\
        );

    \I__4422\ : InMux
    port map (
            O => \N__27700\,
            I => \N__27694\
        );

    \I__4421\ : Span4Mux_v
    port map (
            O => \N__27697\,
            I => \N__27691\
        );

    \I__4420\ : LocalMux
    port map (
            O => \N__27694\,
            I => \N__27686\
        );

    \I__4419\ : Sp12to4
    port map (
            O => \N__27691\,
            I => \N__27686\
        );

    \I__4418\ : Odrv12
    port map (
            O => \N__27686\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__4417\ : InMux
    port map (
            O => \N__27683\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_5\
        );

    \I__4416\ : InMux
    port map (
            O => \N__27680\,
            I => \N__27677\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__27677\,
            I => \N__27674\
        );

    \I__4414\ : Span4Mux_s2_h
    port map (
            O => \N__27674\,
            I => \N__27670\
        );

    \I__4413\ : InMux
    port map (
            O => \N__27673\,
            I => \N__27667\
        );

    \I__4412\ : Span4Mux_h
    port map (
            O => \N__27670\,
            I => \N__27664\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__27667\,
            I => \N__27661\
        );

    \I__4410\ : Span4Mux_h
    port map (
            O => \N__27664\,
            I => \N__27658\
        );

    \I__4409\ : Odrv12
    port map (
            O => \N__27661\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__4408\ : Odrv4
    port map (
            O => \N__27658\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__4407\ : InMux
    port map (
            O => \N__27653\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_6\
        );

    \I__4406\ : InMux
    port map (
            O => \N__27650\,
            I => \N__27646\
        );

    \I__4405\ : InMux
    port map (
            O => \N__27649\,
            I => \N__27643\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__27646\,
            I => \N__27640\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__27643\,
            I => \N__27637\
        );

    \I__4402\ : Span12Mux_s9_h
    port map (
            O => \N__27640\,
            I => \N__27634\
        );

    \I__4401\ : Odrv12
    port map (
            O => \N__27637\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__4400\ : Odrv12
    port map (
            O => \N__27634\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__4399\ : InMux
    port map (
            O => \N__27629\,
            I => \bfn_9_16_0_\
        );

    \I__4398\ : InMux
    port map (
            O => \N__27626\,
            I => \N__27623\
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__27623\,
            I => \N__27619\
        );

    \I__4396\ : InMux
    port map (
            O => \N__27622\,
            I => \N__27616\
        );

    \I__4395\ : Span4Mux_s1_h
    port map (
            O => \N__27619\,
            I => \N__27613\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__27616\,
            I => \N__27610\
        );

    \I__4393\ : Span4Mux_h
    port map (
            O => \N__27613\,
            I => \N__27607\
        );

    \I__4392\ : Span4Mux_h
    port map (
            O => \N__27610\,
            I => \N__27604\
        );

    \I__4391\ : Span4Mux_h
    port map (
            O => \N__27607\,
            I => \N__27601\
        );

    \I__4390\ : Odrv4
    port map (
            O => \N__27604\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__4389\ : Odrv4
    port map (
            O => \N__27601\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__4388\ : InMux
    port map (
            O => \N__27596\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_8\
        );

    \I__4387\ : InMux
    port map (
            O => \N__27593\,
            I => \N__27589\
        );

    \I__4386\ : InMux
    port map (
            O => \N__27592\,
            I => \N__27586\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__27589\,
            I => \N__27583\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__27586\,
            I => \N__27580\
        );

    \I__4383\ : Span4Mux_s2_h
    port map (
            O => \N__27583\,
            I => \N__27577\
        );

    \I__4382\ : Span4Mux_h
    port map (
            O => \N__27580\,
            I => \N__27574\
        );

    \I__4381\ : Span4Mux_h
    port map (
            O => \N__27577\,
            I => \N__27571\
        );

    \I__4380\ : Span4Mux_h
    port map (
            O => \N__27574\,
            I => \N__27568\
        );

    \I__4379\ : Span4Mux_h
    port map (
            O => \N__27571\,
            I => \N__27565\
        );

    \I__4378\ : Odrv4
    port map (
            O => \N__27568\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__4377\ : Odrv4
    port map (
            O => \N__27565\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__4376\ : InMux
    port map (
            O => \N__27560\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_9\
        );

    \I__4375\ : InMux
    port map (
            O => \N__27557\,
            I => \N__27554\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__27554\,
            I => \N__27551\
        );

    \I__4373\ : Span4Mux_s2_h
    port map (
            O => \N__27551\,
            I => \N__27547\
        );

    \I__4372\ : InMux
    port map (
            O => \N__27550\,
            I => \N__27544\
        );

    \I__4371\ : Span4Mux_h
    port map (
            O => \N__27547\,
            I => \N__27541\
        );

    \I__4370\ : LocalMux
    port map (
            O => \N__27544\,
            I => \N__27538\
        );

    \I__4369\ : Span4Mux_h
    port map (
            O => \N__27541\,
            I => \N__27535\
        );

    \I__4368\ : Odrv12
    port map (
            O => \N__27538\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__4367\ : Odrv4
    port map (
            O => \N__27535\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__4366\ : InMux
    port map (
            O => \N__27530\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_10\
        );

    \I__4365\ : InMux
    port map (
            O => \N__27527\,
            I => \N__27524\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__27524\,
            I => \N__27521\
        );

    \I__4363\ : Span4Mux_s1_h
    port map (
            O => \N__27521\,
            I => \N__27517\
        );

    \I__4362\ : InMux
    port map (
            O => \N__27520\,
            I => \N__27514\
        );

    \I__4361\ : Span4Mux_h
    port map (
            O => \N__27517\,
            I => \N__27511\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__27514\,
            I => \N__27508\
        );

    \I__4359\ : Span4Mux_h
    port map (
            O => \N__27511\,
            I => \N__27505\
        );

    \I__4358\ : Odrv12
    port map (
            O => \N__27508\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__4357\ : Odrv4
    port map (
            O => \N__27505\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__4356\ : InMux
    port map (
            O => \N__27500\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_11\
        );

    \I__4355\ : InMux
    port map (
            O => \N__27497\,
            I => \N__27494\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__27494\,
            I => \N__27490\
        );

    \I__4353\ : InMux
    port map (
            O => \N__27493\,
            I => \N__27487\
        );

    \I__4352\ : Span4Mux_v
    port map (
            O => \N__27490\,
            I => \N__27484\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__27487\,
            I => \N__27481\
        );

    \I__4350\ : Sp12to4
    port map (
            O => \N__27484\,
            I => \N__27476\
        );

    \I__4349\ : Span12Mux_v
    port map (
            O => \N__27481\,
            I => \N__27476\
        );

    \I__4348\ : Odrv12
    port map (
            O => \N__27476\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_13\
        );

    \I__4347\ : InMux
    port map (
            O => \N__27473\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_12\
        );

    \I__4346\ : InMux
    port map (
            O => \N__27470\,
            I => \N__27467\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__27467\,
            I => \N__27463\
        );

    \I__4344\ : InMux
    port map (
            O => \N__27466\,
            I => \N__27460\
        );

    \I__4343\ : Span4Mux_s2_h
    port map (
            O => \N__27463\,
            I => \N__27457\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__27460\,
            I => \N__27454\
        );

    \I__4341\ : Span4Mux_v
    port map (
            O => \N__27457\,
            I => \N__27451\
        );

    \I__4340\ : Span4Mux_v
    port map (
            O => \N__27454\,
            I => \N__27446\
        );

    \I__4339\ : Span4Mux_h
    port map (
            O => \N__27451\,
            I => \N__27446\
        );

    \I__4338\ : Odrv4
    port map (
            O => \N__27446\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__4337\ : InMux
    port map (
            O => \N__27443\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_13\
        );

    \I__4336\ : InMux
    port map (
            O => \N__27440\,
            I => \N__27437\
        );

    \I__4335\ : LocalMux
    port map (
            O => \N__27437\,
            I => \N__27434\
        );

    \I__4334\ : Odrv4
    port map (
            O => \N__27434\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\
        );

    \I__4333\ : CascadeMux
    port map (
            O => \N__27431\,
            I => \N__27428\
        );

    \I__4332\ : InMux
    port map (
            O => \N__27428\,
            I => \N__27425\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__27425\,
            I => \N__27422\
        );

    \I__4330\ : Span4Mux_v
    port map (
            O => \N__27422\,
            I => \N__27419\
        );

    \I__4329\ : Odrv4
    port map (
            O => \N__27419\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt30\
        );

    \I__4328\ : InMux
    port map (
            O => \N__27416\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_30\
        );

    \I__4327\ : InMux
    port map (
            O => \N__27413\,
            I => \N__27410\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__27410\,
            I => \N__27405\
        );

    \I__4325\ : InMux
    port map (
            O => \N__27409\,
            I => \N__27400\
        );

    \I__4324\ : InMux
    port map (
            O => \N__27408\,
            I => \N__27400\
        );

    \I__4323\ : Span4Mux_h
    port map (
            O => \N__27405\,
            I => \N__27397\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__27400\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__4321\ : Odrv4
    port map (
            O => \N__27397\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__4320\ : InMux
    port map (
            O => \N__27392\,
            I => \N__27389\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__27389\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axb_0\
        );

    \I__4318\ : InMux
    port map (
            O => \N__27386\,
            I => \N__27382\
        );

    \I__4317\ : InMux
    port map (
            O => \N__27385\,
            I => \N__27379\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__27382\,
            I => \N__27376\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__27379\,
            I => \N__27373\
        );

    \I__4314\ : Span4Mux_h
    port map (
            O => \N__27376\,
            I => \N__27370\
        );

    \I__4313\ : Span12Mux_s9_h
    port map (
            O => \N__27373\,
            I => \N__27367\
        );

    \I__4312\ : Odrv4
    port map (
            O => \N__27370\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_1\
        );

    \I__4311\ : Odrv12
    port map (
            O => \N__27367\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_1\
        );

    \I__4310\ : InMux
    port map (
            O => \N__27362\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_0\
        );

    \I__4309\ : InMux
    port map (
            O => \N__27359\,
            I => \N__27356\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__27356\,
            I => \N__27353\
        );

    \I__4307\ : Span4Mux_s1_h
    port map (
            O => \N__27353\,
            I => \N__27349\
        );

    \I__4306\ : InMux
    port map (
            O => \N__27352\,
            I => \N__27346\
        );

    \I__4305\ : Span4Mux_h
    port map (
            O => \N__27349\,
            I => \N__27343\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__27346\,
            I => \N__27340\
        );

    \I__4303\ : Span4Mux_h
    port map (
            O => \N__27343\,
            I => \N__27337\
        );

    \I__4302\ : Odrv12
    port map (
            O => \N__27340\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__4301\ : Odrv4
    port map (
            O => \N__27337\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__4300\ : InMux
    port map (
            O => \N__27332\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_1\
        );

    \I__4299\ : InMux
    port map (
            O => \N__27329\,
            I => \N__27325\
        );

    \I__4298\ : InMux
    port map (
            O => \N__27328\,
            I => \N__27322\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__27325\,
            I => \N__27319\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__27322\,
            I => \N__27316\
        );

    \I__4295\ : Span4Mux_s1_h
    port map (
            O => \N__27319\,
            I => \N__27313\
        );

    \I__4294\ : Span4Mux_v
    port map (
            O => \N__27316\,
            I => \N__27308\
        );

    \I__4293\ : Span4Mux_h
    port map (
            O => \N__27313\,
            I => \N__27308\
        );

    \I__4292\ : Span4Mux_h
    port map (
            O => \N__27308\,
            I => \N__27305\
        );

    \I__4291\ : Odrv4
    port map (
            O => \N__27305\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__4290\ : InMux
    port map (
            O => \N__27302\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_2\
        );

    \I__4289\ : InMux
    port map (
            O => \N__27299\,
            I => \N__27296\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__27296\,
            I => \N__27292\
        );

    \I__4287\ : InMux
    port map (
            O => \N__27295\,
            I => \N__27289\
        );

    \I__4286\ : Span4Mux_v
    port map (
            O => \N__27292\,
            I => \N__27286\
        );

    \I__4285\ : LocalMux
    port map (
            O => \N__27289\,
            I => \N__27281\
        );

    \I__4284\ : Sp12to4
    port map (
            O => \N__27286\,
            I => \N__27281\
        );

    \I__4283\ : Odrv12
    port map (
            O => \N__27281\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__4282\ : InMux
    port map (
            O => \N__27278\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_3\
        );

    \I__4281\ : InMux
    port map (
            O => \N__27275\,
            I => \N__27272\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__27272\,
            I => \N__27268\
        );

    \I__4279\ : InMux
    port map (
            O => \N__27271\,
            I => \N__27265\
        );

    \I__4278\ : Span4Mux_v
    port map (
            O => \N__27268\,
            I => \N__27262\
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__27265\,
            I => \N__27259\
        );

    \I__4276\ : Sp12to4
    port map (
            O => \N__27262\,
            I => \N__27254\
        );

    \I__4275\ : Span12Mux_v
    port map (
            O => \N__27259\,
            I => \N__27254\
        );

    \I__4274\ : Odrv12
    port map (
            O => \N__27254\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__4273\ : InMux
    port map (
            O => \N__27251\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_4\
        );

    \I__4272\ : InMux
    port map (
            O => \N__27248\,
            I => \N__27244\
        );

    \I__4271\ : InMux
    port map (
            O => \N__27247\,
            I => \N__27241\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__27244\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__27241\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__4268\ : InMux
    port map (
            O => \N__27236\,
            I => \N__27233\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__27233\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\
        );

    \I__4266\ : InMux
    port map (
            O => \N__27230\,
            I => \N__27227\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__27227\,
            I => \N__27224\
        );

    \I__4264\ : Odrv12
    port map (
            O => \N__27224\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22\
        );

    \I__4263\ : CascadeMux
    port map (
            O => \N__27221\,
            I => \N__27218\
        );

    \I__4262\ : InMux
    port map (
            O => \N__27218\,
            I => \N__27215\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__27215\,
            I => \N__27212\
        );

    \I__4260\ : Odrv12
    port map (
            O => \N__27212\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt22\
        );

    \I__4259\ : InMux
    port map (
            O => \N__27209\,
            I => \N__27206\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__27206\,
            I => \N__27203\
        );

    \I__4257\ : Odrv12
    port map (
            O => \N__27203\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24\
        );

    \I__4256\ : CascadeMux
    port map (
            O => \N__27200\,
            I => \N__27197\
        );

    \I__4255\ : InMux
    port map (
            O => \N__27197\,
            I => \N__27194\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__27194\,
            I => \N__27191\
        );

    \I__4253\ : Span4Mux_v
    port map (
            O => \N__27191\,
            I => \N__27188\
        );

    \I__4252\ : Odrv4
    port map (
            O => \N__27188\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt24\
        );

    \I__4251\ : InMux
    port map (
            O => \N__27185\,
            I => \N__27182\
        );

    \I__4250\ : LocalMux
    port map (
            O => \N__27182\,
            I => \N__27179\
        );

    \I__4249\ : Odrv4
    port map (
            O => \N__27179\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt26\
        );

    \I__4248\ : CascadeMux
    port map (
            O => \N__27176\,
            I => \N__27173\
        );

    \I__4247\ : InMux
    port map (
            O => \N__27173\,
            I => \N__27170\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__27170\,
            I => \N__27167\
        );

    \I__4245\ : Odrv4
    port map (
            O => \N__27167\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26\
        );

    \I__4244\ : InMux
    port map (
            O => \N__27164\,
            I => \N__27161\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__27161\,
            I => \N__27158\
        );

    \I__4242\ : Span4Mux_h
    port map (
            O => \N__27158\,
            I => \N__27155\
        );

    \I__4241\ : Odrv4
    port map (
            O => \N__27155\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt28\
        );

    \I__4240\ : CascadeMux
    port map (
            O => \N__27152\,
            I => \N__27149\
        );

    \I__4239\ : InMux
    port map (
            O => \N__27149\,
            I => \N__27146\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__27146\,
            I => \N__27143\
        );

    \I__4237\ : Span4Mux_h
    port map (
            O => \N__27143\,
            I => \N__27140\
        );

    \I__4236\ : Odrv4
    port map (
            O => \N__27140\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28\
        );

    \I__4235\ : InMux
    port map (
            O => \N__27137\,
            I => \N__27134\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__27134\,
            I => \N__27131\
        );

    \I__4233\ : Odrv4
    port map (
            O => \N__27131\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\
        );

    \I__4232\ : InMux
    port map (
            O => \N__27128\,
            I => \N__27124\
        );

    \I__4231\ : InMux
    port map (
            O => \N__27127\,
            I => \N__27121\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__27124\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__4229\ : LocalMux
    port map (
            O => \N__27121\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__4228\ : CascadeMux
    port map (
            O => \N__27116\,
            I => \N__27113\
        );

    \I__4227\ : InMux
    port map (
            O => \N__27113\,
            I => \N__27110\
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__27110\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\
        );

    \I__4225\ : InMux
    port map (
            O => \N__27107\,
            I => \N__27103\
        );

    \I__4224\ : InMux
    port map (
            O => \N__27106\,
            I => \N__27100\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__27103\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__27100\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__4221\ : InMux
    port map (
            O => \N__27095\,
            I => \N__27092\
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__27092\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\
        );

    \I__4219\ : InMux
    port map (
            O => \N__27089\,
            I => \N__27085\
        );

    \I__4218\ : InMux
    port map (
            O => \N__27088\,
            I => \N__27082\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__27085\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__4216\ : LocalMux
    port map (
            O => \N__27082\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__4215\ : InMux
    port map (
            O => \N__27077\,
            I => \N__27074\
        );

    \I__4214\ : LocalMux
    port map (
            O => \N__27074\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\
        );

    \I__4213\ : InMux
    port map (
            O => \N__27071\,
            I => \N__27068\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__27068\,
            I => \N__27065\
        );

    \I__4211\ : Odrv4
    port map (
            O => \N__27065\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\
        );

    \I__4210\ : InMux
    port map (
            O => \N__27062\,
            I => \N__27059\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__27059\,
            I => \N__27055\
        );

    \I__4208\ : InMux
    port map (
            O => \N__27058\,
            I => \N__27052\
        );

    \I__4207\ : Span4Mux_v
    port map (
            O => \N__27055\,
            I => \N__27049\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__27052\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__4205\ : Odrv4
    port map (
            O => \N__27049\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__4204\ : CascadeMux
    port map (
            O => \N__27044\,
            I => \N__27041\
        );

    \I__4203\ : InMux
    port map (
            O => \N__27041\,
            I => \N__27038\
        );

    \I__4202\ : LocalMux
    port map (
            O => \N__27038\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\
        );

    \I__4201\ : InMux
    port map (
            O => \N__27035\,
            I => \N__27032\
        );

    \I__4200\ : LocalMux
    port map (
            O => \N__27032\,
            I => \N__27029\
        );

    \I__4199\ : Odrv4
    port map (
            O => \N__27029\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\
        );

    \I__4198\ : InMux
    port map (
            O => \N__27026\,
            I => \N__27022\
        );

    \I__4197\ : InMux
    port map (
            O => \N__27025\,
            I => \N__27019\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__27022\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__4195\ : LocalMux
    port map (
            O => \N__27019\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__4194\ : CascadeMux
    port map (
            O => \N__27014\,
            I => \N__27011\
        );

    \I__4193\ : InMux
    port map (
            O => \N__27011\,
            I => \N__27008\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__27008\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\
        );

    \I__4191\ : CascadeMux
    port map (
            O => \N__27005\,
            I => \N__27002\
        );

    \I__4190\ : InMux
    port map (
            O => \N__27002\,
            I => \N__26999\
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__26999\,
            I => \N__26996\
        );

    \I__4188\ : Odrv12
    port map (
            O => \N__26996\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\
        );

    \I__4187\ : InMux
    port map (
            O => \N__26993\,
            I => \N__26989\
        );

    \I__4186\ : InMux
    port map (
            O => \N__26992\,
            I => \N__26986\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__26989\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__26986\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__4183\ : InMux
    port map (
            O => \N__26981\,
            I => \N__26978\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__26978\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\
        );

    \I__4181\ : InMux
    port map (
            O => \N__26975\,
            I => \N__26971\
        );

    \I__4180\ : InMux
    port map (
            O => \N__26974\,
            I => \N__26968\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__26971\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__26968\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__4177\ : CascadeMux
    port map (
            O => \N__26963\,
            I => \N__26960\
        );

    \I__4176\ : InMux
    port map (
            O => \N__26960\,
            I => \N__26957\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__26957\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\
        );

    \I__4174\ : CascadeMux
    port map (
            O => \N__26954\,
            I => \N__26951\
        );

    \I__4173\ : InMux
    port map (
            O => \N__26951\,
            I => \N__26948\
        );

    \I__4172\ : LocalMux
    port map (
            O => \N__26948\,
            I => \N__26945\
        );

    \I__4171\ : Odrv4
    port map (
            O => \N__26945\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\
        );

    \I__4170\ : InMux
    port map (
            O => \N__26942\,
            I => \N__26938\
        );

    \I__4169\ : InMux
    port map (
            O => \N__26941\,
            I => \N__26935\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__26938\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__26935\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__4166\ : InMux
    port map (
            O => \N__26930\,
            I => \N__26927\
        );

    \I__4165\ : LocalMux
    port map (
            O => \N__26927\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\
        );

    \I__4164\ : InMux
    port map (
            O => \N__26924\,
            I => \N__26917\
        );

    \I__4163\ : InMux
    port map (
            O => \N__26923\,
            I => \N__26917\
        );

    \I__4162\ : InMux
    port map (
            O => \N__26922\,
            I => \N__26914\
        );

    \I__4161\ : LocalMux
    port map (
            O => \N__26917\,
            I => \N__26911\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__26914\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__4159\ : Odrv4
    port map (
            O => \N__26911\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__4158\ : CascadeMux
    port map (
            O => \N__26906\,
            I => \N__26902\
        );

    \I__4157\ : InMux
    port map (
            O => \N__26905\,
            I => \N__26897\
        );

    \I__4156\ : InMux
    port map (
            O => \N__26902\,
            I => \N__26897\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__26897\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_30\
        );

    \I__4154\ : CascadeMux
    port map (
            O => \N__26894\,
            I => \N__26890\
        );

    \I__4153\ : InMux
    port map (
            O => \N__26893\,
            I => \N__26885\
        );

    \I__4152\ : InMux
    port map (
            O => \N__26890\,
            I => \N__26885\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__26885\,
            I => \N__26881\
        );

    \I__4150\ : InMux
    port map (
            O => \N__26884\,
            I => \N__26878\
        );

    \I__4149\ : Span4Mux_h
    port map (
            O => \N__26881\,
            I => \N__26875\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__26878\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__4147\ : Odrv4
    port map (
            O => \N__26875\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__4146\ : InMux
    port map (
            O => \N__26870\,
            I => \N__26864\
        );

    \I__4145\ : InMux
    port map (
            O => \N__26869\,
            I => \N__26864\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__26864\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_31\
        );

    \I__4143\ : CascadeMux
    port map (
            O => \N__26861\,
            I => \N__26858\
        );

    \I__4142\ : InMux
    port map (
            O => \N__26858\,
            I => \N__26855\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__26855\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\
        );

    \I__4140\ : InMux
    port map (
            O => \N__26852\,
            I => \N__26848\
        );

    \I__4139\ : InMux
    port map (
            O => \N__26851\,
            I => \N__26845\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__26848\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__26845\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__4136\ : CascadeMux
    port map (
            O => \N__26840\,
            I => \N__26837\
        );

    \I__4135\ : InMux
    port map (
            O => \N__26837\,
            I => \N__26834\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__26834\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\
        );

    \I__4133\ : InMux
    port map (
            O => \N__26831\,
            I => \N__26827\
        );

    \I__4132\ : InMux
    port map (
            O => \N__26830\,
            I => \N__26824\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__26827\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__26824\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__4129\ : CascadeMux
    port map (
            O => \N__26819\,
            I => \N__26816\
        );

    \I__4128\ : InMux
    port map (
            O => \N__26816\,
            I => \N__26813\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__26813\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\
        );

    \I__4126\ : InMux
    port map (
            O => \N__26810\,
            I => \N__26806\
        );

    \I__4125\ : InMux
    port map (
            O => \N__26809\,
            I => \N__26803\
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__26806\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__26803\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__4122\ : CascadeMux
    port map (
            O => \N__26798\,
            I => \N__26795\
        );

    \I__4121\ : InMux
    port map (
            O => \N__26795\,
            I => \N__26792\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__26792\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\
        );

    \I__4119\ : CascadeMux
    port map (
            O => \N__26789\,
            I => \N__26786\
        );

    \I__4118\ : InMux
    port map (
            O => \N__26786\,
            I => \N__26783\
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__26783\,
            I => \N__26780\
        );

    \I__4116\ : Odrv12
    port map (
            O => \N__26780\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\
        );

    \I__4115\ : InMux
    port map (
            O => \N__26777\,
            I => \N__26773\
        );

    \I__4114\ : InMux
    port map (
            O => \N__26776\,
            I => \N__26770\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__26773\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__26770\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__4111\ : InMux
    port map (
            O => \N__26765\,
            I => \N__26762\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__26762\,
            I => \N__26759\
        );

    \I__4109\ : Odrv4
    port map (
            O => \N__26759\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\
        );

    \I__4108\ : InMux
    port map (
            O => \N__26756\,
            I => \N__26752\
        );

    \I__4107\ : InMux
    port map (
            O => \N__26755\,
            I => \N__26749\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__26752\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__26749\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__4104\ : CascadeMux
    port map (
            O => \N__26744\,
            I => \N__26741\
        );

    \I__4103\ : InMux
    port map (
            O => \N__26741\,
            I => \N__26738\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__26738\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\
        );

    \I__4101\ : InMux
    port map (
            O => \N__26735\,
            I => \N__26731\
        );

    \I__4100\ : InMux
    port map (
            O => \N__26734\,
            I => \N__26728\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__26731\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__26728\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14\
        );

    \I__4097\ : InMux
    port map (
            O => \N__26723\,
            I => \N__26719\
        );

    \I__4096\ : InMux
    port map (
            O => \N__26722\,
            I => \N__26714\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__26719\,
            I => \N__26711\
        );

    \I__4094\ : InMux
    port map (
            O => \N__26718\,
            I => \N__26706\
        );

    \I__4093\ : InMux
    port map (
            O => \N__26717\,
            I => \N__26706\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__26714\,
            I => \N__26703\
        );

    \I__4091\ : Odrv4
    port map (
            O => \N__26711\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__26706\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\
        );

    \I__4089\ : Odrv4
    port map (
            O => \N__26703\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\
        );

    \I__4088\ : InMux
    port map (
            O => \N__26696\,
            I => \N__26693\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__26693\,
            I => \N__26687\
        );

    \I__4086\ : InMux
    port map (
            O => \N__26692\,
            I => \N__26682\
        );

    \I__4085\ : InMux
    port map (
            O => \N__26691\,
            I => \N__26682\
        );

    \I__4084\ : InMux
    port map (
            O => \N__26690\,
            I => \N__26679\
        );

    \I__4083\ : Odrv4
    port map (
            O => \N__26687\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__4082\ : LocalMux
    port map (
            O => \N__26682\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__4081\ : LocalMux
    port map (
            O => \N__26679\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__4080\ : InMux
    port map (
            O => \N__26672\,
            I => \N__26668\
        );

    \I__4079\ : InMux
    port map (
            O => \N__26671\,
            I => \N__26665\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__26668\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__26665\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18\
        );

    \I__4076\ : InMux
    port map (
            O => \N__26660\,
            I => \N__26654\
        );

    \I__4075\ : InMux
    port map (
            O => \N__26659\,
            I => \N__26654\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__26654\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_24\
        );

    \I__4073\ : InMux
    port map (
            O => \N__26651\,
            I => \N__26644\
        );

    \I__4072\ : InMux
    port map (
            O => \N__26650\,
            I => \N__26644\
        );

    \I__4071\ : InMux
    port map (
            O => \N__26649\,
            I => \N__26641\
        );

    \I__4070\ : LocalMux
    port map (
            O => \N__26644\,
            I => \N__26638\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__26641\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__4068\ : Odrv4
    port map (
            O => \N__26638\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__4067\ : CascadeMux
    port map (
            O => \N__26633\,
            I => \N__26630\
        );

    \I__4066\ : InMux
    port map (
            O => \N__26630\,
            I => \N__26623\
        );

    \I__4065\ : InMux
    port map (
            O => \N__26629\,
            I => \N__26623\
        );

    \I__4064\ : InMux
    port map (
            O => \N__26628\,
            I => \N__26620\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__26623\,
            I => \N__26617\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__26620\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__4061\ : Odrv4
    port map (
            O => \N__26617\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__4060\ : CascadeMux
    port map (
            O => \N__26612\,
            I => \N__26609\
        );

    \I__4059\ : InMux
    port map (
            O => \N__26609\,
            I => \N__26603\
        );

    \I__4058\ : InMux
    port map (
            O => \N__26608\,
            I => \N__26603\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__26603\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\
        );

    \I__4056\ : CascadeMux
    port map (
            O => \N__26600\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18_cascade_\
        );

    \I__4055\ : InMux
    port map (
            O => \N__26597\,
            I => \N__26591\
        );

    \I__4054\ : InMux
    port map (
            O => \N__26596\,
            I => \N__26591\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__26591\,
            I => \N__26588\
        );

    \I__4052\ : Odrv4
    port map (
            O => \N__26588\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\
        );

    \I__4051\ : InMux
    port map (
            O => \N__26585\,
            I => \N__26579\
        );

    \I__4050\ : InMux
    port map (
            O => \N__26584\,
            I => \N__26579\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__26579\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\
        );

    \I__4048\ : CascadeMux
    port map (
            O => \N__26576\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14_cascade_\
        );

    \I__4047\ : CascadeMux
    port map (
            O => \N__26573\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17_cascade_\
        );

    \I__4046\ : InMux
    port map (
            O => \N__26570\,
            I => \N__26567\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__26567\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3\
        );

    \I__4044\ : InMux
    port map (
            O => \N__26564\,
            I => \N__26561\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__26561\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23\
        );

    \I__4042\ : CascadeMux
    port map (
            O => \N__26558\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21_cascade_\
        );

    \I__4041\ : InMux
    port map (
            O => \N__26555\,
            I => \N__26552\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__26552\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\
        );

    \I__4039\ : InMux
    port map (
            O => \N__26549\,
            I => \N__26546\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__26546\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\
        );

    \I__4037\ : InMux
    port map (
            O => \N__26543\,
            I => \N__26540\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__26540\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\
        );

    \I__4035\ : InMux
    port map (
            O => \N__26537\,
            I => \N__26534\
        );

    \I__4034\ : LocalMux
    port map (
            O => \N__26534\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20\
        );

    \I__4033\ : CascadeMux
    port map (
            O => \N__26531\,
            I => \elapsed_time_ns_1_RNIV9PBB_0_21_cascade_\
        );

    \I__4032\ : InMux
    port map (
            O => \N__26528\,
            I => \N__26522\
        );

    \I__4031\ : InMux
    port map (
            O => \N__26527\,
            I => \N__26522\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__26522\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_23\
        );

    \I__4029\ : CascadeMux
    port map (
            O => \N__26519\,
            I => \N__26515\
        );

    \I__4028\ : InMux
    port map (
            O => \N__26518\,
            I => \N__26510\
        );

    \I__4027\ : InMux
    port map (
            O => \N__26515\,
            I => \N__26510\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__26510\,
            I => \N__26507\
        );

    \I__4025\ : Span4Mux_h
    port map (
            O => \N__26507\,
            I => \N__26503\
        );

    \I__4024\ : InMux
    port map (
            O => \N__26506\,
            I => \N__26500\
        );

    \I__4023\ : Span4Mux_v
    port map (
            O => \N__26503\,
            I => \N__26497\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__26500\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__4021\ : Odrv4
    port map (
            O => \N__26497\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__4020\ : InMux
    port map (
            O => \N__26492\,
            I => \N__26486\
        );

    \I__4019\ : InMux
    port map (
            O => \N__26491\,
            I => \N__26486\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__26486\,
            I => \N__26482\
        );

    \I__4017\ : InMux
    port map (
            O => \N__26485\,
            I => \N__26479\
        );

    \I__4016\ : Span4Mux_v
    port map (
            O => \N__26482\,
            I => \N__26476\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__26479\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__4014\ : Odrv4
    port map (
            O => \N__26476\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__4013\ : CascadeMux
    port map (
            O => \N__26471\,
            I => \N__26467\
        );

    \I__4012\ : InMux
    port map (
            O => \N__26470\,
            I => \N__26462\
        );

    \I__4011\ : InMux
    port map (
            O => \N__26467\,
            I => \N__26462\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__26462\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_22\
        );

    \I__4009\ : InMux
    port map (
            O => \N__26459\,
            I => \N__26456\
        );

    \I__4008\ : LocalMux
    port map (
            O => \N__26456\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15\
        );

    \I__4007\ : CascadeMux
    port map (
            O => \N__26453\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22_cascade_\
        );

    \I__4006\ : CascadeMux
    port map (
            O => \N__26450\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\
        );

    \I__4005\ : InMux
    port map (
            O => \N__26447\,
            I => \N__26443\
        );

    \I__4004\ : InMux
    port map (
            O => \N__26446\,
            I => \N__26440\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__26443\,
            I => \phase_controller_inst2.stoper_tr.runningZ0\
        );

    \I__4002\ : LocalMux
    port map (
            O => \N__26440\,
            I => \phase_controller_inst2.stoper_tr.runningZ0\
        );

    \I__4001\ : InMux
    port map (
            O => \N__26435\,
            I => \N__26432\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__26432\,
            I => \phase_controller_inst2.start_timer_hc_0_sqmuxa\
        );

    \I__3999\ : InMux
    port map (
            O => \N__26429\,
            I => \N__26426\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__26426\,
            I => \N__26422\
        );

    \I__3997\ : InMux
    port map (
            O => \N__26425\,
            I => \N__26419\
        );

    \I__3996\ : Span4Mux_v
    port map (
            O => \N__26422\,
            I => \N__26416\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__26419\,
            I => \N__26413\
        );

    \I__3994\ : Odrv4
    port map (
            O => \N__26416\,
            I => \phase_controller_inst2.state_RNIG7JFZ0Z_2\
        );

    \I__3993\ : Odrv12
    port map (
            O => \N__26413\,
            I => \phase_controller_inst2.state_RNIG7JFZ0Z_2\
        );

    \I__3992\ : InMux
    port map (
            O => \N__26408\,
            I => \N__26402\
        );

    \I__3991\ : InMux
    port map (
            O => \N__26407\,
            I => \N__26399\
        );

    \I__3990\ : InMux
    port map (
            O => \N__26406\,
            I => \N__26396\
        );

    \I__3989\ : InMux
    port map (
            O => \N__26405\,
            I => \N__26393\
        );

    \I__3988\ : LocalMux
    port map (
            O => \N__26402\,
            I => \N__26390\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__26399\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__26396\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__26393\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__3984\ : Odrv12
    port map (
            O => \N__26390\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__3983\ : CEMux
    port map (
            O => \N__26381\,
            I => \N__26376\
        );

    \I__3982\ : CEMux
    port map (
            O => \N__26380\,
            I => \N__26373\
        );

    \I__3981\ : CEMux
    port map (
            O => \N__26379\,
            I => \N__26368\
        );

    \I__3980\ : LocalMux
    port map (
            O => \N__26376\,
            I => \N__26365\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__26373\,
            I => \N__26362\
        );

    \I__3978\ : CEMux
    port map (
            O => \N__26372\,
            I => \N__26359\
        );

    \I__3977\ : CEMux
    port map (
            O => \N__26371\,
            I => \N__26356\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__26368\,
            I => \N__26353\
        );

    \I__3975\ : Span4Mux_v
    port map (
            O => \N__26365\,
            I => \N__26346\
        );

    \I__3974\ : Span4Mux_v
    port map (
            O => \N__26362\,
            I => \N__26346\
        );

    \I__3973\ : LocalMux
    port map (
            O => \N__26359\,
            I => \N__26346\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__26356\,
            I => \N__26343\
        );

    \I__3971\ : Span4Mux_v
    port map (
            O => \N__26353\,
            I => \N__26340\
        );

    \I__3970\ : Span4Mux_v
    port map (
            O => \N__26346\,
            I => \N__26337\
        );

    \I__3969\ : Odrv12
    port map (
            O => \N__26343\,
            I => \delay_measurement_inst.delay_tr_timer.N_200_i\
        );

    \I__3968\ : Odrv4
    port map (
            O => \N__26340\,
            I => \delay_measurement_inst.delay_tr_timer.N_200_i\
        );

    \I__3967\ : Odrv4
    port map (
            O => \N__26337\,
            I => \delay_measurement_inst.delay_tr_timer.N_200_i\
        );

    \I__3966\ : InMux
    port map (
            O => \N__26330\,
            I => \N__26324\
        );

    \I__3965\ : InMux
    port map (
            O => \N__26329\,
            I => \N__26319\
        );

    \I__3964\ : InMux
    port map (
            O => \N__26328\,
            I => \N__26319\
        );

    \I__3963\ : InMux
    port map (
            O => \N__26327\,
            I => \N__26316\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__26324\,
            I => \N__26313\
        );

    \I__3961\ : LocalMux
    port map (
            O => \N__26319\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__26316\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__3959\ : Odrv4
    port map (
            O => \N__26313\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__3958\ : CascadeMux
    port map (
            O => \N__26306\,
            I => \N__26303\
        );

    \I__3957\ : InMux
    port map (
            O => \N__26303\,
            I => \N__26299\
        );

    \I__3956\ : InMux
    port map (
            O => \N__26302\,
            I => \N__26295\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__26299\,
            I => \N__26292\
        );

    \I__3954\ : InMux
    port map (
            O => \N__26298\,
            I => \N__26289\
        );

    \I__3953\ : LocalMux
    port map (
            O => \N__26295\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__3952\ : Odrv4
    port map (
            O => \N__26292\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__26289\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__3950\ : ClkMux
    port map (
            O => \N__26282\,
            I => \N__26279\
        );

    \I__3949\ : GlobalMux
    port map (
            O => \N__26279\,
            I => \N__26276\
        );

    \I__3948\ : gio2CtrlBuf
    port map (
            O => \N__26276\,
            I => delay_tr_input_c_g
        );

    \I__3947\ : InMux
    port map (
            O => \N__26273\,
            I => \N__26270\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__26270\,
            I => \N__26265\
        );

    \I__3945\ : CascadeMux
    port map (
            O => \N__26269\,
            I => \N__26261\
        );

    \I__3944\ : CascadeMux
    port map (
            O => \N__26268\,
            I => \N__26258\
        );

    \I__3943\ : Span12Mux_s5_v
    port map (
            O => \N__26265\,
            I => \N__26255\
        );

    \I__3942\ : InMux
    port map (
            O => \N__26264\,
            I => \N__26252\
        );

    \I__3941\ : InMux
    port map (
            O => \N__26261\,
            I => \N__26247\
        );

    \I__3940\ : InMux
    port map (
            O => \N__26258\,
            I => \N__26247\
        );

    \I__3939\ : Span12Mux_v
    port map (
            O => \N__26255\,
            I => \N__26244\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__26252\,
            I => \N__26241\
        );

    \I__3937\ : LocalMux
    port map (
            O => \N__26247\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__3936\ : Odrv12
    port map (
            O => \N__26244\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__3935\ : Odrv4
    port map (
            O => \N__26241\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__3934\ : IoInMux
    port map (
            O => \N__26234\,
            I => \N__26231\
        );

    \I__3933\ : LocalMux
    port map (
            O => \N__26231\,
            I => \N__26228\
        );

    \I__3932\ : Odrv4
    port map (
            O => \N__26228\,
            I => s3_phy_c
        );

    \I__3931\ : InMux
    port map (
            O => \N__26225\,
            I => \N__26222\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__26222\,
            I => \N__26219\
        );

    \I__3929\ : Span4Mux_v
    port map (
            O => \N__26219\,
            I => \N__26214\
        );

    \I__3928\ : InMux
    port map (
            O => \N__26218\,
            I => \N__26211\
        );

    \I__3927\ : CascadeMux
    port map (
            O => \N__26217\,
            I => \N__26208\
        );

    \I__3926\ : Span4Mux_v
    port map (
            O => \N__26214\,
            I => \N__26204\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__26211\,
            I => \N__26201\
        );

    \I__3924\ : InMux
    port map (
            O => \N__26208\,
            I => \N__26198\
        );

    \I__3923\ : InMux
    port map (
            O => \N__26207\,
            I => \N__26195\
        );

    \I__3922\ : Span4Mux_v
    port map (
            O => \N__26204\,
            I => \N__26192\
        );

    \I__3921\ : Span4Mux_h
    port map (
            O => \N__26201\,
            I => \N__26189\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__26198\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__26195\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__3918\ : Odrv4
    port map (
            O => \N__26192\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__3917\ : Odrv4
    port map (
            O => \N__26189\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__3916\ : IoInMux
    port map (
            O => \N__26180\,
            I => \N__26177\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__26177\,
            I => \N__26174\
        );

    \I__3914\ : Odrv4
    port map (
            O => \N__26174\,
            I => s4_phy_c
        );

    \I__3913\ : IoInMux
    port map (
            O => \N__26171\,
            I => \N__26168\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__26168\,
            I => \GB_BUFFER_clock_output_0_THRU_CO\
        );

    \I__3911\ : InMux
    port map (
            O => \N__26165\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\
        );

    \I__3910\ : InMux
    port map (
            O => \N__26162\,
            I => \bfn_8_14_0_\
        );

    \I__3909\ : CascadeMux
    port map (
            O => \N__26159\,
            I => \N__26154\
        );

    \I__3908\ : InMux
    port map (
            O => \N__26158\,
            I => \N__26151\
        );

    \I__3907\ : InMux
    port map (
            O => \N__26157\,
            I => \N__26146\
        );

    \I__3906\ : InMux
    port map (
            O => \N__26154\,
            I => \N__26146\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__26151\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__26146\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__3903\ : InMux
    port map (
            O => \N__26141\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\
        );

    \I__3902\ : InMux
    port map (
            O => \N__26138\,
            I => \N__26133\
        );

    \I__3901\ : InMux
    port map (
            O => \N__26137\,
            I => \N__26128\
        );

    \I__3900\ : InMux
    port map (
            O => \N__26136\,
            I => \N__26128\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__26133\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__26128\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__3897\ : InMux
    port map (
            O => \N__26123\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\
        );

    \I__3896\ : InMux
    port map (
            O => \N__26120\,
            I => \N__26115\
        );

    \I__3895\ : InMux
    port map (
            O => \N__26119\,
            I => \N__26110\
        );

    \I__3894\ : InMux
    port map (
            O => \N__26118\,
            I => \N__26110\
        );

    \I__3893\ : LocalMux
    port map (
            O => \N__26115\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__26110\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__3891\ : InMux
    port map (
            O => \N__26105\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\
        );

    \I__3890\ : CascadeMux
    port map (
            O => \N__26102\,
            I => \N__26097\
        );

    \I__3889\ : InMux
    port map (
            O => \N__26101\,
            I => \N__26094\
        );

    \I__3888\ : InMux
    port map (
            O => \N__26100\,
            I => \N__26089\
        );

    \I__3887\ : InMux
    port map (
            O => \N__26097\,
            I => \N__26089\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__26094\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__26089\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__3884\ : InMux
    port map (
            O => \N__26084\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\
        );

    \I__3883\ : InMux
    port map (
            O => \N__26081\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\
        );

    \I__3882\ : InMux
    port map (
            O => \N__26078\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\
        );

    \I__3881\ : InMux
    port map (
            O => \N__26075\,
            I => \N__26070\
        );

    \I__3880\ : InMux
    port map (
            O => \N__26074\,
            I => \N__26067\
        );

    \I__3879\ : InMux
    port map (
            O => \N__26073\,
            I => \N__26064\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__26070\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__26067\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__26064\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__3875\ : InMux
    port map (
            O => \N__26057\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\
        );

    \I__3874\ : InMux
    port map (
            O => \N__26054\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\
        );

    \I__3873\ : InMux
    port map (
            O => \N__26051\,
            I => \bfn_8_13_0_\
        );

    \I__3872\ : InMux
    port map (
            O => \N__26048\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\
        );

    \I__3871\ : InMux
    port map (
            O => \N__26045\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\
        );

    \I__3870\ : InMux
    port map (
            O => \N__26042\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\
        );

    \I__3869\ : InMux
    port map (
            O => \N__26039\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__3868\ : InMux
    port map (
            O => \N__26036\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\
        );

    \I__3867\ : InMux
    port map (
            O => \N__26033\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\
        );

    \I__3866\ : InMux
    port map (
            O => \N__26030\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\
        );

    \I__3865\ : InMux
    port map (
            O => \N__26027\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\
        );

    \I__3864\ : InMux
    port map (
            O => \N__26024\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\
        );

    \I__3863\ : InMux
    port map (
            O => \N__26021\,
            I => \bfn_8_12_0_\
        );

    \I__3862\ : InMux
    port map (
            O => \N__26018\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\
        );

    \I__3861\ : InMux
    port map (
            O => \N__26015\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\
        );

    \I__3860\ : InMux
    port map (
            O => \N__26012\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\
        );

    \I__3859\ : InMux
    port map (
            O => \N__26009\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\
        );

    \I__3858\ : InMux
    port map (
            O => \N__26006\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\
        );

    \I__3857\ : InMux
    port map (
            O => \N__26003\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__3856\ : InMux
    port map (
            O => \N__26000\,
            I => \N__25996\
        );

    \I__3855\ : InMux
    port map (
            O => \N__25999\,
            I => \N__25993\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__25996\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__25993\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__3852\ : CascadeMux
    port map (
            O => \N__25988\,
            I => \N__25985\
        );

    \I__3851\ : InMux
    port map (
            O => \N__25985\,
            I => \N__25980\
        );

    \I__3850\ : InMux
    port map (
            O => \N__25984\,
            I => \N__25977\
        );

    \I__3849\ : InMux
    port map (
            O => \N__25983\,
            I => \N__25974\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__25980\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__25977\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__25974\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__3845\ : InMux
    port map (
            O => \N__25967\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__3844\ : InMux
    port map (
            O => \N__25964\,
            I => \N__25960\
        );

    \I__3843\ : InMux
    port map (
            O => \N__25963\,
            I => \N__25957\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__25960\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__25957\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__3840\ : CascadeMux
    port map (
            O => \N__25952\,
            I => \N__25949\
        );

    \I__3839\ : InMux
    port map (
            O => \N__25949\,
            I => \N__25944\
        );

    \I__3838\ : InMux
    port map (
            O => \N__25948\,
            I => \N__25941\
        );

    \I__3837\ : InMux
    port map (
            O => \N__25947\,
            I => \N__25938\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__25944\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__25941\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__25938\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__3833\ : InMux
    port map (
            O => \N__25931\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__3832\ : InMux
    port map (
            O => \N__25928\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__3831\ : CascadeMux
    port map (
            O => \N__25925\,
            I => \N__25922\
        );

    \I__3830\ : InMux
    port map (
            O => \N__25922\,
            I => \N__25919\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__25919\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\
        );

    \I__3828\ : InMux
    port map (
            O => \N__25916\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\
        );

    \I__3827\ : CascadeMux
    port map (
            O => \N__25913\,
            I => \N__25910\
        );

    \I__3826\ : InMux
    port map (
            O => \N__25910\,
            I => \N__25907\
        );

    \I__3825\ : LocalMux
    port map (
            O => \N__25907\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1Z0Z_30\
        );

    \I__3824\ : InMux
    port map (
            O => \N__25904\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\
        );

    \I__3823\ : InMux
    port map (
            O => \N__25901\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\
        );

    \I__3822\ : InMux
    port map (
            O => \N__25898\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\
        );

    \I__3821\ : CascadeMux
    port map (
            O => \N__25895\,
            I => \N__25892\
        );

    \I__3820\ : InMux
    port map (
            O => \N__25892\,
            I => \N__25887\
        );

    \I__3819\ : InMux
    port map (
            O => \N__25891\,
            I => \N__25884\
        );

    \I__3818\ : InMux
    port map (
            O => \N__25890\,
            I => \N__25881\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__25887\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__25884\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__3815\ : LocalMux
    port map (
            O => \N__25881\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__3814\ : InMux
    port map (
            O => \N__25874\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__3813\ : CascadeMux
    port map (
            O => \N__25871\,
            I => \N__25868\
        );

    \I__3812\ : InMux
    port map (
            O => \N__25868\,
            I => \N__25863\
        );

    \I__3811\ : InMux
    port map (
            O => \N__25867\,
            I => \N__25860\
        );

    \I__3810\ : InMux
    port map (
            O => \N__25866\,
            I => \N__25857\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__25863\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__25860\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__25857\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__3806\ : InMux
    port map (
            O => \N__25850\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__3805\ : CascadeMux
    port map (
            O => \N__25847\,
            I => \N__25844\
        );

    \I__3804\ : InMux
    port map (
            O => \N__25844\,
            I => \N__25839\
        );

    \I__3803\ : InMux
    port map (
            O => \N__25843\,
            I => \N__25836\
        );

    \I__3802\ : InMux
    port map (
            O => \N__25842\,
            I => \N__25833\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__25839\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__25836\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__25833\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__3798\ : InMux
    port map (
            O => \N__25826\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__3797\ : CascadeMux
    port map (
            O => \N__25823\,
            I => \N__25820\
        );

    \I__3796\ : InMux
    port map (
            O => \N__25820\,
            I => \N__25815\
        );

    \I__3795\ : InMux
    port map (
            O => \N__25819\,
            I => \N__25812\
        );

    \I__3794\ : InMux
    port map (
            O => \N__25818\,
            I => \N__25809\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__25815\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__25812\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__25809\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__3790\ : InMux
    port map (
            O => \N__25802\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__3789\ : CascadeMux
    port map (
            O => \N__25799\,
            I => \N__25796\
        );

    \I__3788\ : InMux
    port map (
            O => \N__25796\,
            I => \N__25791\
        );

    \I__3787\ : InMux
    port map (
            O => \N__25795\,
            I => \N__25788\
        );

    \I__3786\ : InMux
    port map (
            O => \N__25794\,
            I => \N__25785\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__25791\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__25788\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__25785\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__3782\ : InMux
    port map (
            O => \N__25778\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__3781\ : CascadeMux
    port map (
            O => \N__25775\,
            I => \N__25772\
        );

    \I__3780\ : InMux
    port map (
            O => \N__25772\,
            I => \N__25767\
        );

    \I__3779\ : InMux
    port map (
            O => \N__25771\,
            I => \N__25764\
        );

    \I__3778\ : InMux
    port map (
            O => \N__25770\,
            I => \N__25761\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__25767\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__25764\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__3775\ : LocalMux
    port map (
            O => \N__25761\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__3774\ : InMux
    port map (
            O => \N__25754\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__3773\ : CascadeMux
    port map (
            O => \N__25751\,
            I => \N__25748\
        );

    \I__3772\ : InMux
    port map (
            O => \N__25748\,
            I => \N__25743\
        );

    \I__3771\ : InMux
    port map (
            O => \N__25747\,
            I => \N__25740\
        );

    \I__3770\ : InMux
    port map (
            O => \N__25746\,
            I => \N__25737\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__25743\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__25740\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__25737\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__3766\ : InMux
    port map (
            O => \N__25730\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__3765\ : CascadeMux
    port map (
            O => \N__25727\,
            I => \N__25724\
        );

    \I__3764\ : InMux
    port map (
            O => \N__25724\,
            I => \N__25719\
        );

    \I__3763\ : InMux
    port map (
            O => \N__25723\,
            I => \N__25716\
        );

    \I__3762\ : InMux
    port map (
            O => \N__25722\,
            I => \N__25713\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__25719\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__25716\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__25713\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__3758\ : InMux
    port map (
            O => \N__25706\,
            I => \bfn_8_10_0_\
        );

    \I__3757\ : CascadeMux
    port map (
            O => \N__25703\,
            I => \N__25700\
        );

    \I__3756\ : InMux
    port map (
            O => \N__25700\,
            I => \N__25695\
        );

    \I__3755\ : InMux
    port map (
            O => \N__25699\,
            I => \N__25692\
        );

    \I__3754\ : InMux
    port map (
            O => \N__25698\,
            I => \N__25689\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__25695\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__25692\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__25689\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__3750\ : CascadeMux
    port map (
            O => \N__25682\,
            I => \N__25679\
        );

    \I__3749\ : InMux
    port map (
            O => \N__25679\,
            I => \N__25674\
        );

    \I__3748\ : InMux
    port map (
            O => \N__25678\,
            I => \N__25671\
        );

    \I__3747\ : InMux
    port map (
            O => \N__25677\,
            I => \N__25668\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__25674\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__3745\ : LocalMux
    port map (
            O => \N__25671\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__25668\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__3743\ : InMux
    port map (
            O => \N__25661\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__3742\ : CascadeMux
    port map (
            O => \N__25658\,
            I => \N__25655\
        );

    \I__3741\ : InMux
    port map (
            O => \N__25655\,
            I => \N__25650\
        );

    \I__3740\ : InMux
    port map (
            O => \N__25654\,
            I => \N__25647\
        );

    \I__3739\ : InMux
    port map (
            O => \N__25653\,
            I => \N__25644\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__25650\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__25647\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__25644\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__3735\ : InMux
    port map (
            O => \N__25637\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__3734\ : CascadeMux
    port map (
            O => \N__25634\,
            I => \N__25631\
        );

    \I__3733\ : InMux
    port map (
            O => \N__25631\,
            I => \N__25626\
        );

    \I__3732\ : InMux
    port map (
            O => \N__25630\,
            I => \N__25623\
        );

    \I__3731\ : InMux
    port map (
            O => \N__25629\,
            I => \N__25620\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__25626\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__25623\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__25620\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__3727\ : InMux
    port map (
            O => \N__25613\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__3726\ : CascadeMux
    port map (
            O => \N__25610\,
            I => \N__25607\
        );

    \I__3725\ : InMux
    port map (
            O => \N__25607\,
            I => \N__25602\
        );

    \I__3724\ : InMux
    port map (
            O => \N__25606\,
            I => \N__25599\
        );

    \I__3723\ : InMux
    port map (
            O => \N__25605\,
            I => \N__25596\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__25602\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__25599\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__25596\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__3719\ : InMux
    port map (
            O => \N__25589\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__3718\ : CascadeMux
    port map (
            O => \N__25586\,
            I => \N__25583\
        );

    \I__3717\ : InMux
    port map (
            O => \N__25583\,
            I => \N__25578\
        );

    \I__3716\ : InMux
    port map (
            O => \N__25582\,
            I => \N__25575\
        );

    \I__3715\ : InMux
    port map (
            O => \N__25581\,
            I => \N__25572\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__25578\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__25575\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__25572\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__3711\ : InMux
    port map (
            O => \N__25565\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__3710\ : CascadeMux
    port map (
            O => \N__25562\,
            I => \N__25559\
        );

    \I__3709\ : InMux
    port map (
            O => \N__25559\,
            I => \N__25554\
        );

    \I__3708\ : InMux
    port map (
            O => \N__25558\,
            I => \N__25551\
        );

    \I__3707\ : InMux
    port map (
            O => \N__25557\,
            I => \N__25548\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__25554\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__3705\ : LocalMux
    port map (
            O => \N__25551\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__25548\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__3703\ : InMux
    port map (
            O => \N__25541\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__3702\ : CascadeMux
    port map (
            O => \N__25538\,
            I => \N__25535\
        );

    \I__3701\ : InMux
    port map (
            O => \N__25535\,
            I => \N__25530\
        );

    \I__3700\ : InMux
    port map (
            O => \N__25534\,
            I => \N__25527\
        );

    \I__3699\ : InMux
    port map (
            O => \N__25533\,
            I => \N__25524\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__25530\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__25527\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__25524\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__3695\ : InMux
    port map (
            O => \N__25517\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__3694\ : CascadeMux
    port map (
            O => \N__25514\,
            I => \N__25511\
        );

    \I__3693\ : InMux
    port map (
            O => \N__25511\,
            I => \N__25506\
        );

    \I__3692\ : InMux
    port map (
            O => \N__25510\,
            I => \N__25503\
        );

    \I__3691\ : InMux
    port map (
            O => \N__25509\,
            I => \N__25500\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__25506\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__25503\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__25500\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__3687\ : InMux
    port map (
            O => \N__25493\,
            I => \bfn_8_9_0_\
        );

    \I__3686\ : CascadeMux
    port map (
            O => \N__25490\,
            I => \N__25486\
        );

    \I__3685\ : InMux
    port map (
            O => \N__25489\,
            I => \N__25482\
        );

    \I__3684\ : InMux
    port map (
            O => \N__25486\,
            I => \N__25479\
        );

    \I__3683\ : InMux
    port map (
            O => \N__25485\,
            I => \N__25476\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__25482\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__25479\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__25476\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__3679\ : CascadeMux
    port map (
            O => \N__25469\,
            I => \N__25465\
        );

    \I__3678\ : InMux
    port map (
            O => \N__25468\,
            I => \N__25461\
        );

    \I__3677\ : InMux
    port map (
            O => \N__25465\,
            I => \N__25458\
        );

    \I__3676\ : InMux
    port map (
            O => \N__25464\,
            I => \N__25455\
        );

    \I__3675\ : LocalMux
    port map (
            O => \N__25461\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__25458\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__25455\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__3672\ : InMux
    port map (
            O => \N__25448\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__3671\ : CascadeMux
    port map (
            O => \N__25445\,
            I => \N__25442\
        );

    \I__3670\ : InMux
    port map (
            O => \N__25442\,
            I => \N__25437\
        );

    \I__3669\ : InMux
    port map (
            O => \N__25441\,
            I => \N__25434\
        );

    \I__3668\ : InMux
    port map (
            O => \N__25440\,
            I => \N__25431\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__25437\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__3666\ : LocalMux
    port map (
            O => \N__25434\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__25431\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__3664\ : InMux
    port map (
            O => \N__25424\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__3663\ : CascadeMux
    port map (
            O => \N__25421\,
            I => \N__25418\
        );

    \I__3662\ : InMux
    port map (
            O => \N__25418\,
            I => \N__25413\
        );

    \I__3661\ : InMux
    port map (
            O => \N__25417\,
            I => \N__25410\
        );

    \I__3660\ : InMux
    port map (
            O => \N__25416\,
            I => \N__25407\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__25413\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__25410\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__25407\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__3656\ : InMux
    port map (
            O => \N__25400\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__3655\ : CascadeMux
    port map (
            O => \N__25397\,
            I => \N__25394\
        );

    \I__3654\ : InMux
    port map (
            O => \N__25394\,
            I => \N__25389\
        );

    \I__3653\ : InMux
    port map (
            O => \N__25393\,
            I => \N__25386\
        );

    \I__3652\ : InMux
    port map (
            O => \N__25392\,
            I => \N__25383\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__25389\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__25386\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__25383\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__3648\ : InMux
    port map (
            O => \N__25376\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__3647\ : CascadeMux
    port map (
            O => \N__25373\,
            I => \N__25370\
        );

    \I__3646\ : InMux
    port map (
            O => \N__25370\,
            I => \N__25365\
        );

    \I__3645\ : InMux
    port map (
            O => \N__25369\,
            I => \N__25362\
        );

    \I__3644\ : InMux
    port map (
            O => \N__25368\,
            I => \N__25359\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__25365\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__25362\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__25359\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__3640\ : InMux
    port map (
            O => \N__25352\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__3639\ : CascadeMux
    port map (
            O => \N__25349\,
            I => \N__25346\
        );

    \I__3638\ : InMux
    port map (
            O => \N__25346\,
            I => \N__25341\
        );

    \I__3637\ : InMux
    port map (
            O => \N__25345\,
            I => \N__25338\
        );

    \I__3636\ : InMux
    port map (
            O => \N__25344\,
            I => \N__25335\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__25341\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__25338\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__25335\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__3632\ : InMux
    port map (
            O => \N__25328\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__3631\ : CascadeMux
    port map (
            O => \N__25325\,
            I => \N__25322\
        );

    \I__3630\ : InMux
    port map (
            O => \N__25322\,
            I => \N__25317\
        );

    \I__3629\ : InMux
    port map (
            O => \N__25321\,
            I => \N__25314\
        );

    \I__3628\ : InMux
    port map (
            O => \N__25320\,
            I => \N__25311\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__25317\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__25314\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__25311\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__3624\ : InMux
    port map (
            O => \N__25304\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__3623\ : CascadeMux
    port map (
            O => \N__25301\,
            I => \N__25298\
        );

    \I__3622\ : InMux
    port map (
            O => \N__25298\,
            I => \N__25293\
        );

    \I__3621\ : InMux
    port map (
            O => \N__25297\,
            I => \N__25290\
        );

    \I__3620\ : InMux
    port map (
            O => \N__25296\,
            I => \N__25287\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__25293\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__25290\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__25287\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__3616\ : InMux
    port map (
            O => \N__25280\,
            I => \bfn_8_8_0_\
        );

    \I__3615\ : InMux
    port map (
            O => \N__25277\,
            I => \N__25272\
        );

    \I__3614\ : InMux
    port map (
            O => \N__25276\,
            I => \N__25269\
        );

    \I__3613\ : InMux
    port map (
            O => \N__25275\,
            I => \N__25266\
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__25272\,
            I => \N__25259\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__25269\,
            I => \N__25259\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__25266\,
            I => \N__25259\
        );

    \I__3609\ : Span12Mux_v
    port map (
            O => \N__25259\,
            I => \N__25256\
        );

    \I__3608\ : Odrv12
    port map (
            O => \N__25256\,
            I => il_min_comp2_c
        );

    \I__3607\ : InMux
    port map (
            O => \N__25253\,
            I => \N__25249\
        );

    \I__3606\ : InMux
    port map (
            O => \N__25252\,
            I => \N__25246\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__25249\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__25246\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__3603\ : CascadeMux
    port map (
            O => \N__25241\,
            I => \N__25238\
        );

    \I__3602\ : InMux
    port map (
            O => \N__25238\,
            I => \N__25232\
        );

    \I__3601\ : InMux
    port map (
            O => \N__25237\,
            I => \N__25232\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__25232\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_27\
        );

    \I__3599\ : CascadeMux
    port map (
            O => \N__25229\,
            I => \N__25225\
        );

    \I__3598\ : InMux
    port map (
            O => \N__25228\,
            I => \N__25220\
        );

    \I__3597\ : InMux
    port map (
            O => \N__25225\,
            I => \N__25220\
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__25220\,
            I => \N__25217\
        );

    \I__3595\ : Span4Mux_v
    port map (
            O => \N__25217\,
            I => \N__25214\
        );

    \I__3594\ : Span4Mux_v
    port map (
            O => \N__25214\,
            I => \N__25211\
        );

    \I__3593\ : Odrv4
    port map (
            O => \N__25211\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\
        );

    \I__3592\ : InMux
    port map (
            O => \N__25208\,
            I => \N__25202\
        );

    \I__3591\ : InMux
    port map (
            O => \N__25207\,
            I => \N__25202\
        );

    \I__3590\ : LocalMux
    port map (
            O => \N__25202\,
            I => \N__25199\
        );

    \I__3589\ : Span4Mux_h
    port map (
            O => \N__25199\,
            I => \N__25196\
        );

    \I__3588\ : Odrv4
    port map (
            O => \N__25196\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_28\
        );

    \I__3587\ : InMux
    port map (
            O => \N__25193\,
            I => \N__25190\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__25190\,
            I => \N__25187\
        );

    \I__3585\ : Span4Mux_h
    port map (
            O => \N__25187\,
            I => \N__25182\
        );

    \I__3584\ : InMux
    port map (
            O => \N__25186\,
            I => \N__25177\
        );

    \I__3583\ : InMux
    port map (
            O => \N__25185\,
            I => \N__25177\
        );

    \I__3582\ : Span4Mux_v
    port map (
            O => \N__25182\,
            I => \N__25174\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__25177\,
            I => \N__25171\
        );

    \I__3580\ : Sp12to4
    port map (
            O => \N__25174\,
            I => \N__25166\
        );

    \I__3579\ : Span12Mux_h
    port map (
            O => \N__25171\,
            I => \N__25166\
        );

    \I__3578\ : Span12Mux_v
    port map (
            O => \N__25166\,
            I => \N__25163\
        );

    \I__3577\ : Odrv12
    port map (
            O => \N__25163\,
            I => il_max_comp2_c
        );

    \I__3576\ : CEMux
    port map (
            O => \N__25160\,
            I => \N__25157\
        );

    \I__3575\ : LocalMux
    port map (
            O => \N__25157\,
            I => \N__25153\
        );

    \I__3574\ : CEMux
    port map (
            O => \N__25156\,
            I => \N__25150\
        );

    \I__3573\ : Span4Mux_h
    port map (
            O => \N__25153\,
            I => \N__25143\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__25150\,
            I => \N__25143\
        );

    \I__3571\ : CEMux
    port map (
            O => \N__25149\,
            I => \N__25140\
        );

    \I__3570\ : CEMux
    port map (
            O => \N__25148\,
            I => \N__25137\
        );

    \I__3569\ : Span4Mux_v
    port map (
            O => \N__25143\,
            I => \N__25134\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__25140\,
            I => \N__25129\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__25137\,
            I => \N__25129\
        );

    \I__3566\ : Span4Mux_h
    port map (
            O => \N__25134\,
            I => \N__25124\
        );

    \I__3565\ : Span4Mux_v
    port map (
            O => \N__25129\,
            I => \N__25124\
        );

    \I__3564\ : Odrv4
    port map (
            O => \N__25124\,
            I => \delay_measurement_inst.delay_tr_timer.N_201_i\
        );

    \I__3563\ : InMux
    port map (
            O => \N__25121\,
            I => \N__25115\
        );

    \I__3562\ : InMux
    port map (
            O => \N__25120\,
            I => \N__25115\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__25115\,
            I => \N__25112\
        );

    \I__3560\ : Odrv4
    port map (
            O => \N__25112\,
            I => \phase_controller_inst2.state_RNI9M3OZ0Z_0\
        );

    \I__3559\ : InMux
    port map (
            O => \N__25109\,
            I => \N__25103\
        );

    \I__3558\ : InMux
    port map (
            O => \N__25108\,
            I => \N__25103\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__25103\,
            I => \N__25092\
        );

    \I__3556\ : InMux
    port map (
            O => \N__25102\,
            I => \N__25083\
        );

    \I__3555\ : InMux
    port map (
            O => \N__25101\,
            I => \N__25083\
        );

    \I__3554\ : InMux
    port map (
            O => \N__25100\,
            I => \N__25083\
        );

    \I__3553\ : InMux
    port map (
            O => \N__25099\,
            I => \N__25083\
        );

    \I__3552\ : InMux
    port map (
            O => \N__25098\,
            I => \N__25054\
        );

    \I__3551\ : InMux
    port map (
            O => \N__25097\,
            I => \N__25054\
        );

    \I__3550\ : InMux
    port map (
            O => \N__25096\,
            I => \N__25054\
        );

    \I__3549\ : InMux
    port map (
            O => \N__25095\,
            I => \N__25054\
        );

    \I__3548\ : Span4Mux_v
    port map (
            O => \N__25092\,
            I => \N__25049\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__25083\,
            I => \N__25049\
        );

    \I__3546\ : InMux
    port map (
            O => \N__25082\,
            I => \N__25040\
        );

    \I__3545\ : InMux
    port map (
            O => \N__25081\,
            I => \N__25040\
        );

    \I__3544\ : InMux
    port map (
            O => \N__25080\,
            I => \N__25040\
        );

    \I__3543\ : InMux
    port map (
            O => \N__25079\,
            I => \N__25040\
        );

    \I__3542\ : InMux
    port map (
            O => \N__25078\,
            I => \N__25031\
        );

    \I__3541\ : InMux
    port map (
            O => \N__25077\,
            I => \N__25031\
        );

    \I__3540\ : InMux
    port map (
            O => \N__25076\,
            I => \N__25031\
        );

    \I__3539\ : InMux
    port map (
            O => \N__25075\,
            I => \N__25031\
        );

    \I__3538\ : InMux
    port map (
            O => \N__25074\,
            I => \N__25022\
        );

    \I__3537\ : InMux
    port map (
            O => \N__25073\,
            I => \N__25022\
        );

    \I__3536\ : InMux
    port map (
            O => \N__25072\,
            I => \N__25022\
        );

    \I__3535\ : InMux
    port map (
            O => \N__25071\,
            I => \N__25022\
        );

    \I__3534\ : InMux
    port map (
            O => \N__25070\,
            I => \N__25013\
        );

    \I__3533\ : InMux
    port map (
            O => \N__25069\,
            I => \N__25013\
        );

    \I__3532\ : InMux
    port map (
            O => \N__25068\,
            I => \N__25013\
        );

    \I__3531\ : InMux
    port map (
            O => \N__25067\,
            I => \N__25013\
        );

    \I__3530\ : InMux
    port map (
            O => \N__25066\,
            I => \N__25004\
        );

    \I__3529\ : InMux
    port map (
            O => \N__25065\,
            I => \N__25004\
        );

    \I__3528\ : InMux
    port map (
            O => \N__25064\,
            I => \N__25004\
        );

    \I__3527\ : InMux
    port map (
            O => \N__25063\,
            I => \N__25004\
        );

    \I__3526\ : LocalMux
    port map (
            O => \N__25054\,
            I => \N__24997\
        );

    \I__3525\ : Span4Mux_h
    port map (
            O => \N__25049\,
            I => \N__24997\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__25040\,
            I => \N__24997\
        );

    \I__3523\ : LocalMux
    port map (
            O => \N__25031\,
            I => \N__24988\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__25022\,
            I => \N__24988\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__25013\,
            I => \N__24988\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__25004\,
            I => \N__24988\
        );

    \I__3519\ : Odrv4
    port map (
            O => \N__24997\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__3518\ : Odrv12
    port map (
            O => \N__24988\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__3517\ : InMux
    port map (
            O => \N__24983\,
            I => \N__24980\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__24980\,
            I => \phase_controller_inst2.start_timer_tr_RNO_0_0\
        );

    \I__3515\ : CascadeMux
    port map (
            O => \N__24977\,
            I => \N__24971\
        );

    \I__3514\ : InMux
    port map (
            O => \N__24976\,
            I => \N__24968\
        );

    \I__3513\ : InMux
    port map (
            O => \N__24975\,
            I => \N__24963\
        );

    \I__3512\ : InMux
    port map (
            O => \N__24974\,
            I => \N__24963\
        );

    \I__3511\ : InMux
    port map (
            O => \N__24971\,
            I => \N__24960\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__24968\,
            I => \N__24957\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__24963\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__24960\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__3507\ : Odrv4
    port map (
            O => \N__24957\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__3506\ : InMux
    port map (
            O => \N__24950\,
            I => \N__24946\
        );

    \I__3505\ : InMux
    port map (
            O => \N__24949\,
            I => \N__24942\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__24946\,
            I => \N__24939\
        );

    \I__3503\ : InMux
    port map (
            O => \N__24945\,
            I => \N__24936\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__24942\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__3501\ : Odrv4
    port map (
            O => \N__24939\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__3500\ : LocalMux
    port map (
            O => \N__24936\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__3499\ : InMux
    port map (
            O => \N__24929\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_22\
        );

    \I__3498\ : InMux
    port map (
            O => \N__24926\,
            I => \bfn_7_10_0_\
        );

    \I__3497\ : InMux
    port map (
            O => \N__24923\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_24\
        );

    \I__3496\ : InMux
    port map (
            O => \N__24920\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_25\
        );

    \I__3495\ : InMux
    port map (
            O => \N__24917\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_26\
        );

    \I__3494\ : InMux
    port map (
            O => \N__24914\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_27\
        );

    \I__3493\ : InMux
    port map (
            O => \N__24911\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_28\
        );

    \I__3492\ : InMux
    port map (
            O => \N__24908\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_13\
        );

    \I__3491\ : InMux
    port map (
            O => \N__24905\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_14\
        );

    \I__3490\ : InMux
    port map (
            O => \N__24902\,
            I => \bfn_7_9_0_\
        );

    \I__3489\ : InMux
    port map (
            O => \N__24899\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_16\
        );

    \I__3488\ : InMux
    port map (
            O => \N__24896\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_17\
        );

    \I__3487\ : InMux
    port map (
            O => \N__24893\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_18\
        );

    \I__3486\ : InMux
    port map (
            O => \N__24890\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_19\
        );

    \I__3485\ : InMux
    port map (
            O => \N__24887\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_20\
        );

    \I__3484\ : InMux
    port map (
            O => \N__24884\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_21\
        );

    \I__3483\ : InMux
    port map (
            O => \N__24881\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_4\
        );

    \I__3482\ : InMux
    port map (
            O => \N__24878\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_5\
        );

    \I__3481\ : InMux
    port map (
            O => \N__24875\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_6\
        );

    \I__3480\ : InMux
    port map (
            O => \N__24872\,
            I => \bfn_7_8_0_\
        );

    \I__3479\ : InMux
    port map (
            O => \N__24869\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_8\
        );

    \I__3478\ : InMux
    port map (
            O => \N__24866\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_9\
        );

    \I__3477\ : InMux
    port map (
            O => \N__24863\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_10\
        );

    \I__3476\ : InMux
    port map (
            O => \N__24860\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_11\
        );

    \I__3475\ : InMux
    port map (
            O => \N__24857\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_12\
        );

    \I__3474\ : InMux
    port map (
            O => \N__24854\,
            I => \N__24849\
        );

    \I__3473\ : InMux
    port map (
            O => \N__24853\,
            I => \N__24846\
        );

    \I__3472\ : InMux
    port map (
            O => \N__24852\,
            I => \N__24843\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__24849\,
            I => \N__24840\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__24846\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__24843\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__3468\ : Odrv12
    port map (
            O => \N__24840\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__3467\ : InMux
    port map (
            O => \N__24833\,
            I => \pwm_generator_inst.counter_cry_6\
        );

    \I__3466\ : InMux
    port map (
            O => \N__24830\,
            I => \N__24825\
        );

    \I__3465\ : InMux
    port map (
            O => \N__24829\,
            I => \N__24822\
        );

    \I__3464\ : InMux
    port map (
            O => \N__24828\,
            I => \N__24819\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__24825\,
            I => \N__24816\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__24822\,
            I => \N__24813\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__24819\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__3460\ : Odrv4
    port map (
            O => \N__24816\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__3459\ : Odrv4
    port map (
            O => \N__24813\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__3458\ : InMux
    port map (
            O => \N__24806\,
            I => \bfn_5_27_0_\
        );

    \I__3457\ : InMux
    port map (
            O => \N__24803\,
            I => \N__24785\
        );

    \I__3456\ : InMux
    port map (
            O => \N__24802\,
            I => \N__24785\
        );

    \I__3455\ : InMux
    port map (
            O => \N__24801\,
            I => \N__24785\
        );

    \I__3454\ : InMux
    port map (
            O => \N__24800\,
            I => \N__24785\
        );

    \I__3453\ : InMux
    port map (
            O => \N__24799\,
            I => \N__24780\
        );

    \I__3452\ : InMux
    port map (
            O => \N__24798\,
            I => \N__24780\
        );

    \I__3451\ : InMux
    port map (
            O => \N__24797\,
            I => \N__24771\
        );

    \I__3450\ : InMux
    port map (
            O => \N__24796\,
            I => \N__24771\
        );

    \I__3449\ : InMux
    port map (
            O => \N__24795\,
            I => \N__24771\
        );

    \I__3448\ : InMux
    port map (
            O => \N__24794\,
            I => \N__24771\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__24785\,
            I => \N__24766\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__24780\,
            I => \N__24766\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__24771\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__3444\ : Odrv4
    port map (
            O => \N__24766\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__3443\ : InMux
    port map (
            O => \N__24761\,
            I => \pwm_generator_inst.counter_cry_8\
        );

    \I__3442\ : InMux
    port map (
            O => \N__24758\,
            I => \N__24753\
        );

    \I__3441\ : InMux
    port map (
            O => \N__24757\,
            I => \N__24750\
        );

    \I__3440\ : InMux
    port map (
            O => \N__24756\,
            I => \N__24747\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__24753\,
            I => \N__24744\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__24750\,
            I => \N__24741\
        );

    \I__3437\ : LocalMux
    port map (
            O => \N__24747\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__3436\ : Odrv4
    port map (
            O => \N__24744\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__3435\ : Odrv4
    port map (
            O => \N__24741\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__3434\ : InMux
    port map (
            O => \N__24734\,
            I => \bfn_7_7_0_\
        );

    \I__3433\ : InMux
    port map (
            O => \N__24731\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_0\
        );

    \I__3432\ : InMux
    port map (
            O => \N__24728\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_1\
        );

    \I__3431\ : InMux
    port map (
            O => \N__24725\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_2\
        );

    \I__3430\ : InMux
    port map (
            O => \N__24722\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_3\
        );

    \I__3429\ : CascadeMux
    port map (
            O => \N__24719\,
            I => \pwm_generator_inst.un1_counterlto2_0_cascade_\
        );

    \I__3428\ : InMux
    port map (
            O => \N__24716\,
            I => \N__24713\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__24713\,
            I => \pwm_generator_inst.un1_counterlt9\
        );

    \I__3426\ : InMux
    port map (
            O => \N__24710\,
            I => \N__24706\
        );

    \I__3425\ : InMux
    port map (
            O => \N__24709\,
            I => \N__24702\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__24706\,
            I => \N__24699\
        );

    \I__3423\ : InMux
    port map (
            O => \N__24705\,
            I => \N__24696\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__24702\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__3421\ : Odrv4
    port map (
            O => \N__24699\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__24696\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__3419\ : InMux
    port map (
            O => \N__24689\,
            I => \bfn_5_26_0_\
        );

    \I__3418\ : InMux
    port map (
            O => \N__24686\,
            I => \N__24681\
        );

    \I__3417\ : InMux
    port map (
            O => \N__24685\,
            I => \N__24678\
        );

    \I__3416\ : InMux
    port map (
            O => \N__24684\,
            I => \N__24675\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__24681\,
            I => \N__24672\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__24678\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__24675\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__3412\ : Odrv4
    port map (
            O => \N__24672\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__3411\ : InMux
    port map (
            O => \N__24665\,
            I => \pwm_generator_inst.counter_cry_0\
        );

    \I__3410\ : InMux
    port map (
            O => \N__24662\,
            I => \N__24658\
        );

    \I__3409\ : InMux
    port map (
            O => \N__24661\,
            I => \N__24654\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__24658\,
            I => \N__24651\
        );

    \I__3407\ : InMux
    port map (
            O => \N__24657\,
            I => \N__24648\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__24654\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__3405\ : Odrv4
    port map (
            O => \N__24651\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__24648\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__3403\ : InMux
    port map (
            O => \N__24641\,
            I => \pwm_generator_inst.counter_cry_1\
        );

    \I__3402\ : InMux
    port map (
            O => \N__24638\,
            I => \N__24633\
        );

    \I__3401\ : InMux
    port map (
            O => \N__24637\,
            I => \N__24630\
        );

    \I__3400\ : InMux
    port map (
            O => \N__24636\,
            I => \N__24627\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__24633\,
            I => \N__24624\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__24630\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__24627\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__3396\ : Odrv4
    port map (
            O => \N__24624\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__3395\ : InMux
    port map (
            O => \N__24617\,
            I => \pwm_generator_inst.counter_cry_2\
        );

    \I__3394\ : InMux
    port map (
            O => \N__24614\,
            I => \N__24609\
        );

    \I__3393\ : InMux
    port map (
            O => \N__24613\,
            I => \N__24606\
        );

    \I__3392\ : InMux
    port map (
            O => \N__24612\,
            I => \N__24603\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__24609\,
            I => \N__24600\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__24606\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__24603\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__3388\ : Odrv4
    port map (
            O => \N__24600\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__3387\ : InMux
    port map (
            O => \N__24593\,
            I => \pwm_generator_inst.counter_cry_3\
        );

    \I__3386\ : InMux
    port map (
            O => \N__24590\,
            I => \N__24585\
        );

    \I__3385\ : InMux
    port map (
            O => \N__24589\,
            I => \N__24582\
        );

    \I__3384\ : InMux
    port map (
            O => \N__24588\,
            I => \N__24579\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__24585\,
            I => \N__24576\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__24582\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__24579\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__3380\ : Odrv4
    port map (
            O => \N__24576\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__3379\ : InMux
    port map (
            O => \N__24569\,
            I => \pwm_generator_inst.counter_cry_4\
        );

    \I__3378\ : InMux
    port map (
            O => \N__24566\,
            I => \N__24561\
        );

    \I__3377\ : InMux
    port map (
            O => \N__24565\,
            I => \N__24558\
        );

    \I__3376\ : InMux
    port map (
            O => \N__24564\,
            I => \N__24555\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__24561\,
            I => \N__24552\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__24558\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__24555\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__3372\ : Odrv12
    port map (
            O => \N__24552\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__3371\ : InMux
    port map (
            O => \N__24545\,
            I => \pwm_generator_inst.counter_cry_5\
        );

    \I__3370\ : CascadeMux
    port map (
            O => \N__24542\,
            I => \N__24539\
        );

    \I__3369\ : InMux
    port map (
            O => \N__24539\,
            I => \N__24536\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__24536\,
            I => \pwm_generator_inst.un14_counter_6\
        );

    \I__3367\ : InMux
    port map (
            O => \N__24533\,
            I => \N__24530\
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__24530\,
            I => \pwm_generator_inst.counter_i_6\
        );

    \I__3365\ : InMux
    port map (
            O => \N__24527\,
            I => \N__24524\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__24524\,
            I => \pwm_generator_inst.un14_counter_7\
        );

    \I__3363\ : CascadeMux
    port map (
            O => \N__24521\,
            I => \N__24518\
        );

    \I__3362\ : InMux
    port map (
            O => \N__24518\,
            I => \N__24515\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__24515\,
            I => \pwm_generator_inst.counter_i_7\
        );

    \I__3360\ : CascadeMux
    port map (
            O => \N__24512\,
            I => \N__24509\
        );

    \I__3359\ : InMux
    port map (
            O => \N__24509\,
            I => \N__24506\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__24506\,
            I => \pwm_generator_inst.un14_counter_8\
        );

    \I__3357\ : InMux
    port map (
            O => \N__24503\,
            I => \N__24500\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__24500\,
            I => \pwm_generator_inst.counter_i_8\
        );

    \I__3355\ : CascadeMux
    port map (
            O => \N__24497\,
            I => \N__24494\
        );

    \I__3354\ : InMux
    port map (
            O => \N__24494\,
            I => \N__24491\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__24491\,
            I => \N__24488\
        );

    \I__3352\ : Odrv4
    port map (
            O => \N__24488\,
            I => \pwm_generator_inst.threshold_9\
        );

    \I__3351\ : InMux
    port map (
            O => \N__24485\,
            I => \N__24482\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__24482\,
            I => \pwm_generator_inst.counter_i_9\
        );

    \I__3349\ : InMux
    port map (
            O => \N__24479\,
            I => \pwm_generator_inst.un14_counter_cry_9\
        );

    \I__3348\ : IoInMux
    port map (
            O => \N__24476\,
            I => \N__24473\
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__24473\,
            I => \N__24470\
        );

    \I__3346\ : Span4Mux_s1_v
    port map (
            O => \N__24470\,
            I => \N__24467\
        );

    \I__3345\ : Span4Mux_h
    port map (
            O => \N__24467\,
            I => \N__24464\
        );

    \I__3344\ : Sp12to4
    port map (
            O => \N__24464\,
            I => \N__24461\
        );

    \I__3343\ : Span12Mux_h
    port map (
            O => \N__24461\,
            I => \N__24458\
        );

    \I__3342\ : Span12Mux_v
    port map (
            O => \N__24458\,
            I => \N__24455\
        );

    \I__3341\ : Odrv12
    port map (
            O => \N__24455\,
            I => pwm_output_c
        );

    \I__3340\ : InMux
    port map (
            O => \N__24452\,
            I => \N__24449\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__24449\,
            I => \N__24446\
        );

    \I__3338\ : Span4Mux_s3_v
    port map (
            O => \N__24446\,
            I => \N__24443\
        );

    \I__3337\ : Span4Mux_h
    port map (
            O => \N__24443\,
            I => \N__24440\
        );

    \I__3336\ : Odrv4
    port map (
            O => \N__24440\,
            I => \N_38_i_i\
        );

    \I__3335\ : CascadeMux
    port map (
            O => \N__24437\,
            I => \pwm_generator_inst.un1_counterlto9_2_cascade_\
        );

    \I__3334\ : InMux
    port map (
            O => \N__24434\,
            I => \N__24431\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__24431\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\
        );

    \I__3332\ : InMux
    port map (
            O => \N__24428\,
            I => \N__24425\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__24425\,
            I => \N__24422\
        );

    \I__3330\ : Odrv12
    port map (
            O => \N__24422\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\
        );

    \I__3329\ : CascadeMux
    port map (
            O => \N__24419\,
            I => \N__24416\
        );

    \I__3328\ : InMux
    port map (
            O => \N__24416\,
            I => \N__24413\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__24413\,
            I => \pwm_generator_inst.threshold_0\
        );

    \I__3326\ : InMux
    port map (
            O => \N__24410\,
            I => \N__24407\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__24407\,
            I => \pwm_generator_inst.counter_i_0\
        );

    \I__3324\ : CascadeMux
    port map (
            O => \N__24404\,
            I => \N__24401\
        );

    \I__3323\ : InMux
    port map (
            O => \N__24401\,
            I => \N__24398\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__24398\,
            I => \pwm_generator_inst.un14_counter_1\
        );

    \I__3321\ : InMux
    port map (
            O => \N__24395\,
            I => \N__24392\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__24392\,
            I => \pwm_generator_inst.counter_i_1\
        );

    \I__3319\ : CascadeMux
    port map (
            O => \N__24389\,
            I => \N__24386\
        );

    \I__3318\ : InMux
    port map (
            O => \N__24386\,
            I => \N__24383\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__24383\,
            I => \pwm_generator_inst.threshold_2\
        );

    \I__3316\ : InMux
    port map (
            O => \N__24380\,
            I => \N__24377\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__24377\,
            I => \N__24374\
        );

    \I__3314\ : Odrv4
    port map (
            O => \N__24374\,
            I => \pwm_generator_inst.counter_i_2\
        );

    \I__3313\ : CascadeMux
    port map (
            O => \N__24371\,
            I => \N__24368\
        );

    \I__3312\ : InMux
    port map (
            O => \N__24368\,
            I => \N__24365\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__24365\,
            I => \pwm_generator_inst.threshold_3\
        );

    \I__3310\ : InMux
    port map (
            O => \N__24362\,
            I => \N__24359\
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__24359\,
            I => \pwm_generator_inst.counter_i_3\
        );

    \I__3308\ : InMux
    port map (
            O => \N__24356\,
            I => \N__24353\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__24353\,
            I => \pwm_generator_inst.threshold_4\
        );

    \I__3306\ : CascadeMux
    port map (
            O => \N__24350\,
            I => \N__24347\
        );

    \I__3305\ : InMux
    port map (
            O => \N__24347\,
            I => \N__24344\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__24344\,
            I => \pwm_generator_inst.counter_i_4\
        );

    \I__3303\ : CascadeMux
    port map (
            O => \N__24341\,
            I => \N__24338\
        );

    \I__3302\ : InMux
    port map (
            O => \N__24338\,
            I => \N__24335\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__24335\,
            I => \pwm_generator_inst.threshold_5\
        );

    \I__3300\ : InMux
    port map (
            O => \N__24332\,
            I => \N__24329\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__24329\,
            I => \pwm_generator_inst.counter_i_5\
        );

    \I__3298\ : InMux
    port map (
            O => \N__24326\,
            I => \N__24323\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__24323\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\
        );

    \I__3296\ : CascadeMux
    port map (
            O => \N__24320\,
            I => \N__24317\
        );

    \I__3295\ : InMux
    port map (
            O => \N__24317\,
            I => \N__24314\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__24314\,
            I => \N__24311\
        );

    \I__3293\ : Odrv4
    port map (
            O => \N__24311\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_28\
        );

    \I__3292\ : InMux
    port map (
            O => \N__24308\,
            I => \N__24305\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__24305\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_23\
        );

    \I__3290\ : InMux
    port map (
            O => \N__24302\,
            I => \N__24299\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__24299\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_24\
        );

    \I__3288\ : InMux
    port map (
            O => \N__24296\,
            I => \N__24293\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__24293\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_17\
        );

    \I__3286\ : CascadeMux
    port map (
            O => \N__24290\,
            I => \N__24287\
        );

    \I__3285\ : InMux
    port map (
            O => \N__24287\,
            I => \N__24284\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__24284\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_29\
        );

    \I__3283\ : InMux
    port map (
            O => \N__24281\,
            I => \N__24278\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__24278\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_26\
        );

    \I__3281\ : InMux
    port map (
            O => \N__24275\,
            I => \N__24272\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__24272\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_25\
        );

    \I__3279\ : InMux
    port map (
            O => \N__24269\,
            I => \N__24266\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__24266\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_30\
        );

    \I__3277\ : CascadeMux
    port map (
            O => \N__24263\,
            I => \N__24260\
        );

    \I__3276\ : InMux
    port map (
            O => \N__24260\,
            I => \N__24257\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__24257\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\
        );

    \I__3274\ : CascadeMux
    port map (
            O => \N__24254\,
            I => \N__24251\
        );

    \I__3273\ : InMux
    port map (
            O => \N__24251\,
            I => \N__24248\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__24248\,
            I => \N__24245\
        );

    \I__3271\ : Odrv4
    port map (
            O => \N__24245\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\
        );

    \I__3270\ : InMux
    port map (
            O => \N__24242\,
            I => \N__24239\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__24239\,
            I => \N__24235\
        );

    \I__3268\ : InMux
    port map (
            O => \N__24238\,
            I => \N__24232\
        );

    \I__3267\ : Odrv12
    port map (
            O => \N__24235\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__24232\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__3265\ : InMux
    port map (
            O => \N__24227\,
            I => \N__24224\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__24224\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\
        );

    \I__3263\ : InMux
    port map (
            O => \N__24221\,
            I => \N__24218\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__24218\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\
        );

    \I__3261\ : InMux
    port map (
            O => \N__24215\,
            I => \N__24212\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__24212\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\
        );

    \I__3259\ : CascadeMux
    port map (
            O => \N__24209\,
            I => \N__24206\
        );

    \I__3258\ : InMux
    port map (
            O => \N__24206\,
            I => \N__24203\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__24203\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_19\
        );

    \I__3256\ : InMux
    port map (
            O => \N__24200\,
            I => \N__24197\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__24197\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_21\
        );

    \I__3254\ : CascadeMux
    port map (
            O => \N__24194\,
            I => \N__24191\
        );

    \I__3253\ : InMux
    port map (
            O => \N__24191\,
            I => \N__24188\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__24188\,
            I => \N__24185\
        );

    \I__3251\ : Odrv4
    port map (
            O => \N__24185\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_27\
        );

    \I__3250\ : CascadeMux
    port map (
            O => \N__24182\,
            I => \N__24179\
        );

    \I__3249\ : InMux
    port map (
            O => \N__24179\,
            I => \N__24176\
        );

    \I__3248\ : LocalMux
    port map (
            O => \N__24176\,
            I => \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23\
        );

    \I__3247\ : InMux
    port map (
            O => \N__24173\,
            I => \N__24169\
        );

    \I__3246\ : InMux
    port map (
            O => \N__24172\,
            I => \N__24166\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__24169\,
            I => \N__24160\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__24166\,
            I => \N__24160\
        );

    \I__3243\ : InMux
    port map (
            O => \N__24165\,
            I => \N__24157\
        );

    \I__3242\ : Span4Mux_h
    port map (
            O => \N__24160\,
            I => \N__24154\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__24157\,
            I => \N__24151\
        );

    \I__3240\ : Odrv4
    port map (
            O => \N__24154\,
            I => pwm_duty_input_3
        );

    \I__3239\ : Odrv4
    port map (
            O => \N__24151\,
            I => pwm_duty_input_3
        );

    \I__3238\ : CascadeMux
    port map (
            O => \N__24146\,
            I => \N__24143\
        );

    \I__3237\ : InMux
    port map (
            O => \N__24143\,
            I => \N__24139\
        );

    \I__3236\ : InMux
    port map (
            O => \N__24142\,
            I => \N__24136\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__24139\,
            I => \N__24130\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__24136\,
            I => \N__24130\
        );

    \I__3233\ : InMux
    port map (
            O => \N__24135\,
            I => \N__24127\
        );

    \I__3232\ : Span4Mux_h
    port map (
            O => \N__24130\,
            I => \N__24124\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__24127\,
            I => \N__24121\
        );

    \I__3230\ : Odrv4
    port map (
            O => \N__24124\,
            I => pwm_duty_input_4
        );

    \I__3229\ : Odrv4
    port map (
            O => \N__24121\,
            I => pwm_duty_input_4
        );

    \I__3228\ : CascadeMux
    port map (
            O => \N__24116\,
            I => \N__24113\
        );

    \I__3227\ : InMux
    port map (
            O => \N__24113\,
            I => \N__24110\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__24110\,
            I => \N__24105\
        );

    \I__3225\ : InMux
    port map (
            O => \N__24109\,
            I => \N__24102\
        );

    \I__3224\ : InMux
    port map (
            O => \N__24108\,
            I => \N__24099\
        );

    \I__3223\ : Span4Mux_h
    port map (
            O => \N__24105\,
            I => \N__24096\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__24102\,
            I => \N__24093\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__24099\,
            I => \N__24090\
        );

    \I__3220\ : Odrv4
    port map (
            O => \N__24096\,
            I => pwm_duty_input_5
        );

    \I__3219\ : Odrv4
    port map (
            O => \N__24093\,
            I => pwm_duty_input_5
        );

    \I__3218\ : Odrv4
    port map (
            O => \N__24090\,
            I => pwm_duty_input_5
        );

    \I__3217\ : InMux
    port map (
            O => \N__24083\,
            I => \N__24080\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__24080\,
            I => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\
        );

    \I__3215\ : InMux
    port map (
            O => \N__24077\,
            I => \N__24066\
        );

    \I__3214\ : InMux
    port map (
            O => \N__24076\,
            I => \N__24049\
        );

    \I__3213\ : InMux
    port map (
            O => \N__24075\,
            I => \N__24049\
        );

    \I__3212\ : InMux
    port map (
            O => \N__24074\,
            I => \N__24049\
        );

    \I__3211\ : InMux
    port map (
            O => \N__24073\,
            I => \N__24049\
        );

    \I__3210\ : InMux
    port map (
            O => \N__24072\,
            I => \N__24049\
        );

    \I__3209\ : InMux
    port map (
            O => \N__24071\,
            I => \N__24049\
        );

    \I__3208\ : InMux
    port map (
            O => \N__24070\,
            I => \N__24049\
        );

    \I__3207\ : InMux
    port map (
            O => \N__24069\,
            I => \N__24049\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__24066\,
            I => \pwm_generator_inst.N_17\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__24049\,
            I => \pwm_generator_inst.N_17\
        );

    \I__3204\ : CascadeMux
    port map (
            O => \N__24044\,
            I => \N__24035\
        );

    \I__3203\ : CascadeMux
    port map (
            O => \N__24043\,
            I => \N__24030\
        );

    \I__3202\ : CascadeMux
    port map (
            O => \N__24042\,
            I => \N__24027\
        );

    \I__3201\ : CascadeMux
    port map (
            O => \N__24041\,
            I => \N__24023\
        );

    \I__3200\ : InMux
    port map (
            O => \N__24040\,
            I => \N__24020\
        );

    \I__3199\ : InMux
    port map (
            O => \N__24039\,
            I => \N__24017\
        );

    \I__3198\ : InMux
    port map (
            O => \N__24038\,
            I => \N__24000\
        );

    \I__3197\ : InMux
    port map (
            O => \N__24035\,
            I => \N__24000\
        );

    \I__3196\ : InMux
    port map (
            O => \N__24034\,
            I => \N__24000\
        );

    \I__3195\ : InMux
    port map (
            O => \N__24033\,
            I => \N__24000\
        );

    \I__3194\ : InMux
    port map (
            O => \N__24030\,
            I => \N__24000\
        );

    \I__3193\ : InMux
    port map (
            O => \N__24027\,
            I => \N__24000\
        );

    \I__3192\ : InMux
    port map (
            O => \N__24026\,
            I => \N__24000\
        );

    \I__3191\ : InMux
    port map (
            O => \N__24023\,
            I => \N__24000\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__24020\,
            I => \pwm_generator_inst.N_16\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__24017\,
            I => \pwm_generator_inst.N_16\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__24000\,
            I => \pwm_generator_inst.N_16\
        );

    \I__3187\ : InMux
    port map (
            O => \N__23993\,
            I => \N__23990\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__23990\,
            I => \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033\
        );

    \I__3185\ : CascadeMux
    port map (
            O => \N__23987\,
            I => \pwm_generator_inst.N_17_cascade_\
        );

    \I__3184\ : InMux
    port map (
            O => \N__23984\,
            I => \N__23980\
        );

    \I__3183\ : CascadeMux
    port map (
            O => \N__23983\,
            I => \N__23977\
        );

    \I__3182\ : LocalMux
    port map (
            O => \N__23980\,
            I => \N__23973\
        );

    \I__3181\ : InMux
    port map (
            O => \N__23977\,
            I => \N__23970\
        );

    \I__3180\ : InMux
    port map (
            O => \N__23976\,
            I => \N__23967\
        );

    \I__3179\ : Span4Mux_v
    port map (
            O => \N__23973\,
            I => \N__23964\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__23970\,
            I => \N__23961\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__23967\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__3176\ : Odrv4
    port map (
            O => \N__23964\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__3175\ : Odrv4
    port map (
            O => \N__23961\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__3174\ : InMux
    port map (
            O => \N__23954\,
            I => \N__23951\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__23951\,
            I => \N__23948\
        );

    \I__3172\ : Odrv12
    port map (
            O => \N__23948\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\
        );

    \I__3171\ : CascadeMux
    port map (
            O => \N__23945\,
            I => \N__23942\
        );

    \I__3170\ : InMux
    port map (
            O => \N__23942\,
            I => \N__23938\
        );

    \I__3169\ : InMux
    port map (
            O => \N__23941\,
            I => \N__23935\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__23938\,
            I => \N__23932\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__23935\,
            I => \N__23929\
        );

    \I__3166\ : Span4Mux_v
    port map (
            O => \N__23932\,
            I => \N__23926\
        );

    \I__3165\ : Span4Mux_h
    port map (
            O => \N__23929\,
            I => \N__23923\
        );

    \I__3164\ : Odrv4
    port map (
            O => \N__23926\,
            I => \pwm_generator_inst.O_10\
        );

    \I__3163\ : Odrv4
    port map (
            O => \N__23923\,
            I => \pwm_generator_inst.O_10\
        );

    \I__3162\ : InMux
    port map (
            O => \N__23918\,
            I => \N__23915\
        );

    \I__3161\ : LocalMux
    port map (
            O => \N__23915\,
            I => \N__23912\
        );

    \I__3160\ : Span4Mux_h
    port map (
            O => \N__23912\,
            I => \N__23909\
        );

    \I__3159\ : Odrv4
    port map (
            O => \N__23909\,
            I => \pwm_generator_inst.un19_threshold_axb_0\
        );

    \I__3158\ : InMux
    port map (
            O => \N__23906\,
            I => \N__23903\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__23903\,
            I => \N__23900\
        );

    \I__3156\ : Glb2LocalMux
    port map (
            O => \N__23900\,
            I => \N__23897\
        );

    \I__3155\ : GlobalMux
    port map (
            O => \N__23897\,
            I => clk_12mhz
        );

    \I__3154\ : IoInMux
    port map (
            O => \N__23894\,
            I => \N__23891\
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__23891\,
            I => \N__23888\
        );

    \I__3152\ : IoSpan4Mux
    port map (
            O => \N__23888\,
            I => \N__23885\
        );

    \I__3151\ : Span4Mux_s0_v
    port map (
            O => \N__23885\,
            I => \N__23882\
        );

    \I__3150\ : Odrv4
    port map (
            O => \N__23882\,
            I => \GB_BUFFER_clk_12mhz_THRU_CO\
        );

    \I__3149\ : InMux
    port map (
            O => \N__23879\,
            I => \N__23874\
        );

    \I__3148\ : InMux
    port map (
            O => \N__23878\,
            I => \N__23860\
        );

    \I__3147\ : InMux
    port map (
            O => \N__23877\,
            I => \N__23860\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__23874\,
            I => \N__23857\
        );

    \I__3145\ : InMux
    port map (
            O => \N__23873\,
            I => \N__23852\
        );

    \I__3144\ : InMux
    port map (
            O => \N__23872\,
            I => \N__23852\
        );

    \I__3143\ : InMux
    port map (
            O => \N__23871\,
            I => \N__23839\
        );

    \I__3142\ : InMux
    port map (
            O => \N__23870\,
            I => \N__23833\
        );

    \I__3141\ : InMux
    port map (
            O => \N__23869\,
            I => \N__23830\
        );

    \I__3140\ : InMux
    port map (
            O => \N__23868\,
            I => \N__23827\
        );

    \I__3139\ : InMux
    port map (
            O => \N__23867\,
            I => \N__23820\
        );

    \I__3138\ : InMux
    port map (
            O => \N__23866\,
            I => \N__23820\
        );

    \I__3137\ : InMux
    port map (
            O => \N__23865\,
            I => \N__23820\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__23860\,
            I => \N__23813\
        );

    \I__3135\ : Span4Mux_h
    port map (
            O => \N__23857\,
            I => \N__23813\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__23852\,
            I => \N__23813\
        );

    \I__3133\ : InMux
    port map (
            O => \N__23851\,
            I => \N__23810\
        );

    \I__3132\ : InMux
    port map (
            O => \N__23850\,
            I => \N__23805\
        );

    \I__3131\ : InMux
    port map (
            O => \N__23849\,
            I => \N__23805\
        );

    \I__3130\ : InMux
    port map (
            O => \N__23848\,
            I => \N__23785\
        );

    \I__3129\ : InMux
    port map (
            O => \N__23847\,
            I => \N__23785\
        );

    \I__3128\ : InMux
    port map (
            O => \N__23846\,
            I => \N__23785\
        );

    \I__3127\ : InMux
    port map (
            O => \N__23845\,
            I => \N__23785\
        );

    \I__3126\ : InMux
    port map (
            O => \N__23844\,
            I => \N__23785\
        );

    \I__3125\ : InMux
    port map (
            O => \N__23843\,
            I => \N__23785\
        );

    \I__3124\ : InMux
    port map (
            O => \N__23842\,
            I => \N__23785\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__23839\,
            I => \N__23782\
        );

    \I__3122\ : InMux
    port map (
            O => \N__23838\,
            I => \N__23775\
        );

    \I__3121\ : InMux
    port map (
            O => \N__23837\,
            I => \N__23775\
        );

    \I__3120\ : InMux
    port map (
            O => \N__23836\,
            I => \N__23775\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__23833\,
            I => \N__23766\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__23830\,
            I => \N__23766\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__23827\,
            I => \N__23766\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__23820\,
            I => \N__23766\
        );

    \I__3115\ : Span4Mux_h
    port map (
            O => \N__23813\,
            I => \N__23763\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__23810\,
            I => \N__23758\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__23805\,
            I => \N__23755\
        );

    \I__3112\ : InMux
    port map (
            O => \N__23804\,
            I => \N__23752\
        );

    \I__3111\ : InMux
    port map (
            O => \N__23803\,
            I => \N__23743\
        );

    \I__3110\ : InMux
    port map (
            O => \N__23802\,
            I => \N__23743\
        );

    \I__3109\ : InMux
    port map (
            O => \N__23801\,
            I => \N__23743\
        );

    \I__3108\ : InMux
    port map (
            O => \N__23800\,
            I => \N__23743\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__23785\,
            I => \N__23738\
        );

    \I__3106\ : Span4Mux_h
    port map (
            O => \N__23782\,
            I => \N__23738\
        );

    \I__3105\ : LocalMux
    port map (
            O => \N__23775\,
            I => \N__23731\
        );

    \I__3104\ : Span4Mux_v
    port map (
            O => \N__23766\,
            I => \N__23731\
        );

    \I__3103\ : Span4Mux_v
    port map (
            O => \N__23763\,
            I => \N__23731\
        );

    \I__3102\ : InMux
    port map (
            O => \N__23762\,
            I => \N__23728\
        );

    \I__3101\ : InMux
    port map (
            O => \N__23761\,
            I => \N__23725\
        );

    \I__3100\ : Span4Mux_h
    port map (
            O => \N__23758\,
            I => \N__23718\
        );

    \I__3099\ : Span4Mux_v
    port map (
            O => \N__23755\,
            I => \N__23718\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__23752\,
            I => \N__23718\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__23743\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3096\ : Odrv4
    port map (
            O => \N__23738\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3095\ : Odrv4
    port map (
            O => \N__23731\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__23728\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__23725\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3092\ : Odrv4
    port map (
            O => \N__23718\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3091\ : InMux
    port map (
            O => \N__23705\,
            I => \N__23691\
        );

    \I__3090\ : InMux
    port map (
            O => \N__23704\,
            I => \N__23691\
        );

    \I__3089\ : InMux
    port map (
            O => \N__23703\,
            I => \N__23691\
        );

    \I__3088\ : CascadeMux
    port map (
            O => \N__23702\,
            I => \N__23679\
        );

    \I__3087\ : CascadeMux
    port map (
            O => \N__23701\,
            I => \N__23675\
        );

    \I__3086\ : InMux
    port map (
            O => \N__23700\,
            I => \N__23668\
        );

    \I__3085\ : InMux
    port map (
            O => \N__23699\,
            I => \N__23668\
        );

    \I__3084\ : InMux
    port map (
            O => \N__23698\,
            I => \N__23668\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__23691\,
            I => \N__23665\
        );

    \I__3082\ : InMux
    port map (
            O => \N__23690\,
            I => \N__23662\
        );

    \I__3081\ : CascadeMux
    port map (
            O => \N__23689\,
            I => \N__23648\
        );

    \I__3080\ : CascadeMux
    port map (
            O => \N__23688\,
            I => \N__23643\
        );

    \I__3079\ : InMux
    port map (
            O => \N__23687\,
            I => \N__23640\
        );

    \I__3078\ : InMux
    port map (
            O => \N__23686\,
            I => \N__23637\
        );

    \I__3077\ : InMux
    port map (
            O => \N__23685\,
            I => \N__23630\
        );

    \I__3076\ : InMux
    port map (
            O => \N__23684\,
            I => \N__23630\
        );

    \I__3075\ : InMux
    port map (
            O => \N__23683\,
            I => \N__23630\
        );

    \I__3074\ : InMux
    port map (
            O => \N__23682\,
            I => \N__23625\
        );

    \I__3073\ : InMux
    port map (
            O => \N__23679\,
            I => \N__23625\
        );

    \I__3072\ : InMux
    port map (
            O => \N__23678\,
            I => \N__23620\
        );

    \I__3071\ : InMux
    port map (
            O => \N__23675\,
            I => \N__23620\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__23668\,
            I => \N__23617\
        );

    \I__3069\ : Span4Mux_v
    port map (
            O => \N__23665\,
            I => \N__23614\
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__23662\,
            I => \N__23611\
        );

    \I__3067\ : InMux
    port map (
            O => \N__23661\,
            I => \N__23608\
        );

    \I__3066\ : InMux
    port map (
            O => \N__23660\,
            I => \N__23593\
        );

    \I__3065\ : InMux
    port map (
            O => \N__23659\,
            I => \N__23593\
        );

    \I__3064\ : InMux
    port map (
            O => \N__23658\,
            I => \N__23593\
        );

    \I__3063\ : InMux
    port map (
            O => \N__23657\,
            I => \N__23593\
        );

    \I__3062\ : InMux
    port map (
            O => \N__23656\,
            I => \N__23593\
        );

    \I__3061\ : InMux
    port map (
            O => \N__23655\,
            I => \N__23593\
        );

    \I__3060\ : InMux
    port map (
            O => \N__23654\,
            I => \N__23593\
        );

    \I__3059\ : InMux
    port map (
            O => \N__23653\,
            I => \N__23584\
        );

    \I__3058\ : InMux
    port map (
            O => \N__23652\,
            I => \N__23584\
        );

    \I__3057\ : InMux
    port map (
            O => \N__23651\,
            I => \N__23584\
        );

    \I__3056\ : InMux
    port map (
            O => \N__23648\,
            I => \N__23584\
        );

    \I__3055\ : InMux
    port map (
            O => \N__23647\,
            I => \N__23577\
        );

    \I__3054\ : InMux
    port map (
            O => \N__23646\,
            I => \N__23577\
        );

    \I__3053\ : InMux
    port map (
            O => \N__23643\,
            I => \N__23577\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__23640\,
            I => \N__23574\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__23637\,
            I => \N__23571\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__23630\,
            I => \N__23568\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__23625\,
            I => \N__23563\
        );

    \I__3048\ : LocalMux
    port map (
            O => \N__23620\,
            I => \N__23563\
        );

    \I__3047\ : Span4Mux_v
    port map (
            O => \N__23617\,
            I => \N__23556\
        );

    \I__3046\ : Span4Mux_s2_h
    port map (
            O => \N__23614\,
            I => \N__23556\
        );

    \I__3045\ : Span4Mux_v
    port map (
            O => \N__23611\,
            I => \N__23556\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__23608\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__23593\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__23584\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__23577\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__3040\ : Odrv4
    port map (
            O => \N__23574\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__3039\ : Odrv4
    port map (
            O => \N__23571\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__3038\ : Odrv4
    port map (
            O => \N__23568\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__3037\ : Odrv4
    port map (
            O => \N__23563\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__3036\ : Odrv4
    port map (
            O => \N__23556\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__3035\ : CascadeMux
    port map (
            O => \N__23537\,
            I => \N__23534\
        );

    \I__3034\ : InMux
    port map (
            O => \N__23534\,
            I => \N__23531\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__23531\,
            I => \N__23528\
        );

    \I__3032\ : Span4Mux_h
    port map (
            O => \N__23528\,
            I => \N__23525\
        );

    \I__3031\ : Odrv4
    port map (
            O => \N__23525\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\
        );

    \I__3030\ : CascadeMux
    port map (
            O => \N__23522\,
            I => \N__23496\
        );

    \I__3029\ : CascadeMux
    port map (
            O => \N__23521\,
            I => \N__23493\
        );

    \I__3028\ : CascadeMux
    port map (
            O => \N__23520\,
            I => \N__23490\
        );

    \I__3027\ : CascadeMux
    port map (
            O => \N__23519\,
            I => \N__23487\
        );

    \I__3026\ : InMux
    port map (
            O => \N__23518\,
            I => \N__23484\
        );

    \I__3025\ : InMux
    port map (
            O => \N__23517\,
            I => \N__23477\
        );

    \I__3024\ : InMux
    port map (
            O => \N__23516\,
            I => \N__23477\
        );

    \I__3023\ : InMux
    port map (
            O => \N__23515\,
            I => \N__23477\
        );

    \I__3022\ : CascadeMux
    port map (
            O => \N__23514\,
            I => \N__23473\
        );

    \I__3021\ : CascadeMux
    port map (
            O => \N__23513\,
            I => \N__23470\
        );

    \I__3020\ : InMux
    port map (
            O => \N__23512\,
            I => \N__23467\
        );

    \I__3019\ : InMux
    port map (
            O => \N__23511\,
            I => \N__23464\
        );

    \I__3018\ : InMux
    port map (
            O => \N__23510\,
            I => \N__23461\
        );

    \I__3017\ : CascadeMux
    port map (
            O => \N__23509\,
            I => \N__23456\
        );

    \I__3016\ : InMux
    port map (
            O => \N__23508\,
            I => \N__23447\
        );

    \I__3015\ : InMux
    port map (
            O => \N__23507\,
            I => \N__23447\
        );

    \I__3014\ : InMux
    port map (
            O => \N__23506\,
            I => \N__23440\
        );

    \I__3013\ : InMux
    port map (
            O => \N__23505\,
            I => \N__23440\
        );

    \I__3012\ : InMux
    port map (
            O => \N__23504\,
            I => \N__23440\
        );

    \I__3011\ : InMux
    port map (
            O => \N__23503\,
            I => \N__23435\
        );

    \I__3010\ : InMux
    port map (
            O => \N__23502\,
            I => \N__23435\
        );

    \I__3009\ : InMux
    port map (
            O => \N__23501\,
            I => \N__23420\
        );

    \I__3008\ : InMux
    port map (
            O => \N__23500\,
            I => \N__23420\
        );

    \I__3007\ : InMux
    port map (
            O => \N__23499\,
            I => \N__23420\
        );

    \I__3006\ : InMux
    port map (
            O => \N__23496\,
            I => \N__23420\
        );

    \I__3005\ : InMux
    port map (
            O => \N__23493\,
            I => \N__23420\
        );

    \I__3004\ : InMux
    port map (
            O => \N__23490\,
            I => \N__23420\
        );

    \I__3003\ : InMux
    port map (
            O => \N__23487\,
            I => \N__23420\
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__23484\,
            I => \N__23415\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__23477\,
            I => \N__23415\
        );

    \I__3000\ : InMux
    port map (
            O => \N__23476\,
            I => \N__23408\
        );

    \I__2999\ : InMux
    port map (
            O => \N__23473\,
            I => \N__23408\
        );

    \I__2998\ : InMux
    port map (
            O => \N__23470\,
            I => \N__23408\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__23467\,
            I => \N__23401\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__23464\,
            I => \N__23401\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__23461\,
            I => \N__23401\
        );

    \I__2994\ : InMux
    port map (
            O => \N__23460\,
            I => \N__23394\
        );

    \I__2993\ : InMux
    port map (
            O => \N__23459\,
            I => \N__23394\
        );

    \I__2992\ : InMux
    port map (
            O => \N__23456\,
            I => \N__23394\
        );

    \I__2991\ : InMux
    port map (
            O => \N__23455\,
            I => \N__23385\
        );

    \I__2990\ : InMux
    port map (
            O => \N__23454\,
            I => \N__23385\
        );

    \I__2989\ : InMux
    port map (
            O => \N__23453\,
            I => \N__23385\
        );

    \I__2988\ : InMux
    port map (
            O => \N__23452\,
            I => \N__23385\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__23447\,
            I => \N__23382\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__23440\,
            I => \N__23379\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__23435\,
            I => \N__23372\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__23420\,
            I => \N__23372\
        );

    \I__2983\ : Span4Mux_h
    port map (
            O => \N__23415\,
            I => \N__23372\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__23408\,
            I => \N__23367\
        );

    \I__2981\ : Span4Mux_v
    port map (
            O => \N__23401\,
            I => \N__23367\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__23394\,
            I => \N__23364\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__23385\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__2978\ : Odrv4
    port map (
            O => \N__23382\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__2977\ : Odrv4
    port map (
            O => \N__23379\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__2976\ : Odrv4
    port map (
            O => \N__23372\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__2975\ : Odrv4
    port map (
            O => \N__23367\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__2974\ : Odrv12
    port map (
            O => \N__23364\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__2973\ : CascadeMux
    port map (
            O => \N__23351\,
            I => \N__23346\
        );

    \I__2972\ : InMux
    port map (
            O => \N__23350\,
            I => \N__23342\
        );

    \I__2971\ : InMux
    port map (
            O => \N__23349\,
            I => \N__23339\
        );

    \I__2970\ : InMux
    port map (
            O => \N__23346\,
            I => \N__23336\
        );

    \I__2969\ : InMux
    port map (
            O => \N__23345\,
            I => \N__23333\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__23342\,
            I => \N__23330\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__23339\,
            I => \N__23327\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__23336\,
            I => \N__23324\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__23333\,
            I => \N__23321\
        );

    \I__2964\ : Span4Mux_v
    port map (
            O => \N__23330\,
            I => \N__23318\
        );

    \I__2963\ : Span4Mux_v
    port map (
            O => \N__23327\,
            I => \N__23315\
        );

    \I__2962\ : Span4Mux_v
    port map (
            O => \N__23324\,
            I => \N__23312\
        );

    \I__2961\ : Span12Mux_v
    port map (
            O => \N__23321\,
            I => \N__23309\
        );

    \I__2960\ : Odrv4
    port map (
            O => \N__23318\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__2959\ : Odrv4
    port map (
            O => \N__23315\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__2958\ : Odrv4
    port map (
            O => \N__23312\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__2957\ : Odrv12
    port map (
            O => \N__23309\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__2956\ : CascadeMux
    port map (
            O => \N__23300\,
            I => \N__23297\
        );

    \I__2955\ : InMux
    port map (
            O => \N__23297\,
            I => \N__23294\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__23294\,
            I => \N__23290\
        );

    \I__2953\ : InMux
    port map (
            O => \N__23293\,
            I => \N__23285\
        );

    \I__2952\ : Span4Mux_v
    port map (
            O => \N__23290\,
            I => \N__23282\
        );

    \I__2951\ : InMux
    port map (
            O => \N__23289\,
            I => \N__23279\
        );

    \I__2950\ : InMux
    port map (
            O => \N__23288\,
            I => \N__23276\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__23285\,
            I => \N__23273\
        );

    \I__2948\ : Odrv4
    port map (
            O => \N__23282\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__23279\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__23276\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__2945\ : Odrv4
    port map (
            O => \N__23273\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__2944\ : InMux
    port map (
            O => \N__23264\,
            I => \N__23260\
        );

    \I__2943\ : InMux
    port map (
            O => \N__23263\,
            I => \N__23257\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__23260\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__23257\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__2940\ : InMux
    port map (
            O => \N__23252\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\
        );

    \I__2939\ : InMux
    port map (
            O => \N__23249\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\
        );

    \I__2938\ : InMux
    port map (
            O => \N__23246\,
            I => \N__23243\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__23243\,
            I => \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2\
        );

    \I__2936\ : CascadeMux
    port map (
            O => \N__23240\,
            I => \N__23237\
        );

    \I__2935\ : InMux
    port map (
            O => \N__23237\,
            I => \N__23234\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__23234\,
            I => \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2\
        );

    \I__2933\ : InMux
    port map (
            O => \N__23231\,
            I => \N__23228\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__23228\,
            I => \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2\
        );

    \I__2931\ : CascadeMux
    port map (
            O => \N__23225\,
            I => \N__23222\
        );

    \I__2930\ : InMux
    port map (
            O => \N__23222\,
            I => \N__23219\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__23219\,
            I => \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2\
        );

    \I__2928\ : InMux
    port map (
            O => \N__23216\,
            I => \N__23213\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__23213\,
            I => \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23\
        );

    \I__2926\ : CascadeMux
    port map (
            O => \N__23210\,
            I => \N__23207\
        );

    \I__2925\ : InMux
    port map (
            O => \N__23207\,
            I => \N__23204\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__23204\,
            I => \N__23201\
        );

    \I__2923\ : Odrv4
    port map (
            O => \N__23201\,
            I => \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2\
        );

    \I__2922\ : InMux
    port map (
            O => \N__23198\,
            I => \N__23195\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__23195\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93\
        );

    \I__2920\ : InMux
    port map (
            O => \N__23192\,
            I => \N__23189\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__23189\,
            I => \N__23186\
        );

    \I__2918\ : Odrv12
    port map (
            O => \N__23186\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_22\
        );

    \I__2917\ : CascadeMux
    port map (
            O => \N__23183\,
            I => \N__23180\
        );

    \I__2916\ : InMux
    port map (
            O => \N__23180\,
            I => \N__23176\
        );

    \I__2915\ : CascadeMux
    port map (
            O => \N__23179\,
            I => \N__23172\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__23176\,
            I => \N__23169\
        );

    \I__2913\ : CascadeMux
    port map (
            O => \N__23175\,
            I => \N__23165\
        );

    \I__2912\ : InMux
    port map (
            O => \N__23172\,
            I => \N__23162\
        );

    \I__2911\ : Span4Mux_v
    port map (
            O => \N__23169\,
            I => \N__23159\
        );

    \I__2910\ : InMux
    port map (
            O => \N__23168\,
            I => \N__23156\
        );

    \I__2909\ : InMux
    port map (
            O => \N__23165\,
            I => \N__23153\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__23162\,
            I => \N__23150\
        );

    \I__2907\ : Odrv4
    port map (
            O => \N__23159\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__23156\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__23153\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__2904\ : Odrv4
    port map (
            O => \N__23150\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__2903\ : CascadeMux
    port map (
            O => \N__23141\,
            I => \N__23138\
        );

    \I__2902\ : InMux
    port map (
            O => \N__23138\,
            I => \N__23134\
        );

    \I__2901\ : InMux
    port map (
            O => \N__23137\,
            I => \N__23131\
        );

    \I__2900\ : LocalMux
    port map (
            O => \N__23134\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__23131\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__2898\ : InMux
    port map (
            O => \N__23126\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\
        );

    \I__2897\ : CascadeMux
    port map (
            O => \N__23123\,
            I => \N__23120\
        );

    \I__2896\ : InMux
    port map (
            O => \N__23120\,
            I => \N__23117\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__23117\,
            I => \N__23113\
        );

    \I__2894\ : InMux
    port map (
            O => \N__23116\,
            I => \N__23108\
        );

    \I__2893\ : Span4Mux_v
    port map (
            O => \N__23113\,
            I => \N__23105\
        );

    \I__2892\ : InMux
    port map (
            O => \N__23112\,
            I => \N__23102\
        );

    \I__2891\ : InMux
    port map (
            O => \N__23111\,
            I => \N__23099\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__23108\,
            I => \N__23096\
        );

    \I__2889\ : Odrv4
    port map (
            O => \N__23105\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__23102\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__23099\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__2886\ : Odrv12
    port map (
            O => \N__23096\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__2885\ : CascadeMux
    port map (
            O => \N__23087\,
            I => \N__23083\
        );

    \I__2884\ : InMux
    port map (
            O => \N__23086\,
            I => \N__23078\
        );

    \I__2883\ : InMux
    port map (
            O => \N__23083\,
            I => \N__23078\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__23078\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__2881\ : InMux
    port map (
            O => \N__23075\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\
        );

    \I__2880\ : CascadeMux
    port map (
            O => \N__23072\,
            I => \N__23069\
        );

    \I__2879\ : InMux
    port map (
            O => \N__23069\,
            I => \N__23066\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__23066\,
            I => \N__23061\
        );

    \I__2877\ : InMux
    port map (
            O => \N__23065\,
            I => \N__23057\
        );

    \I__2876\ : InMux
    port map (
            O => \N__23064\,
            I => \N__23054\
        );

    \I__2875\ : Span4Mux_v
    port map (
            O => \N__23061\,
            I => \N__23051\
        );

    \I__2874\ : InMux
    port map (
            O => \N__23060\,
            I => \N__23048\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__23057\,
            I => \N__23043\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__23054\,
            I => \N__23043\
        );

    \I__2871\ : Odrv4
    port map (
            O => \N__23051\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__23048\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__2869\ : Odrv12
    port map (
            O => \N__23043\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__2868\ : InMux
    port map (
            O => \N__23036\,
            I => \N__23030\
        );

    \I__2867\ : InMux
    port map (
            O => \N__23035\,
            I => \N__23030\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__23030\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__2865\ : InMux
    port map (
            O => \N__23027\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\
        );

    \I__2864\ : CascadeMux
    port map (
            O => \N__23024\,
            I => \N__23021\
        );

    \I__2863\ : InMux
    port map (
            O => \N__23021\,
            I => \N__23017\
        );

    \I__2862\ : CascadeMux
    port map (
            O => \N__23020\,
            I => \N__23014\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__23017\,
            I => \N__23011\
        );

    \I__2860\ : InMux
    port map (
            O => \N__23014\,
            I => \N__23006\
        );

    \I__2859\ : Span4Mux_v
    port map (
            O => \N__23011\,
            I => \N__23003\
        );

    \I__2858\ : InMux
    port map (
            O => \N__23010\,
            I => \N__23000\
        );

    \I__2857\ : InMux
    port map (
            O => \N__23009\,
            I => \N__22997\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__23006\,
            I => \N__22994\
        );

    \I__2855\ : Odrv4
    port map (
            O => \N__23003\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__23000\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__22997\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__2852\ : Odrv4
    port map (
            O => \N__22994\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__2851\ : InMux
    port map (
            O => \N__22985\,
            I => \N__22979\
        );

    \I__2850\ : InMux
    port map (
            O => \N__22984\,
            I => \N__22979\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__22979\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__2848\ : InMux
    port map (
            O => \N__22976\,
            I => \bfn_4_20_0_\
        );

    \I__2847\ : CascadeMux
    port map (
            O => \N__22973\,
            I => \N__22970\
        );

    \I__2846\ : InMux
    port map (
            O => \N__22970\,
            I => \N__22966\
        );

    \I__2845\ : InMux
    port map (
            O => \N__22969\,
            I => \N__22963\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__22966\,
            I => \N__22959\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__22963\,
            I => \N__22956\
        );

    \I__2842\ : InMux
    port map (
            O => \N__22962\,
            I => \N__22952\
        );

    \I__2841\ : Span4Mux_h
    port map (
            O => \N__22959\,
            I => \N__22947\
        );

    \I__2840\ : Span4Mux_h
    port map (
            O => \N__22956\,
            I => \N__22947\
        );

    \I__2839\ : InMux
    port map (
            O => \N__22955\,
            I => \N__22944\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__22952\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__2837\ : Odrv4
    port map (
            O => \N__22947\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__22944\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__2835\ : InMux
    port map (
            O => \N__22937\,
            I => \N__22931\
        );

    \I__2834\ : InMux
    port map (
            O => \N__22936\,
            I => \N__22931\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__22931\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__2832\ : InMux
    port map (
            O => \N__22928\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\
        );

    \I__2831\ : CascadeMux
    port map (
            O => \N__22925\,
            I => \N__22921\
        );

    \I__2830\ : InMux
    port map (
            O => \N__22924\,
            I => \N__22918\
        );

    \I__2829\ : InMux
    port map (
            O => \N__22921\,
            I => \N__22915\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__22918\,
            I => \N__22912\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__22915\,
            I => \N__22908\
        );

    \I__2826\ : Span4Mux_h
    port map (
            O => \N__22912\,
            I => \N__22904\
        );

    \I__2825\ : InMux
    port map (
            O => \N__22911\,
            I => \N__22901\
        );

    \I__2824\ : Span4Mux_h
    port map (
            O => \N__22908\,
            I => \N__22898\
        );

    \I__2823\ : InMux
    port map (
            O => \N__22907\,
            I => \N__22895\
        );

    \I__2822\ : Odrv4
    port map (
            O => \N__22904\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__22901\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__2820\ : Odrv4
    port map (
            O => \N__22898\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__22895\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__2818\ : InMux
    port map (
            O => \N__22886\,
            I => \N__22882\
        );

    \I__2817\ : InMux
    port map (
            O => \N__22885\,
            I => \N__22879\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__22882\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__22879\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__2814\ : InMux
    port map (
            O => \N__22874\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\
        );

    \I__2813\ : InMux
    port map (
            O => \N__22871\,
            I => \N__22868\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__22868\,
            I => \N__22864\
        );

    \I__2811\ : InMux
    port map (
            O => \N__22867\,
            I => \N__22859\
        );

    \I__2810\ : Span4Mux_v
    port map (
            O => \N__22864\,
            I => \N__22856\
        );

    \I__2809\ : InMux
    port map (
            O => \N__22863\,
            I => \N__22853\
        );

    \I__2808\ : InMux
    port map (
            O => \N__22862\,
            I => \N__22850\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__22859\,
            I => \N__22847\
        );

    \I__2806\ : Odrv4
    port map (
            O => \N__22856\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__22853\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__22850\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__2803\ : Odrv4
    port map (
            O => \N__22847\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__2802\ : InMux
    port map (
            O => \N__22838\,
            I => \N__22832\
        );

    \I__2801\ : InMux
    port map (
            O => \N__22837\,
            I => \N__22832\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__22832\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__2799\ : InMux
    port map (
            O => \N__22829\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\
        );

    \I__2798\ : InMux
    port map (
            O => \N__22826\,
            I => \N__22823\
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__22823\,
            I => \N__22820\
        );

    \I__2796\ : Span4Mux_v
    port map (
            O => \N__22820\,
            I => \N__22814\
        );

    \I__2795\ : InMux
    port map (
            O => \N__22819\,
            I => \N__22811\
        );

    \I__2794\ : InMux
    port map (
            O => \N__22818\,
            I => \N__22808\
        );

    \I__2793\ : InMux
    port map (
            O => \N__22817\,
            I => \N__22805\
        );

    \I__2792\ : Odrv4
    port map (
            O => \N__22814\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__22811\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__22808\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__22805\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__2788\ : CascadeMux
    port map (
            O => \N__22796\,
            I => \N__22792\
        );

    \I__2787\ : CascadeMux
    port map (
            O => \N__22795\,
            I => \N__22789\
        );

    \I__2786\ : InMux
    port map (
            O => \N__22792\,
            I => \N__22786\
        );

    \I__2785\ : InMux
    port map (
            O => \N__22789\,
            I => \N__22783\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__22786\,
            I => \N__22780\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__22783\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__2782\ : Odrv4
    port map (
            O => \N__22780\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__2781\ : InMux
    port map (
            O => \N__22775\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\
        );

    \I__2780\ : CascadeMux
    port map (
            O => \N__22772\,
            I => \N__22769\
        );

    \I__2779\ : InMux
    port map (
            O => \N__22769\,
            I => \N__22766\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__22766\,
            I => \N__22761\
        );

    \I__2777\ : InMux
    port map (
            O => \N__22765\,
            I => \N__22757\
        );

    \I__2776\ : InMux
    port map (
            O => \N__22764\,
            I => \N__22754\
        );

    \I__2775\ : Span4Mux_v
    port map (
            O => \N__22761\,
            I => \N__22751\
        );

    \I__2774\ : InMux
    port map (
            O => \N__22760\,
            I => \N__22748\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__22757\,
            I => \N__22743\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__22754\,
            I => \N__22743\
        );

    \I__2771\ : Odrv4
    port map (
            O => \N__22751\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__22748\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__2769\ : Odrv4
    port map (
            O => \N__22743\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__2768\ : CascadeMux
    port map (
            O => \N__22736\,
            I => \N__22733\
        );

    \I__2767\ : InMux
    port map (
            O => \N__22733\,
            I => \N__22730\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__22730\,
            I => \N__22727\
        );

    \I__2765\ : Span4Mux_v
    port map (
            O => \N__22727\,
            I => \N__22723\
        );

    \I__2764\ : InMux
    port map (
            O => \N__22726\,
            I => \N__22720\
        );

    \I__2763\ : Odrv4
    port map (
            O => \N__22723\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__22720\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__2761\ : InMux
    port map (
            O => \N__22715\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\
        );

    \I__2760\ : CascadeMux
    port map (
            O => \N__22712\,
            I => \N__22709\
        );

    \I__2759\ : InMux
    port map (
            O => \N__22709\,
            I => \N__22706\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__22706\,
            I => \N__22701\
        );

    \I__2757\ : InMux
    port map (
            O => \N__22705\,
            I => \N__22698\
        );

    \I__2756\ : InMux
    port map (
            O => \N__22704\,
            I => \N__22695\
        );

    \I__2755\ : Span4Mux_v
    port map (
            O => \N__22701\,
            I => \N__22691\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__22698\,
            I => \N__22686\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__22695\,
            I => \N__22686\
        );

    \I__2752\ : InMux
    port map (
            O => \N__22694\,
            I => \N__22683\
        );

    \I__2751\ : Odrv4
    port map (
            O => \N__22691\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__2750\ : Odrv4
    port map (
            O => \N__22686\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__22683\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__2748\ : InMux
    port map (
            O => \N__22676\,
            I => \N__22670\
        );

    \I__2747\ : InMux
    port map (
            O => \N__22675\,
            I => \N__22670\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__22670\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__2745\ : InMux
    port map (
            O => \N__22667\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\
        );

    \I__2744\ : CascadeMux
    port map (
            O => \N__22664\,
            I => \N__22661\
        );

    \I__2743\ : InMux
    port map (
            O => \N__22661\,
            I => \N__22657\
        );

    \I__2742\ : InMux
    port map (
            O => \N__22660\,
            I => \N__22652\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__22657\,
            I => \N__22649\
        );

    \I__2740\ : InMux
    port map (
            O => \N__22656\,
            I => \N__22646\
        );

    \I__2739\ : InMux
    port map (
            O => \N__22655\,
            I => \N__22643\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__22652\,
            I => \N__22640\
        );

    \I__2737\ : Span4Mux_h
    port map (
            O => \N__22649\,
            I => \N__22631\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__22646\,
            I => \N__22631\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__22643\,
            I => \N__22631\
        );

    \I__2734\ : Span4Mux_s3_h
    port map (
            O => \N__22640\,
            I => \N__22631\
        );

    \I__2733\ : Odrv4
    port map (
            O => \N__22631\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__2732\ : InMux
    port map (
            O => \N__22628\,
            I => \N__22622\
        );

    \I__2731\ : InMux
    port map (
            O => \N__22627\,
            I => \N__22622\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__22622\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__2729\ : InMux
    port map (
            O => \N__22619\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\
        );

    \I__2728\ : CascadeMux
    port map (
            O => \N__22616\,
            I => \N__22613\
        );

    \I__2727\ : InMux
    port map (
            O => \N__22613\,
            I => \N__22609\
        );

    \I__2726\ : InMux
    port map (
            O => \N__22612\,
            I => \N__22605\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__22609\,
            I => \N__22601\
        );

    \I__2724\ : InMux
    port map (
            O => \N__22608\,
            I => \N__22598\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__22605\,
            I => \N__22595\
        );

    \I__2722\ : InMux
    port map (
            O => \N__22604\,
            I => \N__22592\
        );

    \I__2721\ : Span4Mux_v
    port map (
            O => \N__22601\,
            I => \N__22587\
        );

    \I__2720\ : LocalMux
    port map (
            O => \N__22598\,
            I => \N__22587\
        );

    \I__2719\ : Span4Mux_h
    port map (
            O => \N__22595\,
            I => \N__22584\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__22592\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__2717\ : Odrv4
    port map (
            O => \N__22587\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__2716\ : Odrv4
    port map (
            O => \N__22584\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__2715\ : InMux
    port map (
            O => \N__22577\,
            I => \N__22573\
        );

    \I__2714\ : InMux
    port map (
            O => \N__22576\,
            I => \N__22570\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__22573\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__22570\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__2711\ : InMux
    port map (
            O => \N__22565\,
            I => \bfn_4_19_0_\
        );

    \I__2710\ : InMux
    port map (
            O => \N__22562\,
            I => \N__22559\
        );

    \I__2709\ : LocalMux
    port map (
            O => \N__22559\,
            I => \N__22556\
        );

    \I__2708\ : Odrv4
    port map (
            O => \N__22556\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_18\
        );

    \I__2707\ : CascadeMux
    port map (
            O => \N__22553\,
            I => \N__22550\
        );

    \I__2706\ : InMux
    port map (
            O => \N__22550\,
            I => \N__22547\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__22547\,
            I => \N__22543\
        );

    \I__2704\ : InMux
    port map (
            O => \N__22546\,
            I => \N__22538\
        );

    \I__2703\ : Span4Mux_v
    port map (
            O => \N__22543\,
            I => \N__22535\
        );

    \I__2702\ : InMux
    port map (
            O => \N__22542\,
            I => \N__22532\
        );

    \I__2701\ : InMux
    port map (
            O => \N__22541\,
            I => \N__22529\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__22538\,
            I => \N__22526\
        );

    \I__2699\ : Odrv4
    port map (
            O => \N__22535\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__22532\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__22529\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__2696\ : Odrv4
    port map (
            O => \N__22526\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__2695\ : CascadeMux
    port map (
            O => \N__22517\,
            I => \N__22514\
        );

    \I__2694\ : InMux
    port map (
            O => \N__22514\,
            I => \N__22510\
        );

    \I__2693\ : InMux
    port map (
            O => \N__22513\,
            I => \N__22507\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__22510\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__22507\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__2690\ : InMux
    port map (
            O => \N__22502\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\
        );

    \I__2689\ : InMux
    port map (
            O => \N__22499\,
            I => \N__22496\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__22496\,
            I => \N__22491\
        );

    \I__2687\ : CascadeMux
    port map (
            O => \N__22495\,
            I => \N__22488\
        );

    \I__2686\ : InMux
    port map (
            O => \N__22494\,
            I => \N__22484\
        );

    \I__2685\ : Span4Mux_v
    port map (
            O => \N__22491\,
            I => \N__22481\
        );

    \I__2684\ : InMux
    port map (
            O => \N__22488\,
            I => \N__22478\
        );

    \I__2683\ : InMux
    port map (
            O => \N__22487\,
            I => \N__22475\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__22484\,
            I => \N__22472\
        );

    \I__2681\ : Odrv4
    port map (
            O => \N__22481\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__22478\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__22475\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__2678\ : Odrv4
    port map (
            O => \N__22472\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__2677\ : InMux
    port map (
            O => \N__22463\,
            I => \N__22457\
        );

    \I__2676\ : InMux
    port map (
            O => \N__22462\,
            I => \N__22457\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__22457\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__2674\ : InMux
    port map (
            O => \N__22454\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\
        );

    \I__2673\ : InMux
    port map (
            O => \N__22451\,
            I => \N__22448\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__22448\,
            I => \N__22445\
        );

    \I__2671\ : Odrv12
    port map (
            O => \N__22445\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_20\
        );

    \I__2670\ : CascadeMux
    port map (
            O => \N__22442\,
            I => \N__22439\
        );

    \I__2669\ : InMux
    port map (
            O => \N__22439\,
            I => \N__22436\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__22436\,
            I => \N__22432\
        );

    \I__2667\ : CascadeMux
    port map (
            O => \N__22435\,
            I => \N__22427\
        );

    \I__2666\ : Span4Mux_h
    port map (
            O => \N__22432\,
            I => \N__22424\
        );

    \I__2665\ : InMux
    port map (
            O => \N__22431\,
            I => \N__22421\
        );

    \I__2664\ : InMux
    port map (
            O => \N__22430\,
            I => \N__22418\
        );

    \I__2663\ : InMux
    port map (
            O => \N__22427\,
            I => \N__22415\
        );

    \I__2662\ : Sp12to4
    port map (
            O => \N__22424\,
            I => \N__22408\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__22421\,
            I => \N__22408\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__22418\,
            I => \N__22408\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__22415\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__2658\ : Odrv12
    port map (
            O => \N__22408\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__2657\ : CascadeMux
    port map (
            O => \N__22403\,
            I => \N__22399\
        );

    \I__2656\ : InMux
    port map (
            O => \N__22402\,
            I => \N__22394\
        );

    \I__2655\ : InMux
    port map (
            O => \N__22399\,
            I => \N__22394\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__22394\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__2653\ : InMux
    port map (
            O => \N__22391\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\
        );

    \I__2652\ : CascadeMux
    port map (
            O => \N__22388\,
            I => \N__22385\
        );

    \I__2651\ : InMux
    port map (
            O => \N__22385\,
            I => \N__22381\
        );

    \I__2650\ : CascadeMux
    port map (
            O => \N__22384\,
            I => \N__22378\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__22381\,
            I => \N__22375\
        );

    \I__2648\ : InMux
    port map (
            O => \N__22378\,
            I => \N__22372\
        );

    \I__2647\ : Span4Mux_h
    port map (
            O => \N__22375\,
            I => \N__22368\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__22372\,
            I => \N__22364\
        );

    \I__2645\ : InMux
    port map (
            O => \N__22371\,
            I => \N__22361\
        );

    \I__2644\ : Span4Mux_v
    port map (
            O => \N__22368\,
            I => \N__22358\
        );

    \I__2643\ : InMux
    port map (
            O => \N__22367\,
            I => \N__22355\
        );

    \I__2642\ : Span4Mux_v
    port map (
            O => \N__22364\,
            I => \N__22350\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__22361\,
            I => \N__22350\
        );

    \I__2640\ : Odrv4
    port map (
            O => \N__22358\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__22355\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__2638\ : Odrv4
    port map (
            O => \N__22350\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__2637\ : InMux
    port map (
            O => \N__22343\,
            I => \N__22340\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__22340\,
            I => \N__22336\
        );

    \I__2635\ : InMux
    port map (
            O => \N__22339\,
            I => \N__22333\
        );

    \I__2634\ : Odrv4
    port map (
            O => \N__22336\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__22333\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__2632\ : InMux
    port map (
            O => \N__22328\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\
        );

    \I__2631\ : InMux
    port map (
            O => \N__22325\,
            I => \N__22322\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__22322\,
            I => \N__22319\
        );

    \I__2629\ : Odrv12
    port map (
            O => \N__22319\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\
        );

    \I__2628\ : CascadeMux
    port map (
            O => \N__22316\,
            I => \N__22313\
        );

    \I__2627\ : InMux
    port map (
            O => \N__22313\,
            I => \N__22310\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__22310\,
            I => \N__22305\
        );

    \I__2625\ : InMux
    port map (
            O => \N__22309\,
            I => \N__22302\
        );

    \I__2624\ : InMux
    port map (
            O => \N__22308\,
            I => \N__22299\
        );

    \I__2623\ : Span4Mux_v
    port map (
            O => \N__22305\,
            I => \N__22294\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__22302\,
            I => \N__22294\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__22299\,
            I => \N__22291\
        );

    \I__2620\ : Span4Mux_h
    port map (
            O => \N__22294\,
            I => \N__22288\
        );

    \I__2619\ : Span4Mux_v
    port map (
            O => \N__22291\,
            I => \N__22285\
        );

    \I__2618\ : Odrv4
    port map (
            O => \N__22288\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2617\ : Odrv4
    port map (
            O => \N__22285\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2616\ : InMux
    port map (
            O => \N__22280\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\
        );

    \I__2615\ : InMux
    port map (
            O => \N__22277\,
            I => \N__22273\
        );

    \I__2614\ : InMux
    port map (
            O => \N__22276\,
            I => \N__22270\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__22273\,
            I => \N__22266\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__22270\,
            I => \N__22263\
        );

    \I__2611\ : InMux
    port map (
            O => \N__22269\,
            I => \N__22260\
        );

    \I__2610\ : Span4Mux_v
    port map (
            O => \N__22266\,
            I => \N__22257\
        );

    \I__2609\ : Span4Mux_v
    port map (
            O => \N__22263\,
            I => \N__22251\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__22260\,
            I => \N__22251\
        );

    \I__2607\ : Span4Mux_h
    port map (
            O => \N__22257\,
            I => \N__22248\
        );

    \I__2606\ : InMux
    port map (
            O => \N__22256\,
            I => \N__22245\
        );

    \I__2605\ : Odrv4
    port map (
            O => \N__22251\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__2604\ : Odrv4
    port map (
            O => \N__22248\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__22245\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__2602\ : CascadeMux
    port map (
            O => \N__22238\,
            I => \N__22235\
        );

    \I__2601\ : InMux
    port map (
            O => \N__22235\,
            I => \N__22230\
        );

    \I__2600\ : InMux
    port map (
            O => \N__22234\,
            I => \N__22227\
        );

    \I__2599\ : InMux
    port map (
            O => \N__22233\,
            I => \N__22224\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__22230\,
            I => \N__22221\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__22227\,
            I => \N__22218\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__22224\,
            I => \N__22215\
        );

    \I__2595\ : Span12Mux_v
    port map (
            O => \N__22221\,
            I => \N__22212\
        );

    \I__2594\ : Span4Mux_h
    port map (
            O => \N__22218\,
            I => \N__22209\
        );

    \I__2593\ : Span4Mux_v
    port map (
            O => \N__22215\,
            I => \N__22206\
        );

    \I__2592\ : Odrv12
    port map (
            O => \N__22212\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2591\ : Odrv4
    port map (
            O => \N__22209\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2590\ : Odrv4
    port map (
            O => \N__22206\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2589\ : InMux
    port map (
            O => \N__22199\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\
        );

    \I__2588\ : InMux
    port map (
            O => \N__22196\,
            I => \N__22191\
        );

    \I__2587\ : CascadeMux
    port map (
            O => \N__22195\,
            I => \N__22187\
        );

    \I__2586\ : InMux
    port map (
            O => \N__22194\,
            I => \N__22184\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__22191\,
            I => \N__22181\
        );

    \I__2584\ : CascadeMux
    port map (
            O => \N__22190\,
            I => \N__22178\
        );

    \I__2583\ : InMux
    port map (
            O => \N__22187\,
            I => \N__22175\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__22184\,
            I => \N__22172\
        );

    \I__2581\ : Span4Mux_v
    port map (
            O => \N__22181\,
            I => \N__22169\
        );

    \I__2580\ : InMux
    port map (
            O => \N__22178\,
            I => \N__22166\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__22175\,
            I => \N__22161\
        );

    \I__2578\ : Span4Mux_h
    port map (
            O => \N__22172\,
            I => \N__22161\
        );

    \I__2577\ : Odrv4
    port map (
            O => \N__22169\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__22166\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__2575\ : Odrv4
    port map (
            O => \N__22161\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__2574\ : InMux
    port map (
            O => \N__22154\,
            I => \N__22150\
        );

    \I__2573\ : InMux
    port map (
            O => \N__22153\,
            I => \N__22146\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__22150\,
            I => \N__22143\
        );

    \I__2571\ : InMux
    port map (
            O => \N__22149\,
            I => \N__22140\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__22146\,
            I => \N__22137\
        );

    \I__2569\ : Span4Mux_s3_h
    port map (
            O => \N__22143\,
            I => \N__22132\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__22140\,
            I => \N__22132\
        );

    \I__2567\ : Span4Mux_h
    port map (
            O => \N__22137\,
            I => \N__22129\
        );

    \I__2566\ : Span4Mux_v
    port map (
            O => \N__22132\,
            I => \N__22126\
        );

    \I__2565\ : Odrv4
    port map (
            O => \N__22129\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2564\ : Odrv4
    port map (
            O => \N__22126\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2563\ : InMux
    port map (
            O => \N__22121\,
            I => \bfn_4_18_0_\
        );

    \I__2562\ : InMux
    port map (
            O => \N__22118\,
            I => \N__22115\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__22115\,
            I => \N__22112\
        );

    \I__2560\ : Odrv12
    port map (
            O => \N__22112\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\
        );

    \I__2559\ : CascadeMux
    port map (
            O => \N__22109\,
            I => \N__22106\
        );

    \I__2558\ : InMux
    port map (
            O => \N__22106\,
            I => \N__22101\
        );

    \I__2557\ : CascadeMux
    port map (
            O => \N__22105\,
            I => \N__22098\
        );

    \I__2556\ : CascadeMux
    port map (
            O => \N__22104\,
            I => \N__22095\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__22101\,
            I => \N__22092\
        );

    \I__2554\ : InMux
    port map (
            O => \N__22098\,
            I => \N__22089\
        );

    \I__2553\ : InMux
    port map (
            O => \N__22095\,
            I => \N__22086\
        );

    \I__2552\ : Span4Mux_h
    port map (
            O => \N__22092\,
            I => \N__22081\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__22089\,
            I => \N__22081\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__22086\,
            I => \N__22078\
        );

    \I__2549\ : Span4Mux_v
    port map (
            O => \N__22081\,
            I => \N__22074\
        );

    \I__2548\ : Span12Mux_v
    port map (
            O => \N__22078\,
            I => \N__22071\
        );

    \I__2547\ : InMux
    port map (
            O => \N__22077\,
            I => \N__22068\
        );

    \I__2546\ : Odrv4
    port map (
            O => \N__22074\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__2545\ : Odrv12
    port map (
            O => \N__22071\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__22068\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__2543\ : InMux
    port map (
            O => \N__22061\,
            I => \N__22055\
        );

    \I__2542\ : InMux
    port map (
            O => \N__22060\,
            I => \N__22055\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__22055\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__2540\ : InMux
    port map (
            O => \N__22052\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\
        );

    \I__2539\ : InMux
    port map (
            O => \N__22049\,
            I => \N__22046\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__22046\,
            I => \N__22043\
        );

    \I__2537\ : Odrv12
    port map (
            O => \N__22043\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\
        );

    \I__2536\ : CascadeMux
    port map (
            O => \N__22040\,
            I => \N__22036\
        );

    \I__2535\ : CascadeMux
    port map (
            O => \N__22039\,
            I => \N__22033\
        );

    \I__2534\ : InMux
    port map (
            O => \N__22036\,
            I => \N__22029\
        );

    \I__2533\ : InMux
    port map (
            O => \N__22033\,
            I => \N__22026\
        );

    \I__2532\ : InMux
    port map (
            O => \N__22032\,
            I => \N__22023\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__22029\,
            I => \N__22019\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__22026\,
            I => \N__22016\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__22023\,
            I => \N__22013\
        );

    \I__2528\ : InMux
    port map (
            O => \N__22022\,
            I => \N__22010\
        );

    \I__2527\ : Span4Mux_v
    port map (
            O => \N__22019\,
            I => \N__22007\
        );

    \I__2526\ : Span4Mux_v
    port map (
            O => \N__22016\,
            I => \N__22002\
        );

    \I__2525\ : Span4Mux_s3_h
    port map (
            O => \N__22013\,
            I => \N__22002\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__22010\,
            I => \N__21999\
        );

    \I__2523\ : Odrv4
    port map (
            O => \N__22007\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__2522\ : Odrv4
    port map (
            O => \N__22002\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__2521\ : Odrv12
    port map (
            O => \N__21999\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__2520\ : InMux
    port map (
            O => \N__21992\,
            I => \N__21986\
        );

    \I__2519\ : InMux
    port map (
            O => \N__21991\,
            I => \N__21986\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__21986\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__2517\ : InMux
    port map (
            O => \N__21983\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\
        );

    \I__2516\ : InMux
    port map (
            O => \N__21980\,
            I => \N__21974\
        );

    \I__2515\ : InMux
    port map (
            O => \N__21979\,
            I => \N__21971\
        );

    \I__2514\ : InMux
    port map (
            O => \N__21978\,
            I => \N__21968\
        );

    \I__2513\ : InMux
    port map (
            O => \N__21977\,
            I => \N__21965\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__21974\,
            I => \N__21962\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__21971\,
            I => \N__21959\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__21968\,
            I => \N__21952\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__21965\,
            I => \N__21952\
        );

    \I__2508\ : Span4Mux_s3_h
    port map (
            O => \N__21962\,
            I => \N__21952\
        );

    \I__2507\ : Odrv4
    port map (
            O => \N__21959\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__2506\ : Odrv4
    port map (
            O => \N__21952\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__2505\ : InMux
    port map (
            O => \N__21947\,
            I => \N__21943\
        );

    \I__2504\ : InMux
    port map (
            O => \N__21946\,
            I => \N__21940\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__21943\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__21940\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__2501\ : InMux
    port map (
            O => \N__21935\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\
        );

    \I__2500\ : InMux
    port map (
            O => \N__21932\,
            I => \N__21929\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__21929\,
            I => \N__21926\
        );

    \I__2498\ : Odrv4
    port map (
            O => \N__21926\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\
        );

    \I__2497\ : CascadeMux
    port map (
            O => \N__21923\,
            I => \N__21920\
        );

    \I__2496\ : InMux
    port map (
            O => \N__21920\,
            I => \N__21915\
        );

    \I__2495\ : InMux
    port map (
            O => \N__21919\,
            I => \N__21912\
        );

    \I__2494\ : InMux
    port map (
            O => \N__21918\,
            I => \N__21908\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__21915\,
            I => \N__21905\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__21912\,
            I => \N__21902\
        );

    \I__2491\ : InMux
    port map (
            O => \N__21911\,
            I => \N__21899\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__21908\,
            I => \N__21896\
        );

    \I__2489\ : Span4Mux_v
    port map (
            O => \N__21905\,
            I => \N__21893\
        );

    \I__2488\ : Sp12to4
    port map (
            O => \N__21902\,
            I => \N__21888\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__21899\,
            I => \N__21888\
        );

    \I__2486\ : Span4Mux_s3_h
    port map (
            O => \N__21896\,
            I => \N__21885\
        );

    \I__2485\ : Odrv4
    port map (
            O => \N__21893\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__2484\ : Odrv12
    port map (
            O => \N__21888\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__2483\ : Odrv4
    port map (
            O => \N__21885\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__2482\ : InMux
    port map (
            O => \N__21878\,
            I => \N__21875\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__21875\,
            I => \N__21871\
        );

    \I__2480\ : InMux
    port map (
            O => \N__21874\,
            I => \N__21868\
        );

    \I__2479\ : Odrv4
    port map (
            O => \N__21871\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__21868\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__2477\ : InMux
    port map (
            O => \N__21863\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\
        );

    \I__2476\ : CascadeMux
    port map (
            O => \N__21860\,
            I => \N__21857\
        );

    \I__2475\ : InMux
    port map (
            O => \N__21857\,
            I => \N__21852\
        );

    \I__2474\ : InMux
    port map (
            O => \N__21856\,
            I => \N__21849\
        );

    \I__2473\ : InMux
    port map (
            O => \N__21855\,
            I => \N__21844\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__21852\,
            I => \N__21841\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__21849\,
            I => \N__21838\
        );

    \I__2470\ : InMux
    port map (
            O => \N__21848\,
            I => \N__21835\
        );

    \I__2469\ : InMux
    port map (
            O => \N__21847\,
            I => \N__21832\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__21844\,
            I => \N__21829\
        );

    \I__2467\ : Span4Mux_v
    port map (
            O => \N__21841\,
            I => \N__21826\
        );

    \I__2466\ : Span4Mux_v
    port map (
            O => \N__21838\,
            I => \N__21823\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__21835\,
            I => \N__21820\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__21832\,
            I => \N__21811\
        );

    \I__2463\ : Span4Mux_v
    port map (
            O => \N__21829\,
            I => \N__21811\
        );

    \I__2462\ : Span4Mux_h
    port map (
            O => \N__21826\,
            I => \N__21811\
        );

    \I__2461\ : Span4Mux_s1_h
    port map (
            O => \N__21823\,
            I => \N__21811\
        );

    \I__2460\ : Odrv12
    port map (
            O => \N__21820\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__2459\ : Odrv4
    port map (
            O => \N__21811\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__2458\ : InMux
    port map (
            O => \N__21806\,
            I => \N__21803\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__21803\,
            I => \N__21800\
        );

    \I__2456\ : Odrv4
    port map (
            O => \N__21800\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\
        );

    \I__2455\ : CascadeMux
    port map (
            O => \N__21797\,
            I => \N__21794\
        );

    \I__2454\ : InMux
    port map (
            O => \N__21794\,
            I => \N__21790\
        );

    \I__2453\ : InMux
    port map (
            O => \N__21793\,
            I => \N__21786\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__21790\,
            I => \N__21783\
        );

    \I__2451\ : InMux
    port map (
            O => \N__21789\,
            I => \N__21780\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__21786\,
            I => \N__21777\
        );

    \I__2449\ : Span4Mux_v
    port map (
            O => \N__21783\,
            I => \N__21774\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__21780\,
            I => \N__21771\
        );

    \I__2447\ : Odrv12
    port map (
            O => \N__21777\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__2446\ : Odrv4
    port map (
            O => \N__21774\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__2445\ : Odrv12
    port map (
            O => \N__21771\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__2444\ : InMux
    port map (
            O => \N__21764\,
            I => \N__21761\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__21761\,
            I => \N__21758\
        );

    \I__2442\ : Span4Mux_h
    port map (
            O => \N__21758\,
            I => \N__21755\
        );

    \I__2441\ : Span4Mux_v
    port map (
            O => \N__21755\,
            I => \N__21752\
        );

    \I__2440\ : Odrv4
    port map (
            O => \N__21752\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\
        );

    \I__2439\ : InMux
    port map (
            O => \N__21749\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\
        );

    \I__2438\ : InMux
    port map (
            O => \N__21746\,
            I => \N__21743\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__21743\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\
        );

    \I__2436\ : CascadeMux
    port map (
            O => \N__21740\,
            I => \N__21736\
        );

    \I__2435\ : InMux
    port map (
            O => \N__21739\,
            I => \N__21732\
        );

    \I__2434\ : InMux
    port map (
            O => \N__21736\,
            I => \N__21729\
        );

    \I__2433\ : InMux
    port map (
            O => \N__21735\,
            I => \N__21726\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__21732\,
            I => \N__21721\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__21729\,
            I => \N__21721\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__21726\,
            I => \N__21717\
        );

    \I__2429\ : Span4Mux_h
    port map (
            O => \N__21721\,
            I => \N__21714\
        );

    \I__2428\ : CascadeMux
    port map (
            O => \N__21720\,
            I => \N__21711\
        );

    \I__2427\ : Span4Mux_v
    port map (
            O => \N__21717\,
            I => \N__21708\
        );

    \I__2426\ : Span4Mux_v
    port map (
            O => \N__21714\,
            I => \N__21705\
        );

    \I__2425\ : InMux
    port map (
            O => \N__21711\,
            I => \N__21702\
        );

    \I__2424\ : Odrv4
    port map (
            O => \N__21708\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__2423\ : Odrv4
    port map (
            O => \N__21705\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__21702\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__2421\ : InMux
    port map (
            O => \N__21695\,
            I => \N__21692\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__21692\,
            I => \N__21687\
        );

    \I__2419\ : InMux
    port map (
            O => \N__21691\,
            I => \N__21684\
        );

    \I__2418\ : InMux
    port map (
            O => \N__21690\,
            I => \N__21681\
        );

    \I__2417\ : Span4Mux_v
    port map (
            O => \N__21687\,
            I => \N__21674\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__21684\,
            I => \N__21674\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__21681\,
            I => \N__21674\
        );

    \I__2414\ : Span4Mux_v
    port map (
            O => \N__21674\,
            I => \N__21671\
        );

    \I__2413\ : Odrv4
    port map (
            O => \N__21671\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__2412\ : InMux
    port map (
            O => \N__21668\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\
        );

    \I__2411\ : InMux
    port map (
            O => \N__21665\,
            I => \N__21662\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__21662\,
            I => \N__21659\
        );

    \I__2409\ : Odrv4
    port map (
            O => \N__21659\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\
        );

    \I__2408\ : CascadeMux
    port map (
            O => \N__21656\,
            I => \N__21651\
        );

    \I__2407\ : CascadeMux
    port map (
            O => \N__21655\,
            I => \N__21648\
        );

    \I__2406\ : InMux
    port map (
            O => \N__21654\,
            I => \N__21645\
        );

    \I__2405\ : InMux
    port map (
            O => \N__21651\,
            I => \N__21642\
        );

    \I__2404\ : InMux
    port map (
            O => \N__21648\,
            I => \N__21639\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__21645\,
            I => \N__21633\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__21642\,
            I => \N__21633\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__21639\,
            I => \N__21630\
        );

    \I__2400\ : InMux
    port map (
            O => \N__21638\,
            I => \N__21627\
        );

    \I__2399\ : Span4Mux_v
    port map (
            O => \N__21633\,
            I => \N__21624\
        );

    \I__2398\ : Span4Mux_v
    port map (
            O => \N__21630\,
            I => \N__21621\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__21627\,
            I => \N__21618\
        );

    \I__2396\ : Odrv4
    port map (
            O => \N__21624\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__2395\ : Odrv4
    port map (
            O => \N__21621\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__2394\ : Odrv12
    port map (
            O => \N__21618\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__2393\ : InMux
    port map (
            O => \N__21611\,
            I => \N__21608\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__21608\,
            I => \N__21602\
        );

    \I__2391\ : InMux
    port map (
            O => \N__21607\,
            I => \N__21599\
        );

    \I__2390\ : InMux
    port map (
            O => \N__21606\,
            I => \N__21594\
        );

    \I__2389\ : InMux
    port map (
            O => \N__21605\,
            I => \N__21594\
        );

    \I__2388\ : Span4Mux_v
    port map (
            O => \N__21602\,
            I => \N__21587\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__21599\,
            I => \N__21587\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__21594\,
            I => \N__21587\
        );

    \I__2385\ : Span4Mux_v
    port map (
            O => \N__21587\,
            I => \N__21584\
        );

    \I__2384\ : Odrv4
    port map (
            O => \N__21584\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2383\ : InMux
    port map (
            O => \N__21581\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\
        );

    \I__2382\ : InMux
    port map (
            O => \N__21578\,
            I => \N__21573\
        );

    \I__2381\ : InMux
    port map (
            O => \N__21577\,
            I => \N__21569\
        );

    \I__2380\ : InMux
    port map (
            O => \N__21576\,
            I => \N__21566\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__21573\,
            I => \N__21563\
        );

    \I__2378\ : InMux
    port map (
            O => \N__21572\,
            I => \N__21560\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__21569\,
            I => \N__21557\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__21566\,
            I => \N__21554\
        );

    \I__2375\ : Span4Mux_v
    port map (
            O => \N__21563\,
            I => \N__21551\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__21560\,
            I => \N__21544\
        );

    \I__2373\ : Span4Mux_h
    port map (
            O => \N__21557\,
            I => \N__21544\
        );

    \I__2372\ : Span4Mux_s3_h
    port map (
            O => \N__21554\,
            I => \N__21544\
        );

    \I__2371\ : Odrv4
    port map (
            O => \N__21551\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__2370\ : Odrv4
    port map (
            O => \N__21544\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__2369\ : CascadeMux
    port map (
            O => \N__21539\,
            I => \N__21536\
        );

    \I__2368\ : InMux
    port map (
            O => \N__21536\,
            I => \N__21533\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__21533\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\
        );

    \I__2366\ : CascadeMux
    port map (
            O => \N__21530\,
            I => \N__21527\
        );

    \I__2365\ : InMux
    port map (
            O => \N__21527\,
            I => \N__21524\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__21524\,
            I => \N__21519\
        );

    \I__2363\ : InMux
    port map (
            O => \N__21523\,
            I => \N__21516\
        );

    \I__2362\ : InMux
    port map (
            O => \N__21522\,
            I => \N__21513\
        );

    \I__2361\ : Span4Mux_v
    port map (
            O => \N__21519\,
            I => \N__21506\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__21516\,
            I => \N__21506\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__21513\,
            I => \N__21506\
        );

    \I__2358\ : Span4Mux_v
    port map (
            O => \N__21506\,
            I => \N__21503\
        );

    \I__2357\ : Odrv4
    port map (
            O => \N__21503\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__2356\ : InMux
    port map (
            O => \N__21500\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\
        );

    \I__2355\ : InMux
    port map (
            O => \N__21497\,
            I => \N__21494\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__21494\,
            I => \N__21491\
        );

    \I__2353\ : Odrv4
    port map (
            O => \N__21491\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\
        );

    \I__2352\ : CascadeMux
    port map (
            O => \N__21488\,
            I => \N__21483\
        );

    \I__2351\ : InMux
    port map (
            O => \N__21487\,
            I => \N__21480\
        );

    \I__2350\ : InMux
    port map (
            O => \N__21486\,
            I => \N__21476\
        );

    \I__2349\ : InMux
    port map (
            O => \N__21483\,
            I => \N__21473\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__21480\,
            I => \N__21470\
        );

    \I__2347\ : InMux
    port map (
            O => \N__21479\,
            I => \N__21467\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__21476\,
            I => \N__21464\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__21473\,
            I => \N__21461\
        );

    \I__2344\ : Span4Mux_h
    port map (
            O => \N__21470\,
            I => \N__21454\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__21467\,
            I => \N__21454\
        );

    \I__2342\ : Span4Mux_h
    port map (
            O => \N__21464\,
            I => \N__21454\
        );

    \I__2341\ : Odrv4
    port map (
            O => \N__21461\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__2340\ : Odrv4
    port map (
            O => \N__21454\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__2339\ : CascadeMux
    port map (
            O => \N__21449\,
            I => \N__21446\
        );

    \I__2338\ : InMux
    port map (
            O => \N__21446\,
            I => \N__21443\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__21443\,
            I => \N__21438\
        );

    \I__2336\ : InMux
    port map (
            O => \N__21442\,
            I => \N__21435\
        );

    \I__2335\ : InMux
    port map (
            O => \N__21441\,
            I => \N__21432\
        );

    \I__2334\ : Span4Mux_v
    port map (
            O => \N__21438\,
            I => \N__21425\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__21435\,
            I => \N__21425\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__21432\,
            I => \N__21425\
        );

    \I__2331\ : Span4Mux_v
    port map (
            O => \N__21425\,
            I => \N__21422\
        );

    \I__2330\ : Odrv4
    port map (
            O => \N__21422\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__2329\ : InMux
    port map (
            O => \N__21419\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\
        );

    \I__2328\ : CascadeMux
    port map (
            O => \N__21416\,
            I => \N__21413\
        );

    \I__2327\ : InMux
    port map (
            O => \N__21413\,
            I => \N__21410\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__21410\,
            I => \N__21407\
        );

    \I__2325\ : Span4Mux_h
    port map (
            O => \N__21407\,
            I => \N__21404\
        );

    \I__2324\ : Odrv4
    port map (
            O => \N__21404\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\
        );

    \I__2323\ : CascadeMux
    port map (
            O => \N__21401\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433_cascade_\
        );

    \I__2322\ : InMux
    port map (
            O => \N__21398\,
            I => \N__21394\
        );

    \I__2321\ : InMux
    port map (
            O => \N__21397\,
            I => \N__21390\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__21394\,
            I => \N__21387\
        );

    \I__2319\ : InMux
    port map (
            O => \N__21393\,
            I => \N__21384\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__21390\,
            I => \pwm_generator_inst.un15_threshold_1_axb_13\
        );

    \I__2317\ : Odrv4
    port map (
            O => \N__21387\,
            I => \pwm_generator_inst.un15_threshold_1_axb_13\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__21384\,
            I => \pwm_generator_inst.un15_threshold_1_axb_13\
        );

    \I__2315\ : CascadeMux
    port map (
            O => \N__21377\,
            I => \N__21374\
        );

    \I__2314\ : InMux
    port map (
            O => \N__21374\,
            I => \N__21371\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__21371\,
            I => \N__21368\
        );

    \I__2312\ : Span4Mux_h
    port map (
            O => \N__21368\,
            I => \N__21365\
        );

    \I__2311\ : Odrv4
    port map (
            O => \N__21365\,
            I => \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\
        );

    \I__2310\ : InMux
    port map (
            O => \N__21362\,
            I => \N__21359\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__21359\,
            I => \pwm_generator_inst.un19_threshold_axb_3\
        );

    \I__2308\ : InMux
    port map (
            O => \N__21356\,
            I => \N__21353\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__21353\,
            I => \N__21350\
        );

    \I__2306\ : Odrv4
    port map (
            O => \N__21350\,
            I => \pwm_generator_inst.un1_duty_inputlt3\
        );

    \I__2305\ : InMux
    port map (
            O => \N__21347\,
            I => \N__21344\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__21344\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0\
        );

    \I__2303\ : InMux
    port map (
            O => \N__21341\,
            I => \N__21338\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__21338\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\
        );

    \I__2301\ : InMux
    port map (
            O => \N__21335\,
            I => \N__21329\
        );

    \I__2300\ : InMux
    port map (
            O => \N__21334\,
            I => \N__21329\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__21329\,
            I => \N__21325\
        );

    \I__2298\ : InMux
    port map (
            O => \N__21328\,
            I => \N__21322\
        );

    \I__2297\ : Span4Mux_v
    port map (
            O => \N__21325\,
            I => \N__21319\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__21322\,
            I => \N__21316\
        );

    \I__2295\ : Odrv4
    port map (
            O => \N__21319\,
            I => pwm_duty_input_9
        );

    \I__2294\ : Odrv4
    port map (
            O => \N__21316\,
            I => pwm_duty_input_9
        );

    \I__2293\ : CascadeMux
    port map (
            O => \N__21311\,
            I => \N__21307\
        );

    \I__2292\ : InMux
    port map (
            O => \N__21310\,
            I => \N__21301\
        );

    \I__2291\ : InMux
    port map (
            O => \N__21307\,
            I => \N__21301\
        );

    \I__2290\ : InMux
    port map (
            O => \N__21306\,
            I => \N__21298\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__21301\,
            I => \N__21295\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__21298\,
            I => \N__21292\
        );

    \I__2287\ : Span4Mux_h
    port map (
            O => \N__21295\,
            I => \N__21289\
        );

    \I__2286\ : Span4Mux_s1_h
    port map (
            O => \N__21292\,
            I => \N__21286\
        );

    \I__2285\ : Odrv4
    port map (
            O => \N__21289\,
            I => pwm_duty_input_8
        );

    \I__2284\ : Odrv4
    port map (
            O => \N__21286\,
            I => pwm_duty_input_8
        );

    \I__2283\ : CascadeMux
    port map (
            O => \N__21281\,
            I => \N__21278\
        );

    \I__2282\ : InMux
    port map (
            O => \N__21278\,
            I => \N__21271\
        );

    \I__2281\ : InMux
    port map (
            O => \N__21277\,
            I => \N__21271\
        );

    \I__2280\ : InMux
    port map (
            O => \N__21276\,
            I => \N__21268\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__21271\,
            I => \N__21265\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__21268\,
            I => \N__21262\
        );

    \I__2277\ : Span4Mux_h
    port map (
            O => \N__21265\,
            I => \N__21259\
        );

    \I__2276\ : Span4Mux_v
    port map (
            O => \N__21262\,
            I => \N__21256\
        );

    \I__2275\ : Odrv4
    port map (
            O => \N__21259\,
            I => pwm_duty_input_6
        );

    \I__2274\ : Odrv4
    port map (
            O => \N__21256\,
            I => pwm_duty_input_6
        );

    \I__2273\ : InMux
    port map (
            O => \N__21251\,
            I => \N__21247\
        );

    \I__2272\ : InMux
    port map (
            O => \N__21250\,
            I => \N__21244\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__21247\,
            I => \N__21241\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__21244\,
            I => \N__21237\
        );

    \I__2269\ : Span4Mux_v
    port map (
            O => \N__21241\,
            I => \N__21234\
        );

    \I__2268\ : InMux
    port map (
            O => \N__21240\,
            I => \N__21231\
        );

    \I__2267\ : Span4Mux_s1_h
    port map (
            O => \N__21237\,
            I => \N__21228\
        );

    \I__2266\ : Odrv4
    port map (
            O => \N__21234\,
            I => pwm_duty_input_7
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__21231\,
            I => pwm_duty_input_7
        );

    \I__2264\ : Odrv4
    port map (
            O => \N__21228\,
            I => pwm_duty_input_7
        );

    \I__2263\ : InMux
    port map (
            O => \N__21221\,
            I => \N__21218\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__21218\,
            I => \N__21215\
        );

    \I__2261\ : Odrv4
    port map (
            O => \N__21215\,
            I => \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\
        );

    \I__2260\ : InMux
    port map (
            O => \N__21212\,
            I => \N__21207\
        );

    \I__2259\ : InMux
    port map (
            O => \N__21211\,
            I => \N__21204\
        );

    \I__2258\ : InMux
    port map (
            O => \N__21210\,
            I => \N__21201\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__21207\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__21204\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__21201\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__2254\ : InMux
    port map (
            O => \N__21194\,
            I => \N__21191\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__21191\,
            I => \N__21188\
        );

    \I__2252\ : Odrv4
    port map (
            O => \N__21188\,
            I => \pwm_generator_inst.un19_threshold_axb_2\
        );

    \I__2251\ : CascadeMux
    port map (
            O => \N__21185\,
            I => \N__21182\
        );

    \I__2250\ : InMux
    port map (
            O => \N__21182\,
            I => \N__21179\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__21179\,
            I => \N__21176\
        );

    \I__2248\ : Odrv4
    port map (
            O => \N__21176\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\
        );

    \I__2247\ : CascadeMux
    port map (
            O => \N__21173\,
            I => \N__21170\
        );

    \I__2246\ : InMux
    port map (
            O => \N__21170\,
            I => \N__21167\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__21167\,
            I => \N__21164\
        );

    \I__2244\ : Span4Mux_v
    port map (
            O => \N__21164\,
            I => \N__21161\
        );

    \I__2243\ : Odrv4
    port map (
            O => \N__21161\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\
        );

    \I__2242\ : InMux
    port map (
            O => \N__21158\,
            I => \pwm_generator_inst.un19_threshold_cry_1\
        );

    \I__2241\ : InMux
    port map (
            O => \N__21155\,
            I => \pwm_generator_inst.un19_threshold_cry_2\
        );

    \I__2240\ : InMux
    port map (
            O => \N__21152\,
            I => \N__21149\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__21149\,
            I => \pwm_generator_inst.un19_threshold_axb_4\
        );

    \I__2238\ : InMux
    port map (
            O => \N__21146\,
            I => \pwm_generator_inst.un19_threshold_cry_3\
        );

    \I__2237\ : InMux
    port map (
            O => \N__21143\,
            I => \N__21140\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__21140\,
            I => \pwm_generator_inst.un19_threshold_axb_5\
        );

    \I__2235\ : InMux
    port map (
            O => \N__21137\,
            I => \pwm_generator_inst.un19_threshold_cry_4\
        );

    \I__2234\ : InMux
    port map (
            O => \N__21134\,
            I => \N__21131\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__21131\,
            I => \pwm_generator_inst.un19_threshold_axb_6\
        );

    \I__2232\ : InMux
    port map (
            O => \N__21128\,
            I => \pwm_generator_inst.un19_threshold_cry_5\
        );

    \I__2231\ : InMux
    port map (
            O => \N__21125\,
            I => \N__21122\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__21122\,
            I => \pwm_generator_inst.un19_threshold_axb_7\
        );

    \I__2229\ : InMux
    port map (
            O => \N__21119\,
            I => \pwm_generator_inst.un19_threshold_cry_6\
        );

    \I__2228\ : InMux
    port map (
            O => \N__21116\,
            I => \N__21113\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__21113\,
            I => \pwm_generator_inst.un19_threshold_axb_8\
        );

    \I__2226\ : InMux
    port map (
            O => \N__21110\,
            I => \bfn_3_24_0_\
        );

    \I__2225\ : InMux
    port map (
            O => \N__21107\,
            I => \N__21104\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__21104\,
            I => \N__21101\
        );

    \I__2223\ : Span4Mux_v
    port map (
            O => \N__21101\,
            I => \N__21098\
        );

    \I__2222\ : Odrv4
    port map (
            O => \N__21098\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\
        );

    \I__2221\ : InMux
    port map (
            O => \N__21095\,
            I => \pwm_generator_inst.un19_threshold_cry_8\
        );

    \I__2220\ : CascadeMux
    port map (
            O => \N__21092\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\
        );

    \I__2219\ : InMux
    port map (
            O => \N__21089\,
            I => \N__21086\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__21086\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\
        );

    \I__2217\ : InMux
    port map (
            O => \N__21083\,
            I => \N__21080\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__21080\,
            I => \N__21077\
        );

    \I__2215\ : Odrv4
    port map (
            O => \N__21077\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9\
        );

    \I__2214\ : CascadeMux
    port map (
            O => \N__21074\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_\
        );

    \I__2213\ : InMux
    port map (
            O => \N__21071\,
            I => \N__21068\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__21068\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\
        );

    \I__2211\ : InMux
    port map (
            O => \N__21065\,
            I => \N__21056\
        );

    \I__2210\ : InMux
    port map (
            O => \N__21064\,
            I => \N__21051\
        );

    \I__2209\ : InMux
    port map (
            O => \N__21063\,
            I => \N__21051\
        );

    \I__2208\ : InMux
    port map (
            O => \N__21062\,
            I => \N__21044\
        );

    \I__2207\ : InMux
    port map (
            O => \N__21061\,
            I => \N__21044\
        );

    \I__2206\ : InMux
    port map (
            O => \N__21060\,
            I => \N__21044\
        );

    \I__2205\ : InMux
    port map (
            O => \N__21059\,
            I => \N__21041\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__21056\,
            I => \N__21036\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__21051\,
            I => \N__21036\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__21044\,
            I => \N__21033\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__21041\,
            I => \N__21030\
        );

    \I__2200\ : Span4Mux_v
    port map (
            O => \N__21036\,
            I => \N__21027\
        );

    \I__2199\ : Span4Mux_s3_h
    port map (
            O => \N__21033\,
            I => \N__21024\
        );

    \I__2198\ : Span4Mux_s3_h
    port map (
            O => \N__21030\,
            I => \N__21021\
        );

    \I__2197\ : Odrv4
    port map (
            O => \N__21027\,
            I => \current_shift_inst.PI_CTRL.N_159\
        );

    \I__2196\ : Odrv4
    port map (
            O => \N__21024\,
            I => \current_shift_inst.PI_CTRL.N_159\
        );

    \I__2195\ : Odrv4
    port map (
            O => \N__21021\,
            I => \current_shift_inst.PI_CTRL.N_159\
        );

    \I__2194\ : InMux
    port map (
            O => \N__21014\,
            I => \N__21011\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__21011\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\
        );

    \I__2192\ : CascadeMux
    port map (
            O => \N__21008\,
            I => \N__21005\
        );

    \I__2191\ : InMux
    port map (
            O => \N__21005\,
            I => \N__21002\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__21002\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\
        );

    \I__2189\ : InMux
    port map (
            O => \N__20999\,
            I => \N__20996\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__20996\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\
        );

    \I__2187\ : InMux
    port map (
            O => \N__20993\,
            I => \N__20990\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__20990\,
            I => \N__20987\
        );

    \I__2185\ : Span4Mux_v
    port map (
            O => \N__20987\,
            I => \N__20984\
        );

    \I__2184\ : Odrv4
    port map (
            O => \N__20984\,
            I => \pwm_generator_inst.un19_threshold_axb_1\
        );

    \I__2183\ : InMux
    port map (
            O => \N__20981\,
            I => \pwm_generator_inst.un19_threshold_cry_0\
        );

    \I__2182\ : CascadeMux
    port map (
            O => \N__20978\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_\
        );

    \I__2181\ : InMux
    port map (
            O => \N__20975\,
            I => \N__20972\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__20972\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\
        );

    \I__2179\ : InMux
    port map (
            O => \N__20969\,
            I => \N__20966\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__20966\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_7\
        );

    \I__2177\ : CascadeMux
    port map (
            O => \N__20963\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_\
        );

    \I__2176\ : InMux
    port map (
            O => \N__20960\,
            I => \N__20957\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__20957\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\
        );

    \I__2174\ : InMux
    port map (
            O => \N__20954\,
            I => \N__20951\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__20951\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\
        );

    \I__2172\ : InMux
    port map (
            O => \N__20948\,
            I => \N__20945\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__20945\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\
        );

    \I__2170\ : CascadeMux
    port map (
            O => \N__20942\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_\
        );

    \I__2169\ : InMux
    port map (
            O => \N__20939\,
            I => \N__20936\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__20936\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\
        );

    \I__2167\ : CascadeMux
    port map (
            O => \N__20933\,
            I => \N__20930\
        );

    \I__2166\ : InMux
    port map (
            O => \N__20930\,
            I => \N__20927\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__20927\,
            I => \N__20924\
        );

    \I__2164\ : Odrv4
    port map (
            O => \N__20924\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\
        );

    \I__2163\ : CascadeMux
    port map (
            O => \N__20921\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\
        );

    \I__2162\ : CascadeMux
    port map (
            O => \N__20918\,
            I => \current_shift_inst.PI_CTRL.N_44_cascade_\
        );

    \I__2161\ : InMux
    port map (
            O => \N__20915\,
            I => \N__20912\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__20912\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\
        );

    \I__2159\ : CascadeMux
    port map (
            O => \N__20909\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19_cascade_\
        );

    \I__2158\ : InMux
    port map (
            O => \N__20906\,
            I => \N__20903\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__20903\,
            I => \N__20900\
        );

    \I__2156\ : Odrv4
    port map (
            O => \N__20900\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\
        );

    \I__2155\ : InMux
    port map (
            O => \N__20897\,
            I => \N__20894\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__20894\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\
        );

    \I__2153\ : InMux
    port map (
            O => \N__20891\,
            I => \N__20888\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__20888\,
            I => \current_shift_inst.PI_CTRL.N_77\
        );

    \I__2151\ : InMux
    port map (
            O => \N__20885\,
            I => \N__20881\
        );

    \I__2150\ : InMux
    port map (
            O => \N__20884\,
            I => \N__20877\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__20881\,
            I => \N__20874\
        );

    \I__2148\ : InMux
    port map (
            O => \N__20880\,
            I => \N__20871\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__20877\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__2146\ : Odrv12
    port map (
            O => \N__20874\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__20871\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__2144\ : InMux
    port map (
            O => \N__20864\,
            I => \N__20861\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__20861\,
            I => \N__20858\
        );

    \I__2142\ : Span4Mux_s1_v
    port map (
            O => \N__20858\,
            I => \N__20855\
        );

    \I__2141\ : Odrv4
    port map (
            O => \N__20855\,
            I => \rgb_drv_RNOZ0\
        );

    \I__2140\ : CascadeMux
    port map (
            O => \N__20852\,
            I => \N__20849\
        );

    \I__2139\ : InMux
    port map (
            O => \N__20849\,
            I => \N__20846\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__20846\,
            I => \N__20843\
        );

    \I__2137\ : Span4Mux_h
    port map (
            O => \N__20843\,
            I => \N__20840\
        );

    \I__2136\ : Odrv4
    port map (
            O => \N__20840\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\
        );

    \I__2135\ : InMux
    port map (
            O => \N__20837\,
            I => \N__20834\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__20834\,
            I => \N__20831\
        );

    \I__2133\ : Odrv4
    port map (
            O => \N__20831\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\
        );

    \I__2132\ : CascadeMux
    port map (
            O => \N__20828\,
            I => \N__20825\
        );

    \I__2131\ : InMux
    port map (
            O => \N__20825\,
            I => \N__20822\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__20822\,
            I => \N__20819\
        );

    \I__2129\ : Span4Mux_h
    port map (
            O => \N__20819\,
            I => \N__20816\
        );

    \I__2128\ : Odrv4
    port map (
            O => \N__20816\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\
        );

    \I__2127\ : CascadeMux
    port map (
            O => \N__20813\,
            I => \N__20810\
        );

    \I__2126\ : InMux
    port map (
            O => \N__20810\,
            I => \N__20807\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__20807\,
            I => \N__20804\
        );

    \I__2124\ : Span4Mux_v
    port map (
            O => \N__20804\,
            I => \N__20801\
        );

    \I__2123\ : Odrv4
    port map (
            O => \N__20801\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\
        );

    \I__2122\ : InMux
    port map (
            O => \N__20798\,
            I => \N__20794\
        );

    \I__2121\ : CascadeMux
    port map (
            O => \N__20797\,
            I => \N__20791\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__20794\,
            I => \N__20788\
        );

    \I__2119\ : InMux
    port map (
            O => \N__20791\,
            I => \N__20785\
        );

    \I__2118\ : Span4Mux_h
    port map (
            O => \N__20788\,
            I => \N__20780\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__20785\,
            I => \N__20780\
        );

    \I__2116\ : Span4Mux_v
    port map (
            O => \N__20780\,
            I => \N__20777\
        );

    \I__2115\ : Odrv4
    port map (
            O => \N__20777\,
            I => \current_shift_inst.PI_CTRL.un1_integrator\
        );

    \I__2114\ : CascadeMux
    port map (
            O => \N__20774\,
            I => \N__20771\
        );

    \I__2113\ : InMux
    port map (
            O => \N__20771\,
            I => \N__20768\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__20768\,
            I => \N__20765\
        );

    \I__2111\ : Span4Mux_h
    port map (
            O => \N__20765\,
            I => \N__20762\
        );

    \I__2110\ : Odrv4
    port map (
            O => \N__20762\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\
        );

    \I__2109\ : InMux
    port map (
            O => \N__20759\,
            I => \N__20756\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__20756\,
            I => \N__20753\
        );

    \I__2107\ : Span4Mux_v
    port map (
            O => \N__20753\,
            I => \N__20750\
        );

    \I__2106\ : Odrv4
    port map (
            O => \N__20750\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\
        );

    \I__2105\ : InMux
    port map (
            O => \N__20747\,
            I => \N__20744\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__20744\,
            I => \N__20741\
        );

    \I__2103\ : Odrv4
    port map (
            O => \N__20741\,
            I => \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\
        );

    \I__2102\ : InMux
    port map (
            O => \N__20738\,
            I => \N__20735\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__20735\,
            I => \N__20732\
        );

    \I__2100\ : Odrv4
    port map (
            O => \N__20732\,
            I => \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\
        );

    \I__2099\ : InMux
    port map (
            O => \N__20729\,
            I => \N__20726\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__20726\,
            I => \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\
        );

    \I__2097\ : InMux
    port map (
            O => \N__20723\,
            I => \N__20718\
        );

    \I__2096\ : InMux
    port map (
            O => \N__20722\,
            I => \N__20715\
        );

    \I__2095\ : InMux
    port map (
            O => \N__20721\,
            I => \N__20712\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__20718\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__20715\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__20712\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__2091\ : CascadeMux
    port map (
            O => \N__20705\,
            I => \N__20702\
        );

    \I__2090\ : InMux
    port map (
            O => \N__20702\,
            I => \N__20698\
        );

    \I__2089\ : InMux
    port map (
            O => \N__20701\,
            I => \N__20694\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__20698\,
            I => \N__20691\
        );

    \I__2087\ : InMux
    port map (
            O => \N__20697\,
            I => \N__20688\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__20694\,
            I => \pwm_generator_inst.un15_threshold_1_axb_16\
        );

    \I__2085\ : Odrv4
    port map (
            O => \N__20691\,
            I => \pwm_generator_inst.un15_threshold_1_axb_16\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__20688\,
            I => \pwm_generator_inst.un15_threshold_1_axb_16\
        );

    \I__2083\ : InMux
    port map (
            O => \N__20681\,
            I => \N__20677\
        );

    \I__2082\ : InMux
    port map (
            O => \N__20680\,
            I => \N__20673\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__20677\,
            I => \N__20670\
        );

    \I__2080\ : InMux
    port map (
            O => \N__20676\,
            I => \N__20667\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__20673\,
            I => \pwm_generator_inst.un15_threshold_1_axb_17\
        );

    \I__2078\ : Odrv4
    port map (
            O => \N__20670\,
            I => \pwm_generator_inst.un15_threshold_1_axb_17\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__20667\,
            I => \pwm_generator_inst.un15_threshold_1_axb_17\
        );

    \I__2076\ : InMux
    port map (
            O => \N__20660\,
            I => \N__20657\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__20657\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\
        );

    \I__2074\ : CascadeMux
    port map (
            O => \N__20654\,
            I => \N__20647\
        );

    \I__2073\ : InMux
    port map (
            O => \N__20653\,
            I => \N__20640\
        );

    \I__2072\ : InMux
    port map (
            O => \N__20652\,
            I => \N__20640\
        );

    \I__2071\ : InMux
    port map (
            O => \N__20651\,
            I => \N__20640\
        );

    \I__2070\ : InMux
    port map (
            O => \N__20650\,
            I => \N__20632\
        );

    \I__2069\ : InMux
    port map (
            O => \N__20647\,
            I => \N__20632\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__20640\,
            I => \N__20629\
        );

    \I__2067\ : InMux
    port map (
            O => \N__20639\,
            I => \N__20622\
        );

    \I__2066\ : InMux
    port map (
            O => \N__20638\,
            I => \N__20622\
        );

    \I__2065\ : InMux
    port map (
            O => \N__20637\,
            I => \N__20622\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__20632\,
            I => \N__20615\
        );

    \I__2063\ : Span4Mux_v
    port map (
            O => \N__20629\,
            I => \N__20615\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__20622\,
            I => \N__20615\
        );

    \I__2061\ : Odrv4
    port map (
            O => \N__20615\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\
        );

    \I__2060\ : CascadeMux
    port map (
            O => \N__20612\,
            I => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\
        );

    \I__2059\ : CascadeMux
    port map (
            O => \N__20609\,
            I => \N__20605\
        );

    \I__2058\ : CascadeMux
    port map (
            O => \N__20608\,
            I => \N__20602\
        );

    \I__2057\ : InMux
    port map (
            O => \N__20605\,
            I => \N__20598\
        );

    \I__2056\ : InMux
    port map (
            O => \N__20602\,
            I => \N__20593\
        );

    \I__2055\ : InMux
    port map (
            O => \N__20601\,
            I => \N__20593\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__20598\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__20593\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__2052\ : InMux
    port map (
            O => \N__20588\,
            I => \N__20584\
        );

    \I__2051\ : InMux
    port map (
            O => \N__20587\,
            I => \N__20581\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__20584\,
            I => \N__20578\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__20581\,
            I => pwm_duty_input_0
        );

    \I__2048\ : Odrv4
    port map (
            O => \N__20578\,
            I => pwm_duty_input_0
        );

    \I__2047\ : InMux
    port map (
            O => \N__20573\,
            I => \N__20570\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__20570\,
            I => \N__20566\
        );

    \I__2045\ : InMux
    port map (
            O => \N__20569\,
            I => \N__20563\
        );

    \I__2044\ : Span4Mux_v
    port map (
            O => \N__20566\,
            I => \N__20560\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__20563\,
            I => pwm_duty_input_1
        );

    \I__2042\ : Odrv4
    port map (
            O => \N__20560\,
            I => pwm_duty_input_1
        );

    \I__2041\ : InMux
    port map (
            O => \N__20555\,
            I => \N__20551\
        );

    \I__2040\ : InMux
    port map (
            O => \N__20554\,
            I => \N__20548\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__20551\,
            I => \N__20545\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__20548\,
            I => \N__20540\
        );

    \I__2037\ : Span4Mux_v
    port map (
            O => \N__20545\,
            I => \N__20540\
        );

    \I__2036\ : Odrv4
    port map (
            O => \N__20540\,
            I => pwm_duty_input_2
        );

    \I__2035\ : InMux
    port map (
            O => \N__20537\,
            I => \N__20534\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__20534\,
            I => \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\
        );

    \I__2033\ : CascadeMux
    port map (
            O => \N__20531\,
            I => \N__20527\
        );

    \I__2032\ : InMux
    port map (
            O => \N__20530\,
            I => \N__20524\
        );

    \I__2031\ : InMux
    port map (
            O => \N__20527\,
            I => \N__20521\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__20524\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__20521\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__2028\ : InMux
    port map (
            O => \N__20516\,
            I => \N__20513\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__20513\,
            I => \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\
        );

    \I__2026\ : CascadeMux
    port map (
            O => \N__20510\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15_cascade_\
        );

    \I__2025\ : CascadeMux
    port map (
            O => \N__20507\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_2_cascade_\
        );

    \I__2024\ : CascadeMux
    port map (
            O => \N__20504\,
            I => \current_shift_inst.PI_CTRL.N_43_cascade_\
        );

    \I__2023\ : InMux
    port map (
            O => \N__20501\,
            I => \N__20498\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__20498\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\
        );

    \I__2021\ : InMux
    port map (
            O => \N__20495\,
            I => \N__20492\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__20492\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\
        );

    \I__2019\ : CascadeMux
    port map (
            O => \N__20489\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_\
        );

    \I__2018\ : InMux
    port map (
            O => \N__20486\,
            I => \N__20483\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__20483\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\
        );

    \I__2016\ : CascadeMux
    port map (
            O => \N__20480\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_\
        );

    \I__2015\ : InMux
    port map (
            O => \N__20477\,
            I => \N__20474\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__20474\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\
        );

    \I__2013\ : InMux
    port map (
            O => \N__20471\,
            I => \N__20468\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__20468\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\
        );

    \I__2011\ : InMux
    port map (
            O => \N__20465\,
            I => \N__20462\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__20462\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\
        );

    \I__2009\ : CascadeMux
    port map (
            O => \N__20459\,
            I => \N__20456\
        );

    \I__2008\ : InMux
    port map (
            O => \N__20456\,
            I => \N__20453\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__20453\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\
        );

    \I__2006\ : InMux
    port map (
            O => \N__20450\,
            I => \N__20447\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__20447\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\
        );

    \I__2004\ : CascadeMux
    port map (
            O => \N__20444\,
            I => \N__20441\
        );

    \I__2003\ : InMux
    port map (
            O => \N__20441\,
            I => \N__20438\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__20438\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\
        );

    \I__2001\ : CascadeMux
    port map (
            O => \N__20435\,
            I => \N__20432\
        );

    \I__2000\ : InMux
    port map (
            O => \N__20432\,
            I => \N__20429\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__20429\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\
        );

    \I__1998\ : CascadeMux
    port map (
            O => \N__20426\,
            I => \N__20423\
        );

    \I__1997\ : InMux
    port map (
            O => \N__20423\,
            I => \N__20420\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__20420\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\
        );

    \I__1995\ : InMux
    port map (
            O => \N__20417\,
            I => \N__20414\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__20414\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\
        );

    \I__1993\ : CascadeMux
    port map (
            O => \N__20411\,
            I => \N__20408\
        );

    \I__1992\ : InMux
    port map (
            O => \N__20408\,
            I => \N__20405\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__20405\,
            I => \N__20402\
        );

    \I__1990\ : Odrv4
    port map (
            O => \N__20402\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\
        );

    \I__1989\ : InMux
    port map (
            O => \N__20399\,
            I => \pwm_generator_inst.un15_threshold_1_cry_17\
        );

    \I__1988\ : InMux
    port map (
            O => \N__20396\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18\
        );

    \I__1987\ : InMux
    port map (
            O => \N__20393\,
            I => \N__20390\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__20390\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\
        );

    \I__1985\ : InMux
    port map (
            O => \N__20387\,
            I => \N__20384\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__20384\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\
        );

    \I__1983\ : CascadeMux
    port map (
            O => \N__20381\,
            I => \N__20378\
        );

    \I__1982\ : InMux
    port map (
            O => \N__20378\,
            I => \N__20375\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__20375\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\
        );

    \I__1980\ : CascadeMux
    port map (
            O => \N__20372\,
            I => \N__20369\
        );

    \I__1979\ : InMux
    port map (
            O => \N__20369\,
            I => \N__20366\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__20366\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\
        );

    \I__1977\ : InMux
    port map (
            O => \N__20363\,
            I => \N__20360\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__20360\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\
        );

    \I__1975\ : InMux
    port map (
            O => \N__20357\,
            I => \N__20354\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__20354\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\
        );

    \I__1973\ : CascadeMux
    port map (
            O => \N__20351\,
            I => \N__20348\
        );

    \I__1972\ : InMux
    port map (
            O => \N__20348\,
            I => \N__20345\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__20345\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\
        );

    \I__1970\ : InMux
    port map (
            O => \N__20342\,
            I => \N__20339\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__20339\,
            I => \pwm_generator_inst.O_9\
        );

    \I__1968\ : InMux
    port map (
            O => \N__20336\,
            I => \N__20333\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__20333\,
            I => \pwm_generator_inst.un15_threshold_1_axb_9\
        );

    \I__1966\ : InMux
    port map (
            O => \N__20330\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9\
        );

    \I__1965\ : InMux
    port map (
            O => \N__20327\,
            I => \pwm_generator_inst.un15_threshold_1_cry_10\
        );

    \I__1964\ : InMux
    port map (
            O => \N__20324\,
            I => \pwm_generator_inst.un15_threshold_1_cry_11\
        );

    \I__1963\ : InMux
    port map (
            O => \N__20321\,
            I => \pwm_generator_inst.un15_threshold_1_cry_12\
        );

    \I__1962\ : InMux
    port map (
            O => \N__20318\,
            I => \pwm_generator_inst.un15_threshold_1_cry_13\
        );

    \I__1961\ : InMux
    port map (
            O => \N__20315\,
            I => \pwm_generator_inst.un15_threshold_1_cry_14\
        );

    \I__1960\ : InMux
    port map (
            O => \N__20312\,
            I => \bfn_1_26_0_\
        );

    \I__1959\ : InMux
    port map (
            O => \N__20309\,
            I => \pwm_generator_inst.un15_threshold_1_cry_16\
        );

    \I__1958\ : InMux
    port map (
            O => \N__20306\,
            I => \N__20303\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__20303\,
            I => \pwm_generator_inst.O_1\
        );

    \I__1956\ : InMux
    port map (
            O => \N__20300\,
            I => \N__20297\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__20297\,
            I => \pwm_generator_inst.un15_threshold_1_axb_1\
        );

    \I__1954\ : InMux
    port map (
            O => \N__20294\,
            I => \N__20291\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__20291\,
            I => \pwm_generator_inst.O_2\
        );

    \I__1952\ : InMux
    port map (
            O => \N__20288\,
            I => \N__20285\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__20285\,
            I => \pwm_generator_inst.un15_threshold_1_axb_2\
        );

    \I__1950\ : InMux
    port map (
            O => \N__20282\,
            I => \N__20279\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__20279\,
            I => \pwm_generator_inst.O_3\
        );

    \I__1948\ : InMux
    port map (
            O => \N__20276\,
            I => \N__20273\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__20273\,
            I => \pwm_generator_inst.un15_threshold_1_axb_3\
        );

    \I__1946\ : InMux
    port map (
            O => \N__20270\,
            I => \N__20267\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__20267\,
            I => \pwm_generator_inst.O_4\
        );

    \I__1944\ : InMux
    port map (
            O => \N__20264\,
            I => \N__20261\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__20261\,
            I => \pwm_generator_inst.un15_threshold_1_axb_4\
        );

    \I__1942\ : InMux
    port map (
            O => \N__20258\,
            I => \N__20255\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__20255\,
            I => \pwm_generator_inst.O_5\
        );

    \I__1940\ : InMux
    port map (
            O => \N__20252\,
            I => \N__20249\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__20249\,
            I => \pwm_generator_inst.un15_threshold_1_axb_5\
        );

    \I__1938\ : InMux
    port map (
            O => \N__20246\,
            I => \N__20243\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__20243\,
            I => \pwm_generator_inst.O_6\
        );

    \I__1936\ : InMux
    port map (
            O => \N__20240\,
            I => \N__20237\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__20237\,
            I => \pwm_generator_inst.un15_threshold_1_axb_6\
        );

    \I__1934\ : InMux
    port map (
            O => \N__20234\,
            I => \N__20231\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__20231\,
            I => \pwm_generator_inst.O_7\
        );

    \I__1932\ : InMux
    port map (
            O => \N__20228\,
            I => \N__20225\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__20225\,
            I => \pwm_generator_inst.un15_threshold_1_axb_7\
        );

    \I__1930\ : InMux
    port map (
            O => \N__20222\,
            I => \N__20219\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__20219\,
            I => \pwm_generator_inst.O_8\
        );

    \I__1928\ : InMux
    port map (
            O => \N__20216\,
            I => \N__20213\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__20213\,
            I => \pwm_generator_inst.un15_threshold_1_axb_8\
        );

    \I__1926\ : InMux
    port map (
            O => \N__20210\,
            I => \N__20207\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__20207\,
            I => \current_shift_inst.PI_CTRL.N_96\
        );

    \I__1924\ : InMux
    port map (
            O => \N__20204\,
            I => \N__20200\
        );

    \I__1923\ : InMux
    port map (
            O => \N__20203\,
            I => \N__20197\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__20200\,
            I => \current_shift_inst.PI_CTRL.N_94\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__20197\,
            I => \current_shift_inst.PI_CTRL.N_94\
        );

    \I__1920\ : CascadeMux
    port map (
            O => \N__20192\,
            I => \N__20189\
        );

    \I__1919\ : InMux
    port map (
            O => \N__20189\,
            I => \N__20186\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__20186\,
            I => \N__20182\
        );

    \I__1917\ : InMux
    port map (
            O => \N__20185\,
            I => \N__20179\
        );

    \I__1916\ : Odrv4
    port map (
            O => \N__20182\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__20179\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__1914\ : InMux
    port map (
            O => \N__20174\,
            I => \N__20171\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__20171\,
            I => \current_shift_inst.PI_CTRL.N_91\
        );

    \I__1912\ : InMux
    port map (
            O => \N__20168\,
            I => \N__20159\
        );

    \I__1911\ : InMux
    port map (
            O => \N__20167\,
            I => \N__20159\
        );

    \I__1910\ : InMux
    port map (
            O => \N__20166\,
            I => \N__20159\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__20159\,
            I => \current_shift_inst.PI_CTRL.N_161\
        );

    \I__1908\ : InMux
    port map (
            O => \N__20156\,
            I => \N__20153\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__20153\,
            I => \pwm_generator_inst.O_0\
        );

    \I__1906\ : InMux
    port map (
            O => \N__20150\,
            I => \N__20147\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__20147\,
            I => \pwm_generator_inst.un15_threshold_1_axb_0\
        );

    \I__1904\ : CascadeMux
    port map (
            O => \N__20144\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_\
        );

    \I__1903\ : CascadeMux
    port map (
            O => \N__20141\,
            I => \current_shift_inst.PI_CTRL.N_98_cascade_\
        );

    \I__1902\ : CascadeMux
    port map (
            O => \N__20138\,
            I => \current_shift_inst.PI_CTRL.N_96_cascade_\
        );

    \I__1901\ : InMux
    port map (
            O => \N__20135\,
            I => \N__20132\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__20132\,
            I => \current_shift_inst.PI_CTRL.N_97\
        );

    \I__1899\ : InMux
    port map (
            O => \N__20129\,
            I => \N__20126\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__20126\,
            I => \N__20123\
        );

    \I__1897\ : Odrv12
    port map (
            O => \N__20123\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\
        );

    \I__1896\ : CascadeMux
    port map (
            O => \N__20120\,
            I => \N__20117\
        );

    \I__1895\ : InMux
    port map (
            O => \N__20117\,
            I => \N__20114\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__20114\,
            I => \N__20111\
        );

    \I__1893\ : Span4Mux_v
    port map (
            O => \N__20111\,
            I => \N__20108\
        );

    \I__1892\ : Odrv4
    port map (
            O => \N__20108\,
            I => \current_shift_inst.PI_CTRL.integrator_1_28\
        );

    \I__1891\ : InMux
    port map (
            O => \N__20105\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\
        );

    \I__1890\ : CascadeMux
    port map (
            O => \N__20102\,
            I => \N__20099\
        );

    \I__1889\ : InMux
    port map (
            O => \N__20099\,
            I => \N__20096\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__20096\,
            I => \N__20093\
        );

    \I__1887\ : Odrv12
    port map (
            O => \N__20093\,
            I => \current_shift_inst.PI_CTRL.integrator_1_29\
        );

    \I__1886\ : InMux
    port map (
            O => \N__20090\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\
        );

    \I__1885\ : CascadeMux
    port map (
            O => \N__20087\,
            I => \N__20084\
        );

    \I__1884\ : InMux
    port map (
            O => \N__20084\,
            I => \N__20081\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__20081\,
            I => \N__20078\
        );

    \I__1882\ : Span4Mux_v
    port map (
            O => \N__20078\,
            I => \N__20075\
        );

    \I__1881\ : Odrv4
    port map (
            O => \N__20075\,
            I => \current_shift_inst.PI_CTRL.integrator_1_30\
        );

    \I__1880\ : InMux
    port map (
            O => \N__20072\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\
        );

    \I__1879\ : InMux
    port map (
            O => \N__20069\,
            I => \N__20066\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__20066\,
            I => \N__20063\
        );

    \I__1877\ : Span4Mux_v
    port map (
            O => \N__20063\,
            I => \N__20060\
        );

    \I__1876\ : Odrv4
    port map (
            O => \N__20060\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\
        );

    \I__1875\ : CascadeMux
    port map (
            O => \N__20057\,
            I => \N__20054\
        );

    \I__1874\ : InMux
    port map (
            O => \N__20054\,
            I => \N__20051\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__20051\,
            I => \N__20048\
        );

    \I__1872\ : Odrv12
    port map (
            O => \N__20048\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30\
        );

    \I__1871\ : InMux
    port map (
            O => \N__20045\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\
        );

    \I__1870\ : InMux
    port map (
            O => \N__20042\,
            I => \N__20039\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__20039\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\
        );

    \I__1868\ : CascadeMux
    port map (
            O => \N__20036\,
            I => \N__20033\
        );

    \I__1867\ : InMux
    port map (
            O => \N__20033\,
            I => \N__20030\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__20030\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\
        );

    \I__1865\ : InMux
    port map (
            O => \N__20027\,
            I => \N__20024\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__20024\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\
        );

    \I__1863\ : InMux
    port map (
            O => \N__20021\,
            I => \N__20018\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__20018\,
            I => \N__20015\
        );

    \I__1861\ : Span4Mux_v
    port map (
            O => \N__20015\,
            I => \N__20012\
        );

    \I__1860\ : Odrv4
    port map (
            O => \N__20012\,
            I => \current_shift_inst.PI_CTRL.integrator_1_19\
        );

    \I__1859\ : InMux
    port map (
            O => \N__20009\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\
        );

    \I__1858\ : InMux
    port map (
            O => \N__20006\,
            I => \N__20003\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__20003\,
            I => \N__20000\
        );

    \I__1856\ : Odrv12
    port map (
            O => \N__20000\,
            I => \current_shift_inst.PI_CTRL.integrator_1_20\
        );

    \I__1855\ : InMux
    port map (
            O => \N__19997\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\
        );

    \I__1854\ : CascadeMux
    port map (
            O => \N__19994\,
            I => \N__19991\
        );

    \I__1853\ : InMux
    port map (
            O => \N__19991\,
            I => \N__19988\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__19988\,
            I => \N__19985\
        );

    \I__1851\ : Span4Mux_v
    port map (
            O => \N__19985\,
            I => \N__19982\
        );

    \I__1850\ : Odrv4
    port map (
            O => \N__19982\,
            I => \current_shift_inst.PI_CTRL.integrator_1_21\
        );

    \I__1849\ : InMux
    port map (
            O => \N__19979\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\
        );

    \I__1848\ : CascadeMux
    port map (
            O => \N__19976\,
            I => \N__19973\
        );

    \I__1847\ : InMux
    port map (
            O => \N__19973\,
            I => \N__19970\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__19970\,
            I => \N__19967\
        );

    \I__1845\ : Span4Mux_v
    port map (
            O => \N__19967\,
            I => \N__19964\
        );

    \I__1844\ : Odrv4
    port map (
            O => \N__19964\,
            I => \current_shift_inst.PI_CTRL.integrator_1_22\
        );

    \I__1843\ : InMux
    port map (
            O => \N__19961\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\
        );

    \I__1842\ : CascadeMux
    port map (
            O => \N__19958\,
            I => \N__19955\
        );

    \I__1841\ : InMux
    port map (
            O => \N__19955\,
            I => \N__19952\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__19952\,
            I => \N__19949\
        );

    \I__1839\ : Span4Mux_v
    port map (
            O => \N__19949\,
            I => \N__19946\
        );

    \I__1838\ : Odrv4
    port map (
            O => \N__19946\,
            I => \current_shift_inst.PI_CTRL.integrator_1_23\
        );

    \I__1837\ : InMux
    port map (
            O => \N__19943\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\
        );

    \I__1836\ : CascadeMux
    port map (
            O => \N__19940\,
            I => \N__19937\
        );

    \I__1835\ : InMux
    port map (
            O => \N__19937\,
            I => \N__19934\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__19934\,
            I => \N__19931\
        );

    \I__1833\ : Span4Mux_v
    port map (
            O => \N__19931\,
            I => \N__19928\
        );

    \I__1832\ : Odrv4
    port map (
            O => \N__19928\,
            I => \current_shift_inst.PI_CTRL.integrator_1_24\
        );

    \I__1831\ : InMux
    port map (
            O => \N__19925\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\
        );

    \I__1830\ : CascadeMux
    port map (
            O => \N__19922\,
            I => \N__19919\
        );

    \I__1829\ : InMux
    port map (
            O => \N__19919\,
            I => \N__19916\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__19916\,
            I => \N__19913\
        );

    \I__1827\ : Span4Mux_v
    port map (
            O => \N__19913\,
            I => \N__19910\
        );

    \I__1826\ : Odrv4
    port map (
            O => \N__19910\,
            I => \current_shift_inst.PI_CTRL.integrator_1_25\
        );

    \I__1825\ : InMux
    port map (
            O => \N__19907\,
            I => \bfn_1_16_0_\
        );

    \I__1824\ : CascadeMux
    port map (
            O => \N__19904\,
            I => \N__19901\
        );

    \I__1823\ : InMux
    port map (
            O => \N__19901\,
            I => \N__19898\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__19898\,
            I => \N__19895\
        );

    \I__1821\ : Span4Mux_v
    port map (
            O => \N__19895\,
            I => \N__19892\
        );

    \I__1820\ : Odrv4
    port map (
            O => \N__19892\,
            I => \current_shift_inst.PI_CTRL.integrator_1_26\
        );

    \I__1819\ : InMux
    port map (
            O => \N__19889\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\
        );

    \I__1818\ : CascadeMux
    port map (
            O => \N__19886\,
            I => \N__19883\
        );

    \I__1817\ : InMux
    port map (
            O => \N__19883\,
            I => \N__19880\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__19880\,
            I => \N__19877\
        );

    \I__1815\ : Span4Mux_v
    port map (
            O => \N__19877\,
            I => \N__19874\
        );

    \I__1814\ : Odrv4
    port map (
            O => \N__19874\,
            I => \current_shift_inst.PI_CTRL.integrator_1_27\
        );

    \I__1813\ : InMux
    port map (
            O => \N__19871\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\
        );

    \I__1812\ : CascadeMux
    port map (
            O => \N__19868\,
            I => \N__19865\
        );

    \I__1811\ : InMux
    port map (
            O => \N__19865\,
            I => \N__19862\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__19862\,
            I => \N__19859\
        );

    \I__1809\ : Odrv4
    port map (
            O => \N__19859\,
            I => \current_shift_inst.PI_CTRL.integrator_1_11\
        );

    \I__1808\ : InMux
    port map (
            O => \N__19856\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\
        );

    \I__1807\ : CascadeMux
    port map (
            O => \N__19853\,
            I => \N__19850\
        );

    \I__1806\ : InMux
    port map (
            O => \N__19850\,
            I => \N__19847\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__19847\,
            I => \N__19844\
        );

    \I__1804\ : Odrv4
    port map (
            O => \N__19844\,
            I => \current_shift_inst.PI_CTRL.integrator_1_12\
        );

    \I__1803\ : InMux
    port map (
            O => \N__19841\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\
        );

    \I__1802\ : CascadeMux
    port map (
            O => \N__19838\,
            I => \N__19835\
        );

    \I__1801\ : InMux
    port map (
            O => \N__19835\,
            I => \N__19832\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__19832\,
            I => \N__19829\
        );

    \I__1799\ : Span4Mux_v
    port map (
            O => \N__19829\,
            I => \N__19826\
        );

    \I__1798\ : Odrv4
    port map (
            O => \N__19826\,
            I => \current_shift_inst.PI_CTRL.integrator_1_13\
        );

    \I__1797\ : InMux
    port map (
            O => \N__19823\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\
        );

    \I__1796\ : CascadeMux
    port map (
            O => \N__19820\,
            I => \N__19817\
        );

    \I__1795\ : InMux
    port map (
            O => \N__19817\,
            I => \N__19814\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__19814\,
            I => \N__19811\
        );

    \I__1793\ : Odrv4
    port map (
            O => \N__19811\,
            I => \current_shift_inst.PI_CTRL.integrator_1_14\
        );

    \I__1792\ : InMux
    port map (
            O => \N__19808\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\
        );

    \I__1791\ : CascadeMux
    port map (
            O => \N__19805\,
            I => \N__19802\
        );

    \I__1790\ : InMux
    port map (
            O => \N__19802\,
            I => \N__19799\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__19799\,
            I => \N__19796\
        );

    \I__1788\ : Span4Mux_h
    port map (
            O => \N__19796\,
            I => \N__19793\
        );

    \I__1787\ : Odrv4
    port map (
            O => \N__19793\,
            I => \current_shift_inst.PI_CTRL.integrator_1_15\
        );

    \I__1786\ : InMux
    port map (
            O => \N__19790\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\
        );

    \I__1785\ : CascadeMux
    port map (
            O => \N__19787\,
            I => \N__19784\
        );

    \I__1784\ : InMux
    port map (
            O => \N__19784\,
            I => \N__19781\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__19781\,
            I => \N__19778\
        );

    \I__1782\ : Odrv12
    port map (
            O => \N__19778\,
            I => \current_shift_inst.PI_CTRL.integrator_1_16\
        );

    \I__1781\ : InMux
    port map (
            O => \N__19775\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\
        );

    \I__1780\ : CascadeMux
    port map (
            O => \N__19772\,
            I => \N__19769\
        );

    \I__1779\ : InMux
    port map (
            O => \N__19769\,
            I => \N__19766\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__19766\,
            I => \N__19763\
        );

    \I__1777\ : Span4Mux_v
    port map (
            O => \N__19763\,
            I => \N__19760\
        );

    \I__1776\ : Odrv4
    port map (
            O => \N__19760\,
            I => \current_shift_inst.PI_CTRL.integrator_1_17\
        );

    \I__1775\ : InMux
    port map (
            O => \N__19757\,
            I => \bfn_1_15_0_\
        );

    \I__1774\ : CascadeMux
    port map (
            O => \N__19754\,
            I => \N__19751\
        );

    \I__1773\ : InMux
    port map (
            O => \N__19751\,
            I => \N__19748\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__19748\,
            I => \N__19745\
        );

    \I__1771\ : Span4Mux_v
    port map (
            O => \N__19745\,
            I => \N__19742\
        );

    \I__1770\ : Odrv4
    port map (
            O => \N__19742\,
            I => \current_shift_inst.PI_CTRL.integrator_1_18\
        );

    \I__1769\ : InMux
    port map (
            O => \N__19739\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\
        );

    \I__1768\ : CascadeMux
    port map (
            O => \N__19736\,
            I => \N__19733\
        );

    \I__1767\ : InMux
    port map (
            O => \N__19733\,
            I => \N__19730\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__19730\,
            I => \N__19727\
        );

    \I__1765\ : Span4Mux_v
    port map (
            O => \N__19727\,
            I => \N__19724\
        );

    \I__1764\ : Odrv4
    port map (
            O => \N__19724\,
            I => \current_shift_inst.PI_CTRL.integrator_1_2\
        );

    \I__1763\ : InMux
    port map (
            O => \N__19721\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\
        );

    \I__1762\ : InMux
    port map (
            O => \N__19718\,
            I => \N__19715\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__19715\,
            I => \N__19712\
        );

    \I__1760\ : Odrv4
    port map (
            O => \N__19712\,
            I => \current_shift_inst.PI_CTRL.integrator_1_3\
        );

    \I__1759\ : InMux
    port map (
            O => \N__19709\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\
        );

    \I__1758\ : CascadeMux
    port map (
            O => \N__19706\,
            I => \N__19703\
        );

    \I__1757\ : InMux
    port map (
            O => \N__19703\,
            I => \N__19700\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__19700\,
            I => \N__19697\
        );

    \I__1755\ : Odrv4
    port map (
            O => \N__19697\,
            I => \current_shift_inst.PI_CTRL.integrator_1_4\
        );

    \I__1754\ : InMux
    port map (
            O => \N__19694\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\
        );

    \I__1753\ : CascadeMux
    port map (
            O => \N__19691\,
            I => \N__19688\
        );

    \I__1752\ : InMux
    port map (
            O => \N__19688\,
            I => \N__19685\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__19685\,
            I => \N__19682\
        );

    \I__1750\ : Span4Mux_h
    port map (
            O => \N__19682\,
            I => \N__19679\
        );

    \I__1749\ : Odrv4
    port map (
            O => \N__19679\,
            I => \current_shift_inst.PI_CTRL.integrator_1_5\
        );

    \I__1748\ : InMux
    port map (
            O => \N__19676\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\
        );

    \I__1747\ : CascadeMux
    port map (
            O => \N__19673\,
            I => \N__19670\
        );

    \I__1746\ : InMux
    port map (
            O => \N__19670\,
            I => \N__19667\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__19667\,
            I => \N__19664\
        );

    \I__1744\ : Odrv4
    port map (
            O => \N__19664\,
            I => \current_shift_inst.PI_CTRL.integrator_1_6\
        );

    \I__1743\ : InMux
    port map (
            O => \N__19661\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\
        );

    \I__1742\ : CascadeMux
    port map (
            O => \N__19658\,
            I => \N__19655\
        );

    \I__1741\ : InMux
    port map (
            O => \N__19655\,
            I => \N__19652\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__19652\,
            I => \N__19649\
        );

    \I__1739\ : Span4Mux_v
    port map (
            O => \N__19649\,
            I => \N__19646\
        );

    \I__1738\ : Odrv4
    port map (
            O => \N__19646\,
            I => \current_shift_inst.PI_CTRL.integrator_1_7\
        );

    \I__1737\ : InMux
    port map (
            O => \N__19643\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\
        );

    \I__1736\ : CascadeMux
    port map (
            O => \N__19640\,
            I => \N__19637\
        );

    \I__1735\ : InMux
    port map (
            O => \N__19637\,
            I => \N__19634\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__19634\,
            I => \N__19631\
        );

    \I__1733\ : Span4Mux_v
    port map (
            O => \N__19631\,
            I => \N__19628\
        );

    \I__1732\ : Odrv4
    port map (
            O => \N__19628\,
            I => \current_shift_inst.PI_CTRL.integrator_1_8\
        );

    \I__1731\ : InMux
    port map (
            O => \N__19625\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\
        );

    \I__1730\ : CascadeMux
    port map (
            O => \N__19622\,
            I => \N__19619\
        );

    \I__1729\ : InMux
    port map (
            O => \N__19619\,
            I => \N__19616\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__19616\,
            I => \N__19613\
        );

    \I__1727\ : Span4Mux_v
    port map (
            O => \N__19613\,
            I => \N__19610\
        );

    \I__1726\ : Odrv4
    port map (
            O => \N__19610\,
            I => \current_shift_inst.PI_CTRL.integrator_1_9\
        );

    \I__1725\ : InMux
    port map (
            O => \N__19607\,
            I => \bfn_1_14_0_\
        );

    \I__1724\ : CascadeMux
    port map (
            O => \N__19604\,
            I => \N__19601\
        );

    \I__1723\ : InMux
    port map (
            O => \N__19601\,
            I => \N__19598\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__19598\,
            I => \N__19595\
        );

    \I__1721\ : Span4Mux_v
    port map (
            O => \N__19595\,
            I => \N__19592\
        );

    \I__1720\ : Odrv4
    port map (
            O => \N__19592\,
            I => \current_shift_inst.PI_CTRL.integrator_1_10\
        );

    \I__1719\ : InMux
    port map (
            O => \N__19589\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\
        );

    \I__1718\ : InMux
    port map (
            O => \N__19586\,
            I => \N__19583\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__19583\,
            I => \N__19580\
        );

    \I__1716\ : Span4Mux_v
    port map (
            O => \N__19580\,
            I => \N__19577\
        );

    \I__1715\ : Odrv4
    port map (
            O => \N__19577\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_9\
        );

    \I__1714\ : InMux
    port map (
            O => \N__19574\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\
        );

    \I__1713\ : InMux
    port map (
            O => \N__19571\,
            I => \N__19568\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__19568\,
            I => \N__19565\
        );

    \I__1711\ : Span4Mux_v
    port map (
            O => \N__19565\,
            I => \N__19562\
        );

    \I__1710\ : Odrv4
    port map (
            O => \N__19562\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_10\
        );

    \I__1709\ : InMux
    port map (
            O => \N__19559\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\
        );

    \I__1708\ : InMux
    port map (
            O => \N__19556\,
            I => \N__19553\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__19553\,
            I => \N__19550\
        );

    \I__1706\ : Span4Mux_v
    port map (
            O => \N__19550\,
            I => \N__19547\
        );

    \I__1705\ : Odrv4
    port map (
            O => \N__19547\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_11\
        );

    \I__1704\ : InMux
    port map (
            O => \N__19544\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\
        );

    \I__1703\ : InMux
    port map (
            O => \N__19541\,
            I => \N__19538\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__19538\,
            I => \N__19535\
        );

    \I__1701\ : Span4Mux_h
    port map (
            O => \N__19535\,
            I => \N__19532\
        );

    \I__1700\ : Span4Mux_v
    port map (
            O => \N__19532\,
            I => \N__19529\
        );

    \I__1699\ : Odrv4
    port map (
            O => \N__19529\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_12\
        );

    \I__1698\ : InMux
    port map (
            O => \N__19526\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\
        );

    \I__1697\ : InMux
    port map (
            O => \N__19523\,
            I => \N__19520\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__19520\,
            I => \N__19517\
        );

    \I__1695\ : Span4Mux_v
    port map (
            O => \N__19517\,
            I => \N__19514\
        );

    \I__1694\ : Span4Mux_s1_h
    port map (
            O => \N__19514\,
            I => \N__19511\
        );

    \I__1693\ : Odrv4
    port map (
            O => \N__19511\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_13\
        );

    \I__1692\ : InMux
    port map (
            O => \N__19508\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\
        );

    \I__1691\ : InMux
    port map (
            O => \N__19505\,
            I => \N__19502\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__19502\,
            I => \N__19499\
        );

    \I__1689\ : Span4Mux_v
    port map (
            O => \N__19499\,
            I => \N__19496\
        );

    \I__1688\ : Odrv4
    port map (
            O => \N__19496\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_14\
        );

    \I__1687\ : InMux
    port map (
            O => \N__19493\,
            I => \N__19479\
        );

    \I__1686\ : CascadeMux
    port map (
            O => \N__19492\,
            I => \N__19476\
        );

    \I__1685\ : CascadeMux
    port map (
            O => \N__19491\,
            I => \N__19473\
        );

    \I__1684\ : CascadeMux
    port map (
            O => \N__19490\,
            I => \N__19470\
        );

    \I__1683\ : CascadeMux
    port map (
            O => \N__19489\,
            I => \N__19467\
        );

    \I__1682\ : CascadeMux
    port map (
            O => \N__19488\,
            I => \N__19464\
        );

    \I__1681\ : CascadeMux
    port map (
            O => \N__19487\,
            I => \N__19461\
        );

    \I__1680\ : CascadeMux
    port map (
            O => \N__19486\,
            I => \N__19458\
        );

    \I__1679\ : CascadeMux
    port map (
            O => \N__19485\,
            I => \N__19455\
        );

    \I__1678\ : CascadeMux
    port map (
            O => \N__19484\,
            I => \N__19452\
        );

    \I__1677\ : CascadeMux
    port map (
            O => \N__19483\,
            I => \N__19449\
        );

    \I__1676\ : CascadeMux
    port map (
            O => \N__19482\,
            I => \N__19446\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__19479\,
            I => \N__19443\
        );

    \I__1674\ : InMux
    port map (
            O => \N__19476\,
            I => \N__19436\
        );

    \I__1673\ : InMux
    port map (
            O => \N__19473\,
            I => \N__19436\
        );

    \I__1672\ : InMux
    port map (
            O => \N__19470\,
            I => \N__19436\
        );

    \I__1671\ : InMux
    port map (
            O => \N__19467\,
            I => \N__19427\
        );

    \I__1670\ : InMux
    port map (
            O => \N__19464\,
            I => \N__19427\
        );

    \I__1669\ : InMux
    port map (
            O => \N__19461\,
            I => \N__19427\
        );

    \I__1668\ : InMux
    port map (
            O => \N__19458\,
            I => \N__19427\
        );

    \I__1667\ : InMux
    port map (
            O => \N__19455\,
            I => \N__19422\
        );

    \I__1666\ : InMux
    port map (
            O => \N__19452\,
            I => \N__19422\
        );

    \I__1665\ : InMux
    port map (
            O => \N__19449\,
            I => \N__19417\
        );

    \I__1664\ : InMux
    port map (
            O => \N__19446\,
            I => \N__19417\
        );

    \I__1663\ : Odrv4
    port map (
            O => \N__19443\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_19\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__19436\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_19\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__19427\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_19\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__19422\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_19\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__19417\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_19\
        );

    \I__1658\ : InMux
    port map (
            O => \N__19406\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\
        );

    \I__1657\ : InMux
    port map (
            O => \N__19403\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\
        );

    \I__1656\ : InMux
    port map (
            O => \N__19400\,
            I => \N__19397\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__19397\,
            I => \N__19394\
        );

    \I__1654\ : Span4Mux_v
    port map (
            O => \N__19394\,
            I => \N__19391\
        );

    \I__1653\ : Odrv4
    port map (
            O => \N__19391\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_1\
        );

    \I__1652\ : CascadeMux
    port map (
            O => \N__19388\,
            I => \N__19385\
        );

    \I__1651\ : InMux
    port map (
            O => \N__19385\,
            I => \N__19382\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__19382\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_16\
        );

    \I__1649\ : InMux
    port map (
            O => \N__19379\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\
        );

    \I__1648\ : InMux
    port map (
            O => \N__19376\,
            I => \N__19373\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__19373\,
            I => \N__19370\
        );

    \I__1646\ : Span4Mux_v
    port map (
            O => \N__19370\,
            I => \N__19367\
        );

    \I__1645\ : Odrv4
    port map (
            O => \N__19367\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_2\
        );

    \I__1644\ : CascadeMux
    port map (
            O => \N__19364\,
            I => \N__19361\
        );

    \I__1643\ : InMux
    port map (
            O => \N__19361\,
            I => \N__19358\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__19358\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_17\
        );

    \I__1641\ : InMux
    port map (
            O => \N__19355\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\
        );

    \I__1640\ : InMux
    port map (
            O => \N__19352\,
            I => \N__19349\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__19349\,
            I => \N__19346\
        );

    \I__1638\ : Span4Mux_v
    port map (
            O => \N__19346\,
            I => \N__19343\
        );

    \I__1637\ : Odrv4
    port map (
            O => \N__19343\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_3\
        );

    \I__1636\ : CascadeMux
    port map (
            O => \N__19340\,
            I => \N__19337\
        );

    \I__1635\ : InMux
    port map (
            O => \N__19337\,
            I => \N__19334\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__19334\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_18\
        );

    \I__1633\ : InMux
    port map (
            O => \N__19331\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\
        );

    \I__1632\ : InMux
    port map (
            O => \N__19328\,
            I => \N__19325\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__19325\,
            I => \N__19322\
        );

    \I__1630\ : Span4Mux_v
    port map (
            O => \N__19322\,
            I => \N__19319\
        );

    \I__1629\ : Odrv4
    port map (
            O => \N__19319\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_4\
        );

    \I__1628\ : InMux
    port map (
            O => \N__19316\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\
        );

    \I__1627\ : InMux
    port map (
            O => \N__19313\,
            I => \N__19310\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__19310\,
            I => \N__19307\
        );

    \I__1625\ : Span4Mux_v
    port map (
            O => \N__19307\,
            I => \N__19304\
        );

    \I__1624\ : Odrv4
    port map (
            O => \N__19304\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_5\
        );

    \I__1623\ : InMux
    port map (
            O => \N__19301\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\
        );

    \I__1622\ : InMux
    port map (
            O => \N__19298\,
            I => \N__19295\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__19295\,
            I => \N__19292\
        );

    \I__1620\ : Span4Mux_v
    port map (
            O => \N__19292\,
            I => \N__19289\
        );

    \I__1619\ : Odrv4
    port map (
            O => \N__19289\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_6\
        );

    \I__1618\ : InMux
    port map (
            O => \N__19286\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\
        );

    \I__1617\ : InMux
    port map (
            O => \N__19283\,
            I => \N__19280\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__19280\,
            I => \N__19277\
        );

    \I__1615\ : Span4Mux_v
    port map (
            O => \N__19277\,
            I => \N__19274\
        );

    \I__1614\ : Odrv4
    port map (
            O => \N__19274\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_7\
        );

    \I__1613\ : InMux
    port map (
            O => \N__19271\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\
        );

    \I__1612\ : InMux
    port map (
            O => \N__19268\,
            I => \N__19265\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__19265\,
            I => \N__19262\
        );

    \I__1610\ : Span4Mux_v
    port map (
            O => \N__19262\,
            I => \N__19259\
        );

    \I__1609\ : Odrv4
    port map (
            O => \N__19259\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_8\
        );

    \I__1608\ : InMux
    port map (
            O => \N__19256\,
            I => \bfn_1_12_0_\
        );

    \I__1607\ : InMux
    port map (
            O => \N__19253\,
            I => \N__19250\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__19250\,
            I => \N__19247\
        );

    \I__1605\ : Span4Mux_v
    port map (
            O => \N__19247\,
            I => \N__19244\
        );

    \I__1604\ : Odrv4
    port map (
            O => \N__19244\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_15\
        );

    \I__1603\ : InMux
    port map (
            O => \N__19241\,
            I => \N__19238\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__19238\,
            I => \N__19235\
        );

    \I__1601\ : Span4Mux_v
    port map (
            O => \N__19235\,
            I => \N__19232\
        );

    \I__1600\ : Odrv4
    port map (
            O => \N__19232\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_0\
        );

    \I__1599\ : CascadeMux
    port map (
            O => \N__19229\,
            I => \N__19226\
        );

    \I__1598\ : InMux
    port map (
            O => \N__19226\,
            I => \N__19223\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__19223\,
            I => \N__19220\
        );

    \I__1596\ : Odrv4
    port map (
            O => \N__19220\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_15\
        );

    \I__1595\ : IoInMux
    port map (
            O => \N__19217\,
            I => \N__19214\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__19214\,
            I => \N__19211\
        );

    \I__1593\ : Span4Mux_s3_v
    port map (
            O => \N__19211\,
            I => \N__19208\
        );

    \I__1592\ : Span4Mux_h
    port map (
            O => \N__19208\,
            I => \N__19205\
        );

    \I__1591\ : Sp12to4
    port map (
            O => \N__19205\,
            I => \N__19202\
        );

    \I__1590\ : Span12Mux_v
    port map (
            O => \N__19202\,
            I => \N__19199\
        );

    \I__1589\ : Span12Mux_v
    port map (
            O => \N__19199\,
            I => \N__19196\
        );

    \I__1588\ : Odrv12
    port map (
            O => \N__19196\,
            I => delay_tr_input_ibuf_gb_io_gb_input
        );

    \I__1587\ : IoInMux
    port map (
            O => \N__19193\,
            I => \N__19190\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__19190\,
            I => \N__19187\
        );

    \I__1585\ : IoSpan4Mux
    port map (
            O => \N__19187\,
            I => \N__19184\
        );

    \I__1584\ : IoSpan4Mux
    port map (
            O => \N__19184\,
            I => \N__19181\
        );

    \I__1583\ : Odrv4
    port map (
            O => \N__19181\,
            I => delay_hc_input_ibuf_gb_io_gb_input
        );

    \IN_MUX_bfv_9_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_26_0_\
        );

    \IN_MUX_bfv_9_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_cry_7\,
            carryinitout => \bfn_9_27_0_\
        );

    \IN_MUX_bfv_9_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_cry_15\,
            carryinitout => \bfn_9_28_0_\
        );

    \IN_MUX_bfv_8_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_11_0_\
        );

    \IN_MUX_bfv_8_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_8_12_0_\
        );

    \IN_MUX_bfv_8_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_8_13_0_\
        );

    \IN_MUX_bfv_8_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_8_14_0_\
        );

    \IN_MUX_bfv_14_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_11_0_\
        );

    \IN_MUX_bfv_14_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_14_12_0_\
        );

    \IN_MUX_bfv_14_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_14_13_0_\
        );

    \IN_MUX_bfv_14_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_14_14_0_\
        );

    \IN_MUX_bfv_12_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_7_0_\
        );

    \IN_MUX_bfv_12_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_12_8_0_\
        );

    \IN_MUX_bfv_12_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_12_9_0_\
        );

    \IN_MUX_bfv_12_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_12_10_0_\
        );

    \IN_MUX_bfv_18_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_11_0_\
        );

    \IN_MUX_bfv_18_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_18_12_0_\
        );

    \IN_MUX_bfv_18_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_18_13_0_\
        );

    \IN_MUX_bfv_18_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_18_14_0_\
        );

    \IN_MUX_bfv_14_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_15_0_\
        );

    \IN_MUX_bfv_14_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s1\,
            carryinitout => \bfn_14_16_0_\
        );

    \IN_MUX_bfv_14_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s1\,
            carryinitout => \bfn_14_17_0_\
        );

    \IN_MUX_bfv_14_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s1\,
            carryinitout => \bfn_14_18_0_\
        );

    \IN_MUX_bfv_12_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_16_0_\
        );

    \IN_MUX_bfv_12_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s0\,
            carryinitout => \bfn_12_17_0_\
        );

    \IN_MUX_bfv_12_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s0\,
            carryinitout => \bfn_12_18_0_\
        );

    \IN_MUX_bfv_12_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s0\,
            carryinitout => \bfn_12_19_0_\
        );

    \IN_MUX_bfv_17_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_20_0_\
        );

    \IN_MUX_bfv_17_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_7\,
            carryinitout => \bfn_17_21_0_\
        );

    \IN_MUX_bfv_17_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_15\,
            carryinitout => \bfn_17_22_0_\
        );

    \IN_MUX_bfv_17_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_23\,
            carryinitout => \bfn_17_23_0_\
        );

    \IN_MUX_bfv_1_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_13_0_\
        );

    \IN_MUX_bfv_1_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            carryinitout => \bfn_1_14_0_\
        );

    \IN_MUX_bfv_1_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            carryinitout => \bfn_1_15_0_\
        );

    \IN_MUX_bfv_1_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            carryinitout => \bfn_1_16_0_\
        );

    \IN_MUX_bfv_4_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_17_0_\
        );

    \IN_MUX_bfv_4_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            carryinitout => \bfn_4_18_0_\
        );

    \IN_MUX_bfv_4_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            carryinitout => \bfn_4_19_0_\
        );

    \IN_MUX_bfv_4_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            carryinitout => \bfn_4_20_0_\
        );

    \IN_MUX_bfv_10_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_26_0_\
        );

    \IN_MUX_bfv_10_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_add_1_cry_7\,
            carryinitout => \bfn_10_27_0_\
        );

    \IN_MUX_bfv_10_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_add_1_cry_15\,
            carryinitout => \bfn_10_28_0_\
        );

    \IN_MUX_bfv_3_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_23_0_\
        );

    \IN_MUX_bfv_3_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un19_threshold_cry_7\,
            carryinitout => \bfn_3_24_0_\
        );

    \IN_MUX_bfv_1_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_24_0_\
        );

    \IN_MUX_bfv_1_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_1_cry_7\,
            carryinitout => \bfn_1_25_0_\
        );

    \IN_MUX_bfv_1_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_1_cry_15\,
            carryinitout => \bfn_1_26_0_\
        );

    \IN_MUX_bfv_5_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_23_0_\
        );

    \IN_MUX_bfv_5_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un14_counter_cry_7\,
            carryinitout => \bfn_5_24_0_\
        );

    \IN_MUX_bfv_5_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_26_0_\
        );

    \IN_MUX_bfv_5_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.counter_cry_7\,
            carryinitout => \bfn_5_27_0_\
        );

    \IN_MUX_bfv_9_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_12_0_\
        );

    \IN_MUX_bfv_9_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un4_running_cry_8\,
            carryinitout => \bfn_9_13_0_\
        );

    \IN_MUX_bfv_9_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un4_running_cry_16\,
            carryinitout => \bfn_9_14_0_\
        );

    \IN_MUX_bfv_15_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_13_0_\
        );

    \IN_MUX_bfv_15_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un4_running_cry_8\,
            carryinitout => \bfn_15_14_0_\
        );

    \IN_MUX_bfv_15_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un4_running_cry_16\,
            carryinitout => \bfn_15_15_0_\
        );

    \IN_MUX_bfv_11_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_8_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un4_running_cry_8\,
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_11_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un4_running_cry_16\,
            carryinitout => \bfn_11_10_0_\
        );

    \IN_MUX_bfv_17_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_10_0_\
        );

    \IN_MUX_bfv_17_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un4_running_cry_8\,
            carryinitout => \bfn_17_11_0_\
        );

    \IN_MUX_bfv_17_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un4_running_cry_16\,
            carryinitout => \bfn_17_12_0_\
        );

    \IN_MUX_bfv_8_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_7_0_\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_8_8_0_\
        );

    \IN_MUX_bfv_8_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_8_9_0_\
        );

    \IN_MUX_bfv_8_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_8_10_0_\
        );

    \IN_MUX_bfv_7_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_7_0_\
        );

    \IN_MUX_bfv_7_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            carryinitout => \bfn_7_8_0_\
        );

    \IN_MUX_bfv_7_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            carryinitout => \bfn_7_9_0_\
        );

    \IN_MUX_bfv_7_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            carryinitout => \bfn_7_10_0_\
        );

    \IN_MUX_bfv_16_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_9_0_\
        );

    \IN_MUX_bfv_16_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_16_10_0_\
        );

    \IN_MUX_bfv_16_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_16_11_0_\
        );

    \IN_MUX_bfv_16_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_16_12_0_\
        );

    \IN_MUX_bfv_16_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_5_0_\
        );

    \IN_MUX_bfv_16_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            carryinitout => \bfn_16_6_0_\
        );

    \IN_MUX_bfv_16_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            carryinitout => \bfn_16_7_0_\
        );

    \IN_MUX_bfv_16_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            carryinitout => \bfn_16_8_0_\
        );

    \IN_MUX_bfv_11_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_15_0_\
        );

    \IN_MUX_bfv_11_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_7\,
            carryinitout => \bfn_11_16_0_\
        );

    \IN_MUX_bfv_11_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_15\,
            carryinitout => \bfn_11_17_0_\
        );

    \IN_MUX_bfv_11_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_23\,
            carryinitout => \bfn_11_18_0_\
        );

    \IN_MUX_bfv_16_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_19_0_\
        );

    \IN_MUX_bfv_16_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_16_20_0_\
        );

    \IN_MUX_bfv_16_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_16_21_0_\
        );

    \IN_MUX_bfv_16_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_16_22_0_\
        );

    \IN_MUX_bfv_16_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_15_0_\
        );

    \IN_MUX_bfv_16_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_8\,
            carryinitout => \bfn_16_16_0_\
        );

    \IN_MUX_bfv_16_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_16\,
            carryinitout => \bfn_16_17_0_\
        );

    \IN_MUX_bfv_16_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_24\,
            carryinitout => \bfn_16_18_0_\
        );

    \IN_MUX_bfv_18_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_17_0_\
        );

    \IN_MUX_bfv_18_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_7\,
            carryinitout => \bfn_18_18_0_\
        );

    \IN_MUX_bfv_18_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_15\,
            carryinitout => \bfn_18_19_0_\
        );

    \IN_MUX_bfv_18_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_23\,
            carryinitout => \bfn_18_20_0_\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_11_0_\
        );

    \IN_MUX_bfv_1_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\,
            carryinitout => \bfn_1_12_0_\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_15_0_\
        );

    \IN_MUX_bfv_9_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            carryinitout => \bfn_9_16_0_\
        );

    \IN_MUX_bfv_9_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_15\,
            carryinitout => \bfn_9_17_0_\
        );

    \IN_MUX_bfv_9_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_23\,
            carryinitout => \bfn_9_18_0_\
        );

    \delay_tr_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__19217\,
            GLOBALBUFFEROUTPUT => delay_tr_input_c_g
        );

    \delay_hc_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__19193\,
            GLOBALBUFFEROUTPUT => delay_hc_input_c_g
        );

    \current_shift_inst.timer_s1.running_RNII51H_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__35558\,
            GLOBALBUFFEROUTPUT => \current_shift_inst.timer_s1.N_162_i_g\
        );

    \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__31541\,
            GLOBALBUFFEROUTPUT => \phase_controller_inst2.stoper_tr.un1_start_g\
        );

    \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__36230\,
            GLOBALBUFFEROUTPUT => \phase_controller_inst2.stoper_hc.un1_start_g\
        );

    \osc\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b10"
        )
    port map (
            CLKHFPU => \N__48437\,
            CLKHFEN => \N__48439\,
            CLKHF => clk_12mhz
        );

    \rgb_drv\ : SB_RGBA_DRV
    generic map (
            RGB2_CURRENT => "0b111111",
            CURRENT_MODE => "0b0",
            RGB0_CURRENT => "0b111111",
            RGB1_CURRENT => "0b111111"
        )
    port map (
            RGBLEDEN => \N__48438\,
            RGB2PWM => \N__24452\,
            RGB1 => rgb_g_wire,
            CURREN => \N__48404\,
            RGB2 => rgb_b_wire,
            RGB1PWM => \N__20864\,
            RGB0PWM => \N__49574\,
            RGB0 => rgb_r_wire
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19253\,
            in2 => \_gnd_net_\,
            in3 => \N__19493\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19241\,
            in2 => \N__19229\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_16\,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19400\,
            in2 => \N__19388\,
            in3 => \N__19379\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19376\,
            in2 => \N__19364\,
            in3 => \N__19355\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19352\,
            in2 => \N__19340\,
            in3 => \N__19331\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19328\,
            in2 => \N__19482\,
            in3 => \N__19316\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19313\,
            in2 => \N__19484\,
            in3 => \N__19301\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19298\,
            in2 => \N__19483\,
            in3 => \N__19286\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19283\,
            in2 => \N__19485\,
            in3 => \N__19271\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19268\,
            in2 => \N__19486\,
            in3 => \N__19256\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_24\,
            ltout => OPEN,
            carryin => \bfn_1_12_0_\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19586\,
            in2 => \N__19490\,
            in3 => \N__19574\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19571\,
            in2 => \N__19487\,
            in3 => \N__19559\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19556\,
            in2 => \N__19491\,
            in3 => \N__19544\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19541\,
            in2 => \N__19488\,
            in3 => \N__19526\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19523\,
            in2 => \N__19492\,
            in3 => \N__19508\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19505\,
            in2 => \N__19489\,
            in3 => \N__19406\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19403\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21856\,
            in2 => \N__20797\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_13_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21789\,
            in2 => \N__19736\,
            in3 => \N__19721\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19718\,
            in2 => \N__21720\,
            in3 => \N__19709\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21638\,
            in2 => \N__19706\,
            in3 => \N__19694\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21576\,
            in2 => \N__19691\,
            in3 => \N__19676\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21486\,
            in2 => \N__19673\,
            in3 => \N__19661\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23345\,
            in2 => \N__19658\,
            in3 => \N__19643\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22256\,
            in2 => \N__19640\,
            in3 => \N__19625\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22194\,
            in2 => \N__19622\,
            in3 => \N__19607\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_1_14_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22077\,
            in2 => \N__19604\,
            in3 => \N__19589\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22032\,
            in2 => \N__19868\,
            in3 => \N__19856\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21980\,
            in2 => \N__19853\,
            in3 => \N__19841\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21918\,
            in2 => \N__19838\,
            in3 => \N__19823\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22760\,
            in2 => \N__19820\,
            in3 => \N__19808\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22694\,
            in2 => \N__19805\,
            in3 => \N__19790\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22660\,
            in2 => \N__19787\,
            in3 => \N__19775\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22608\,
            in2 => \N__19772\,
            in3 => \N__19757\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_1_15_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22542\,
            in2 => \N__19754\,
            in3 => \N__19739\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20021\,
            in2 => \N__22495\,
            in3 => \N__20009\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20006\,
            in2 => \N__22435\,
            in3 => \N__19997\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22367\,
            in2 => \N__19994\,
            in3 => \N__19979\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23168\,
            in2 => \N__19976\,
            in3 => \N__19961\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23111\,
            in2 => \N__19958\,
            in3 => \N__19943\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23060\,
            in2 => \N__19940\,
            in3 => \N__19925\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23010\,
            in2 => \N__19922\,
            in3 => \N__19907\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\,
            ltout => OPEN,
            carryin => \bfn_1_16_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22962\,
            in2 => \N__19904\,
            in3 => \N__19889\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22911\,
            in2 => \N__19886\,
            in3 => \N__19871\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22863\,
            in2 => \N__20120\,
            in3 => \N__20105\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22819\,
            in2 => \N__20102\,
            in3 => \N__20090\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23289\,
            in2 => \N__20087\,
            in3 => \N__20072\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20069\,
            in1 => \N__23762\,
            in2 => \N__20057\,
            in3 => \N__20045\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24242\,
            in2 => \_gnd_net_\,
            in3 => \N__21855\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50267\,
            ce => 'H',
            sr => \N__49536\
        );

    \current_shift_inst.PI_CTRL.integrator_27_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000100010"
        )
    port map (
            in0 => \N__23836\,
            in1 => \N__23704\,
            in2 => \N__23513\,
            in3 => \N__20042\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50267\,
            ce => 'H',
            sr => \N__49536\
        );

    \current_shift_inst.PI_CTRL.integrator_26_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010111100000"
        )
    port map (
            in0 => \N__23703\,
            in1 => \N__23476\,
            in2 => \N__20036\,
            in3 => \N__23838\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50267\,
            ce => 'H',
            sr => \N__49536\
        );

    \current_shift_inst.PI_CTRL.integrator_31_LC_1_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000100010"
        )
    port map (
            in0 => \N__23837\,
            in1 => \N__23705\,
            in2 => \N__23514\,
            in3 => \N__20027\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50267\,
            ce => 'H',
            sr => \N__49536\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_1_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21442\,
            in2 => \_gnd_net_\,
            in3 => \N__22153\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_1_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21523\,
            in1 => \N__22234\,
            in2 => \N__20144\,
            in3 => \N__22309\,
            lcout => \current_shift_inst.PI_CTRL.N_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_1_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21605\,
            in2 => \_gnd_net_\,
            in3 => \N__21690\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_98_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_1_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__20185\,
            in1 => \N__28452\,
            in2 => \N__20141\,
            in3 => \N__21059\,
            lcout => \current_shift_inst.PI_CTRL.N_96\,
            ltout => \current_shift_inst.PI_CTRL.N_96_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_1_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__21691\,
            in1 => \N__20135\,
            in2 => \N__20138\,
            in3 => \N__20203\,
            lcout => \current_shift_inst.PI_CTRL.N_161\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_1_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010001"
        )
    port map (
            in0 => \N__20638\,
            in1 => \N__21607\,
            in2 => \N__20609\,
            in3 => \N__28451\,
            lcout => \current_shift_inst.PI_CTRL.N_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_1_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010101"
        )
    port map (
            in0 => \N__28453\,
            in1 => \N__21606\,
            in2 => \N__20608\,
            in3 => \N__20639\,
            lcout => \current_shift_inst.PI_CTRL.N_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_1_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__20637\,
            in1 => \N__28450\,
            in2 => \_gnd_net_\,
            in3 => \N__20601\,
            lcout => \current_shift_inst.PI_CTRL.N_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_1_LC_1_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__20167\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20129\,
            lcout => pwm_duty_input_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50212\,
            ce => 'H',
            sr => \N__49548\
        );

    \current_shift_inst.PI_CTRL.control_out_2_LC_1_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21764\,
            in2 => \_gnd_net_\,
            in3 => \N__20168\,
            lcout => pwm_duty_input_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50212\,
            ce => 'H',
            sr => \N__49548\
        );

    \current_shift_inst.PI_CTRL.control_out_9_LC_1_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101100110000"
        )
    port map (
            in0 => \N__21061\,
            in1 => \N__28465\,
            in2 => \N__20654\,
            in3 => \N__22154\,
            lcout => pwm_duty_input_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50212\,
            ce => 'H',
            sr => \N__49548\
        );

    \current_shift_inst.PI_CTRL.control_out_3_LC_1_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__21695\,
            in1 => \N__20210\,
            in2 => \_gnd_net_\,
            in3 => \N__20204\,
            lcout => pwm_duty_input_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50212\,
            ce => 'H',
            sr => \N__49548\
        );

    \current_shift_inst.PI_CTRL.control_out_5_LC_1_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111010000"
        )
    port map (
            in0 => \N__28464\,
            in1 => \N__21060\,
            in2 => \N__21530\,
            in3 => \N__20650\,
            lcout => pwm_duty_input_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50212\,
            ce => 'H',
            sr => \N__49548\
        );

    \current_shift_inst.PI_CTRL.control_out_4_LC_1_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011011111"
        )
    port map (
            in0 => \N__21062\,
            in1 => \N__21611\,
            in2 => \N__20192\,
            in3 => \N__20174\,
            lcout => pwm_duty_input_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50212\,
            ce => 'H',
            sr => \N__49548\
        );

    \current_shift_inst.PI_CTRL.control_out_0_LC_1_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24428\,
            in2 => \_gnd_net_\,
            in3 => \N__20166\,
            lcout => pwm_duty_input_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50212\,
            ce => 'H',
            sr => \N__49548\
        );

    \current_shift_inst.PI_CTRL.control_out_8_LC_1_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001000110010"
        )
    port map (
            in0 => \N__20651\,
            in1 => \N__28469\,
            in2 => \N__22238\,
            in3 => \N__21065\,
            lcout => pwm_duty_input_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50202\,
            ce => 'H',
            sr => \N__49551\
        );

    \current_shift_inst.PI_CTRL.control_out_6_LC_1_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111010000"
        )
    port map (
            in0 => \N__28467\,
            in1 => \N__21063\,
            in2 => \N__21449\,
            in3 => \N__20652\,
            lcout => pwm_duty_input_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50202\,
            ce => 'H',
            sr => \N__49551\
        );

    \current_shift_inst.PI_CTRL.control_out_7_LC_1_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111010000"
        )
    port map (
            in0 => \N__28468\,
            in1 => \N__21064\,
            in2 => \N__22316\,
            in3 => \N__20653\,
            lcout => pwm_duty_input_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50202\,
            ce => 'H',
            sr => \N__49551\
        );

    \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_1_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20156\,
            in1 => \N__20150\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_1_24_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_1_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20306\,
            in1 => \N__20300\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_0\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_1_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20288\,
            in2 => \_gnd_net_\,
            in3 => \N__20294\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_1\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_1_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20276\,
            in2 => \_gnd_net_\,
            in3 => \N__20282\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_2\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_1_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20264\,
            in2 => \_gnd_net_\,
            in3 => \N__20270\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_3\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_1_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20252\,
            in2 => \_gnd_net_\,
            in3 => \N__20258\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_4\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_1_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20240\,
            in2 => \_gnd_net_\,
            in3 => \N__20246\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_5\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_1_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20228\,
            in2 => \_gnd_net_\,
            in3 => \N__20234\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_6\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_1_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20216\,
            in2 => \_gnd_net_\,
            in3 => \N__20222\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_8\,
            ltout => OPEN,
            carryin => \bfn_1_25_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_1_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20342\,
            in1 => \N__20336\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_8\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_1_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23983\,
            in3 => \N__20330\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_9\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_1_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__30519\,
            in1 => \N__28393\,
            in2 => \_gnd_net_\,
            in3 => \N__20327\,
            lcout => \pwm_generator_inst.un19_threshold_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_10\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_1_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21210\,
            in2 => \_gnd_net_\,
            in3 => \N__20324\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_11\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_1_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21393\,
            in2 => \_gnd_net_\,
            in3 => \N__20321\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_12\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_1_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20880\,
            in2 => \_gnd_net_\,
            in3 => \N__20318\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_13\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_1_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20531\,
            in3 => \N__20315\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_14\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_1_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20697\,
            in2 => \_gnd_net_\,
            in3 => \N__20312\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_1_26_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_1_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20676\,
            in2 => \_gnd_net_\,
            in3 => \N__20309\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_16\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_1_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20722\,
            in2 => \_gnd_net_\,
            in3 => \N__20399\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_17\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_1_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20396\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_3_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__23699\,
            in1 => \N__20393\,
            in2 => \_gnd_net_\,
            in3 => \N__23460\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50305\,
            ce => 'H',
            sr => \N__49517\
        );

    \current_shift_inst.PI_CTRL.integrator_8_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110001000101"
        )
    port map (
            in0 => \N__23877\,
            in1 => \N__20387\,
            in2 => \N__23509\,
            in3 => \N__23700\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50305\,
            ce => 'H',
            sr => \N__49517\
        );

    \current_shift_inst.PI_CTRL.integrator_10_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010011100100"
        )
    port map (
            in0 => \N__23698\,
            in1 => \N__23878\,
            in2 => \N__20381\,
            in3 => \N__23459\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50305\,
            ce => 'H',
            sr => \N__49517\
        );

    \current_shift_inst.PI_CTRL.integrator_14_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011100010"
        )
    port map (
            in0 => \N__23849\,
            in1 => \N__23678\,
            in2 => \N__20372\,
            in3 => \N__23503\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50294\,
            ce => 'H',
            sr => \N__49522\
        );

    \current_shift_inst.PI_CTRL.integrator_15_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001100"
        )
    port map (
            in0 => \N__23502\,
            in1 => \N__23850\,
            in2 => \N__23701\,
            in3 => \N__20363\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50294\,
            ce => 'H',
            sr => \N__49522\
        );

    \current_shift_inst.PI_CTRL.integrator_20_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000100010"
        )
    port map (
            in0 => \N__23843\,
            in1 => \N__23658\,
            in2 => \N__23520\,
            in3 => \N__20357\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50281\,
            ce => 'H',
            sr => \N__49526\
        );

    \current_shift_inst.PI_CTRL.integrator_23_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010011100100"
        )
    port map (
            in0 => \N__23656\,
            in1 => \N__23848\,
            in2 => \N__20351\,
            in3 => \N__23501\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50281\,
            ce => 'H',
            sr => \N__49526\
        );

    \current_shift_inst.PI_CTRL.integrator_19_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000100010"
        )
    port map (
            in0 => \N__23842\,
            in1 => \N__23657\,
            in2 => \N__23519\,
            in3 => \N__20471\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50281\,
            ce => 'H',
            sr => \N__49526\
        );

    \current_shift_inst.PI_CTRL.integrator_21_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000100010"
        )
    port map (
            in0 => \N__23844\,
            in1 => \N__23659\,
            in2 => \N__23521\,
            in3 => \N__20465\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50281\,
            ce => 'H',
            sr => \N__49526\
        );

    \current_shift_inst.PI_CTRL.integrator_18_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010011100100"
        )
    port map (
            in0 => \N__23654\,
            in1 => \N__23846\,
            in2 => \N__20459\,
            in3 => \N__23499\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50281\,
            ce => 'H',
            sr => \N__49526\
        );

    \current_shift_inst.PI_CTRL.integrator_24_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000100010"
        )
    port map (
            in0 => \N__23845\,
            in1 => \N__23660\,
            in2 => \N__23522\,
            in3 => \N__20450\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50281\,
            ce => 'H',
            sr => \N__49526\
        );

    \current_shift_inst.PI_CTRL.integrator_22_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010011100100"
        )
    port map (
            in0 => \N__23655\,
            in1 => \N__23847\,
            in2 => \N__20444\,
            in3 => \N__23500\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50281\,
            ce => 'H',
            sr => \N__49526\
        );

    \current_shift_inst.PI_CTRL.integrator_29_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101100"
        )
    port map (
            in0 => \N__23454\,
            in1 => \N__23803\,
            in2 => \N__20435\,
            in3 => \N__23653\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50269\,
            ce => 'H',
            sr => \N__49530\
        );

    \current_shift_inst.PI_CTRL.integrator_25_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101100"
        )
    port map (
            in0 => \N__23452\,
            in1 => \N__23801\,
            in2 => \N__20426\,
            in3 => \N__23651\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50269\,
            ce => 'H',
            sr => \N__49530\
        );

    \current_shift_inst.PI_CTRL.integrator_30_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001010"
        )
    port map (
            in0 => \N__23800\,
            in1 => \N__23455\,
            in2 => \N__23689\,
            in3 => \N__20417\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50269\,
            ce => 'H',
            sr => \N__49530\
        );

    \current_shift_inst.PI_CTRL.integrator_28_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101100"
        )
    port map (
            in0 => \N__23453\,
            in1 => \N__23802\,
            in2 => \N__20411\,
            in3 => \N__23652\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50269\,
            ce => 'H',
            sr => \N__49530\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__23350\,
            in1 => \N__22276\,
            in2 => \_gnd_net_\,
            in3 => \N__21572\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_2_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__20891\,
            in1 => \N__22196\,
            in2 => \N__20507\,
            in3 => \N__21487\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_43_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20501\,
            in1 => \N__20495\,
            in2 => \N__20504\,
            in3 => \N__20660\,
            lcout => \current_shift_inst.PI_CTRL.N_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_2_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22765\,
            in1 => \N__22656\,
            in2 => \N__22039\,
            in3 => \N__21977\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22817\,
            in1 => \N__21919\,
            in2 => \N__22109\,
            in3 => \N__22705\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_2_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22612\,
            in1 => \N__22494\,
            in2 => \N__23179\,
            in3 => \N__22546\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_2_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22867\,
            in1 => \N__22907\,
            in2 => \N__23020\,
            in3 => \N__23293\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__22371\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22955\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_2_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__22430\,
            in1 => \N__23064\,
            in2 => \N__20489\,
            in3 => \N__20486\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_2_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__23116\,
            in1 => \N__23761\,
            in2 => \N__20480\,
            in3 => \N__20477\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_2_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22431\,
            in1 => \N__23065\,
            in2 => \N__22384\,
            in3 => \N__23804\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_2_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20948\,
            in1 => \N__20954\,
            in2 => \N__21008\,
            in3 => \N__21089\,
            lcout => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22149\,
            in2 => \_gnd_net_\,
            in3 => \N__21522\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__22233\,
            in1 => \N__22308\,
            in2 => \N__20612\,
            in3 => \N__21441\,
            lcout => \current_shift_inst.PI_CTRL.N_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un1_duty_inputlto2_LC_2_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__20587\,
            in1 => \N__20569\,
            in2 => \_gnd_net_\,
            in3 => \N__20554\,
            lcout => \pwm_generator_inst.un1_duty_inputlt3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_2_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23976\,
            in2 => \_gnd_net_\,
            in3 => \N__23941\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_2_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110001011100"
        )
    port map (
            in0 => \N__20537\,
            in1 => \N__28280\,
            in2 => \N__30520\,
            in3 => \N__20885\,
            lcout => \pwm_generator_inst.un19_threshold_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_2_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20530\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28255\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_15\,
            ltout => \pwm_generator_inst.un15_threshold_1_axb_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_2_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010111001100"
        )
    port map (
            in0 => \N__20516\,
            in1 => \N__28256\,
            in2 => \N__20510\,
            in3 => \N__30503\,
            lcout => \pwm_generator_inst.un19_threshold_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_2_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011011110000100"
        )
    port map (
            in0 => \N__20747\,
            in1 => \N__30502\,
            in2 => \N__20705\,
            in3 => \N__28232\,
            lcout => \pwm_generator_inst.un19_threshold_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21240\,
            in2 => \_gnd_net_\,
            in3 => \N__24109\,
            lcout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_2_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110001011100"
        )
    port map (
            in0 => \N__20738\,
            in1 => \N__28559\,
            in2 => \N__30521\,
            in3 => \N__20681\,
            lcout => \pwm_generator_inst.un19_threshold_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_2_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100001110100"
        )
    port map (
            in0 => \N__20721\,
            in1 => \N__30500\,
            in2 => \N__28535\,
            in3 => \N__20729\,
            lcout => \pwm_generator_inst.un19_threshold_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_2_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28525\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20723\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_2_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20701\,
            in2 => \_gnd_net_\,
            in3 => \N__28225\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_2_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \N__20680\,
            in1 => \N__28552\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_2_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28318\,
            in2 => \_gnd_net_\,
            in3 => \N__21397\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_2_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28357\,
            in2 => \_gnd_net_\,
            in3 => \N__21212\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_2_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28273\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20884\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_drv_RNO_LC_2_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__49573\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33560\,
            lcout => \rgb_drv_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_13_LC_3_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011100010"
        )
    port map (
            in0 => \N__23873\,
            in1 => \N__23684\,
            in2 => \N__20852\,
            in3 => \N__23516\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50295\,
            ce => 'H',
            sr => \N__49515\
        );

    \current_shift_inst.PI_CTRL.integrator_2_LC_3_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__20837\,
            in1 => \N__23685\,
            in2 => \_gnd_net_\,
            in3 => \N__23517\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50295\,
            ce => 'H',
            sr => \N__49515\
        );

    \current_shift_inst.PI_CTRL.integrator_11_LC_3_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011100010"
        )
    port map (
            in0 => \N__23872\,
            in1 => \N__23683\,
            in2 => \N__20828\,
            in3 => \N__23515\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50295\,
            ce => 'H',
            sr => \N__49515\
        );

    \current_shift_inst.PI_CTRL.integrator_5_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101000011010001"
        )
    port map (
            in0 => \N__23868\,
            in1 => \N__23682\,
            in2 => \N__20813\,
            in3 => \N__23508\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50282\,
            ce => 'H',
            sr => \N__49518\
        );

    \current_shift_inst.PI_CTRL.integrator_1_LC_3_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001011001000"
        )
    port map (
            in0 => \N__23507\,
            in1 => \N__21847\,
            in2 => \N__23702\,
            in3 => \N__20798\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50282\,
            ce => 'H',
            sr => \N__49518\
        );

    \current_shift_inst.PI_CTRL.integrator_12_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011100010"
        )
    port map (
            in0 => \N__23865\,
            in1 => \N__23646\,
            in2 => \N__20774\,
            in3 => \N__23506\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50270\,
            ce => 'H',
            sr => \N__49523\
        );

    \current_shift_inst.PI_CTRL.integrator_16_LC_3_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001100"
        )
    port map (
            in0 => \N__23504\,
            in1 => \N__23867\,
            in2 => \N__23688\,
            in3 => \N__20759\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50270\,
            ce => 'H',
            sr => \N__49523\
        );

    \current_shift_inst.PI_CTRL.integrator_17_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101010"
        )
    port map (
            in0 => \N__23866\,
            in1 => \N__23505\,
            in2 => \N__20933\,
            in3 => \N__23647\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50270\,
            ce => 'H',
            sr => \N__49523\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_3_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22487\,
            in1 => \N__22541\,
            in2 => \N__23175\,
            in3 => \N__22604\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_3_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22269\,
            in1 => \N__23349\,
            in2 => \N__22190\,
            in3 => \N__21479\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_3_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__21654\,
            in1 => \N__21578\,
            in2 => \N__20921\,
            in3 => \N__21735\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_44_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22818\,
            in1 => \N__23112\,
            in2 => \N__20918\,
            in3 => \N__20915\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_3_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20975\,
            in1 => \N__20897\,
            in2 => \N__20909\,
            in3 => \N__20906\,
            lcout => \current_shift_inst.PI_CTRL.N_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_3_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22862\,
            in1 => \N__23009\,
            in2 => \N__22925\,
            in3 => \N__22969\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000111"
        )
    port map (
            in0 => \N__21848\,
            in1 => \N__21739\,
            in2 => \N__21656\,
            in3 => \N__21793\,
            lcout => \current_shift_inst.PI_CTRL.N_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_3_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22704\,
            in1 => \N__21911\,
            in2 => \N__22105\,
            in3 => \N__22655\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_3_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21978\,
            in1 => \N__20969\,
            in2 => \N__20978\,
            in3 => \N__23288\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22764\,
            in2 => \_gnd_net_\,
            in3 => \N__22022\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22627\,
            in1 => \N__22675\,
            in2 => \N__22796\,
            in3 => \N__22060\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_3_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22628\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22676\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_3_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21946\,
            in2 => \_gnd_net_\,
            in3 => \N__22061\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22513\,
            in2 => \_gnd_net_\,
            in3 => \N__22576\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_3_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21991\,
            in1 => \N__21947\,
            in2 => \N__20963\,
            in3 => \N__20960\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23036\,
            in1 => \N__22726\,
            in2 => \N__23087\,
            in3 => \N__21874\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22343\,
            in1 => \N__23086\,
            in2 => \N__22795\,
            in3 => \N__23035\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_3_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22838\,
            in1 => \N__21992\,
            in2 => \N__20942\,
            in3 => \N__20939\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__22339\,
            in1 => \N__23137\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_3_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22885\,
            in1 => \N__22837\,
            in2 => \N__21092\,
            in3 => \N__23263\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_3_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22985\,
            in1 => \N__21083\,
            in2 => \N__23141\,
            in3 => \N__22937\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_3_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20999\,
            in1 => \N__21014\,
            in2 => \N__21074\,
            in3 => \N__21071\,
            lcout => \current_shift_inst.PI_CTRL.N_159\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_3_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22463\,
            in1 => \N__21878\,
            in2 => \N__22736\,
            in3 => \N__22402\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_3_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22936\,
            in1 => \N__22984\,
            in2 => \N__22403\,
            in3 => \N__22462\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_3_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23264\,
            in1 => \N__22577\,
            in2 => \N__22517\,
            in3 => \N__22886\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_3_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23918\,
            in2 => \N__30529\,
            in3 => \N__30525\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93\,
            ltout => OPEN,
            carryin => \bfn_3_23_0_\,
            carryout => \pwm_generator_inst.un19_threshold_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_3_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20993\,
            in2 => \_gnd_net_\,
            in3 => \N__20981\,
            lcout => \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_0\,
            carryout => \pwm_generator_inst.un19_threshold_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_3_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21194\,
            in2 => \_gnd_net_\,
            in3 => \N__21158\,
            lcout => \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_1\,
            carryout => \pwm_generator_inst.un19_threshold_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_3_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21362\,
            in2 => \_gnd_net_\,
            in3 => \N__21155\,
            lcout => \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_2\,
            carryout => \pwm_generator_inst.un19_threshold_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_3_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21152\,
            in2 => \_gnd_net_\,
            in3 => \N__21146\,
            lcout => \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_3\,
            carryout => \pwm_generator_inst.un19_threshold_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_3_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21143\,
            in2 => \_gnd_net_\,
            in3 => \N__21137\,
            lcout => \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_4\,
            carryout => \pwm_generator_inst.un19_threshold_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_3_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21134\,
            in2 => \_gnd_net_\,
            in3 => \N__21128\,
            lcout => \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_5\,
            carryout => \pwm_generator_inst.un19_threshold_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_3_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21125\,
            in2 => \_gnd_net_\,
            in3 => \N__21119\,
            lcout => \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_6\,
            carryout => \pwm_generator_inst.un19_threshold_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_3_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21116\,
            in2 => \_gnd_net_\,
            in3 => \N__21110\,
            lcout => \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033\,
            ltout => OPEN,
            carryin => \bfn_3_24_0_\,
            carryout => \pwm_generator_inst.un19_threshold_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_3_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__21107\,
            in1 => \N__28508\,
            in2 => \N__30530\,
            in3 => \N__21095\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_3_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__32424\,
            in1 => \N__24077\,
            in2 => \N__21401\,
            in3 => \N__24040\,
            lcout => \pwm_generator_inst.threshold_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_3_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__28319\,
            in1 => \N__21398\,
            in2 => \N__21377\,
            in3 => \N__30501\,
            lcout => \pwm_generator_inst.un19_threshold_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_LC_3_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101011"
        )
    port map (
            in0 => \N__21341\,
            in1 => \N__24172\,
            in2 => \N__24146\,
            in3 => \N__21356\,
            lcout => \pwm_generator_inst.N_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__21347\,
            in1 => \N__21334\,
            in2 => \N__21311\,
            in3 => \N__21277\,
            lcout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_3_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21335\,
            in1 => \N__21310\,
            in2 => \N__21281\,
            in3 => \N__21251\,
            lcout => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_3_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__21221\,
            in1 => \N__21211\,
            in2 => \N__28364\,
            in3 => \N__30499\,
            lcout => \pwm_generator_inst.un19_threshold_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_4_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011100010"
        )
    port map (
            in0 => \N__23879\,
            in1 => \N__23687\,
            in2 => \N__21185\,
            in3 => \N__23518\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50283\,
            ce => 'H',
            sr => \N__49510\
        );

    \current_shift_inst.PI_CTRL.integrator_6_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101000011010001"
        )
    port map (
            in0 => \N__23870\,
            in1 => \N__23686\,
            in2 => \N__21173\,
            in3 => \N__23511\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50271\,
            ce => 'H',
            sr => \N__49516\
        );

    \current_shift_inst.PI_CTRL.prop_term_7_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27673\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50259\,
            ce => 'H',
            sr => \N__49519\
        );

    \current_shift_inst.PI_CTRL.prop_term_4_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27295\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50259\,
            ce => 'H',
            sr => \N__49519\
        );

    \current_shift_inst.PI_CTRL.prop_term_6_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27700\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50259\,
            ce => 'H',
            sr => \N__49519\
        );

    \current_shift_inst.PI_CTRL.prop_term_2_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27352\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50259\,
            ce => 'H',
            sr => \N__49519\
        );

    \current_shift_inst.PI_CTRL.prop_term_10_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27592\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50259\,
            ce => 'H',
            sr => \N__49519\
        );

    \current_shift_inst.PI_CTRL.prop_term_13_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27497\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50259\,
            ce => 'H',
            sr => \N__49519\
        );

    \current_shift_inst.PI_CTRL.integrator_9_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000001010001"
        )
    port map (
            in0 => \N__23869\,
            in1 => \N__23510\,
            in2 => \N__21416\,
            in3 => \N__23661\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50259\,
            ce => 'H',
            sr => \N__49519\
        );

    \current_shift_inst.PI_CTRL.prop_term_3_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27328\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50247\,
            ce => 'H',
            sr => \N__49524\
        );

    \current_shift_inst.PI_CTRL.prop_term_5_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27275\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50247\,
            ce => 'H',
            sr => \N__49524\
        );

    \current_shift_inst.PI_CTRL.prop_term_22_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27733\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50247\,
            ce => 'H',
            sr => \N__49524\
        );

    \current_shift_inst.PI_CTRL.prop_term_20_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27799\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50247\,
            ce => 'H',
            sr => \N__49524\
        );

    \current_shift_inst.PI_CTRL.prop_term_11_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27550\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50247\,
            ce => 'H',
            sr => \N__49524\
        );

    \current_shift_inst.PI_CTRL.prop_term_18_LC_4_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27863\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50247\,
            ce => 'H',
            sr => \N__49524\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24238\,
            in2 => \N__21860\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_17_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_2_LC_4_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21806\,
            in2 => \N__21797\,
            in3 => \N__21749\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            clk => \N__50235\,
            ce => 'H',
            sr => \N__49527\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_3_LC_4_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21746\,
            in2 => \N__21740\,
            in3 => \N__21668\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            clk => \N__50235\,
            ce => 'H',
            sr => \N__49527\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_4_LC_4_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21665\,
            in2 => \N__21655\,
            in3 => \N__21581\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            clk => \N__50235\,
            ce => 'H',
            sr => \N__49527\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_5_LC_4_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21577\,
            in2 => \N__21539\,
            in3 => \N__21500\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            clk => \N__50235\,
            ce => 'H',
            sr => \N__49527\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_6_LC_4_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21497\,
            in2 => \N__21488\,
            in3 => \N__21419\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            clk => \N__50235\,
            ce => 'H',
            sr => \N__49527\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_7_LC_4_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22325\,
            in2 => \N__23351\,
            in3 => \N__22280\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            clk => \N__50235\,
            ce => 'H',
            sr => \N__49527\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_8_LC_4_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22277\,
            in2 => \N__24263\,
            in3 => \N__22199\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            clk => \N__50235\,
            ce => 'H',
            sr => \N__49527\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_9_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24227\,
            in2 => \N__22195\,
            in3 => \N__22121\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_4_18_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            clk => \N__50224\,
            ce => 'H',
            sr => \N__49531\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_10_LC_4_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22118\,
            in2 => \N__22104\,
            in3 => \N__22052\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            clk => \N__50224\,
            ce => 'H',
            sr => \N__49531\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_11_LC_4_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22049\,
            in2 => \N__22040\,
            in3 => \N__21983\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            clk => \N__50224\,
            ce => 'H',
            sr => \N__49531\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_12_LC_4_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21979\,
            in2 => \N__24254\,
            in3 => \N__21935\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            clk => \N__50224\,
            ce => 'H',
            sr => \N__49531\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_13_LC_4_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21932\,
            in2 => \N__21923\,
            in3 => \N__21863\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            clk => \N__50224\,
            ce => 'H',
            sr => \N__49531\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_14_LC_4_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24221\,
            in2 => \N__22772\,
            in3 => \N__22715\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            clk => \N__50224\,
            ce => 'H',
            sr => \N__49531\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_15_LC_4_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24326\,
            in2 => \N__22712\,
            in3 => \N__22667\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            clk => \N__50224\,
            ce => 'H',
            sr => \N__49531\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_16_LC_4_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24215\,
            in2 => \N__22664\,
            in3 => \N__22619\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            clk => \N__50224\,
            ce => 'H',
            sr => \N__49531\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_17_LC_4_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24296\,
            in2 => \N__22616\,
            in3 => \N__22565\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_4_19_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            clk => \N__50213\,
            ce => 'H',
            sr => \N__49534\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_18_LC_4_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22562\,
            in2 => \N__22553\,
            in3 => \N__22502\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            clk => \N__50213\,
            ce => 'H',
            sr => \N__49534\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_19_LC_4_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22499\,
            in2 => \N__24209\,
            in3 => \N__22454\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            clk => \N__50213\,
            ce => 'H',
            sr => \N__49534\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_20_LC_4_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22451\,
            in2 => \N__22442\,
            in3 => \N__22391\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            clk => \N__50213\,
            ce => 'H',
            sr => \N__49534\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_21_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24200\,
            in2 => \N__22388\,
            in3 => \N__22328\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            clk => \N__50213\,
            ce => 'H',
            sr => \N__49534\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_22_LC_4_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23192\,
            in2 => \N__23183\,
            in3 => \N__23126\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            clk => \N__50213\,
            ce => 'H',
            sr => \N__49534\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_23_LC_4_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24308\,
            in2 => \N__23123\,
            in3 => \N__23075\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            clk => \N__50213\,
            ce => 'H',
            sr => \N__49534\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_24_LC_4_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24302\,
            in2 => \N__23072\,
            in3 => \N__23027\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            clk => \N__50213\,
            ce => 'H',
            sr => \N__49534\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_25_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24275\,
            in2 => \N__23024\,
            in3 => \N__22976\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_4_20_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            clk => \N__50203\,
            ce => 'H',
            sr => \N__49537\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_26_LC_4_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24281\,
            in2 => \N__22973\,
            in3 => \N__22928\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            clk => \N__50203\,
            ce => 'H',
            sr => \N__49537\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_27_LC_4_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22924\,
            in2 => \N__24194\,
            in3 => \N__22874\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            clk => \N__50203\,
            ce => 'H',
            sr => \N__49537\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_28_LC_4_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22871\,
            in2 => \N__24320\,
            in3 => \N__22829\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            clk => \N__50203\,
            ce => 'H',
            sr => \N__49537\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_29_LC_4_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22826\,
            in2 => \N__24290\,
            in3 => \N__22775\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            clk => \N__50203\,
            ce => 'H',
            sr => \N__49537\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_30_LC_4_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24269\,
            in2 => \N__23300\,
            in3 => \N__23252\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\,
            clk => \N__50203\,
            ce => 'H',
            sr => \N__49537\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_31_LC_4_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23851\,
            in1 => \N__28478\,
            in2 => \_gnd_net_\,
            in3 => \N__23249\,
            lcout => \current_shift_inst.PI_CTRL.un8_enablelto31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50203\,
            ce => 'H',
            sr => \N__49537\
        );

    \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_4_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__24071\,
            in1 => \N__32391\,
            in2 => \N__24042\,
            in3 => \N__23246\,
            lcout => \pwm_generator_inst.threshold_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_4_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__32393\,
            in1 => \N__24073\,
            in2 => \N__23240\,
            in3 => \N__24033\,
            lcout => \pwm_generator_inst.threshold_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_4_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__24072\,
            in1 => \N__32392\,
            in2 => \N__24043\,
            in3 => \N__23231\,
            lcout => \pwm_generator_inst.threshold_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_4_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__32394\,
            in1 => \N__24074\,
            in2 => \N__23225\,
            in3 => \N__24034\,
            lcout => \pwm_generator_inst.threshold_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_4_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000111"
        )
    port map (
            in0 => \N__24075\,
            in1 => \N__32395\,
            in2 => \N__24044\,
            in3 => \N__23216\,
            lcout => \pwm_generator_inst.un14_counter_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_4_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110111"
        )
    port map (
            in0 => \N__32390\,
            in1 => \N__24070\,
            in2 => \N__23210\,
            in3 => \N__24026\,
            lcout => \pwm_generator_inst.un14_counter_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_4_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__24069\,
            in1 => \N__32389\,
            in2 => \N__24041\,
            in3 => \N__23198\,
            lcout => \pwm_generator_inst.threshold_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_4_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110111"
        )
    port map (
            in0 => \N__32396\,
            in1 => \N__24076\,
            in2 => \N__24182\,
            in3 => \N__24038\,
            lcout => \pwm_generator_inst.un14_counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_LC_4_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__24173\,
            in1 => \N__24142\,
            in2 => \N__24116\,
            in3 => \N__24083\,
            lcout => \pwm_generator_inst.N_17\,
            ltout => \pwm_generator_inst.N_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_4_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111011101"
        )
    port map (
            in0 => \N__24039\,
            in1 => \N__23993\,
            in2 => \N__23987\,
            in3 => \N__32423\,
            lcout => \pwm_generator_inst.un14_counter_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_4_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__23984\,
            in1 => \N__23954\,
            in2 => \N__23945\,
            in3 => \N__30498\,
            lcout => \pwm_generator_inst.un19_threshold_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_4_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23906\,
            lcout => \GB_BUFFER_clk_12mhz_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29074\,
            in1 => \N__29106\,
            in2 => \_gnd_net_\,
            in3 => \N__34816\,
            lcout => \elapsed_time_ns_1_RNI6HPBB_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_28_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29111\,
            in1 => \N__29070\,
            in2 => \_gnd_net_\,
            in3 => \N__34817\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50296\,
            ce => \N__29767\,
            sr => \N__49499\
        );

    \current_shift_inst.PI_CTRL.integrator_7_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101000011010001"
        )
    port map (
            in0 => \N__23871\,
            in1 => \N__23690\,
            in2 => \N__23537\,
            in3 => \N__23512\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50260\,
            ce => 'H',
            sr => \N__49511\
        );

    \current_shift_inst.PI_CTRL.prop_term_8_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27649\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50236\,
            ce => 'H',
            sr => \N__49520\
        );

    \current_shift_inst.PI_CTRL.prop_term_12_LC_5_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27520\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50236\,
            ce => 'H',
            sr => \N__49520\
        );

    \current_shift_inst.PI_CTRL.prop_term_1_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27386\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50225\,
            ce => 'H',
            sr => \N__49525\
        );

    \current_shift_inst.PI_CTRL.prop_term_9_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27622\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50225\,
            ce => 'H',
            sr => \N__49525\
        );

    \current_shift_inst.PI_CTRL.prop_term_14_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27466\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50225\,
            ce => 'H',
            sr => \N__49525\
        );

    \current_shift_inst.PI_CTRL.prop_term_16_LC_5_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27922\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50225\,
            ce => 'H',
            sr => \N__49525\
        );

    \current_shift_inst.PI_CTRL.prop_term_19_LC_5_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27826\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50214\,
            ce => 'H',
            sr => \N__49528\
        );

    \current_shift_inst.PI_CTRL.prop_term_21_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27764\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50214\,
            ce => 'H',
            sr => \N__49528\
        );

    \current_shift_inst.PI_CTRL.prop_term_27_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28075\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50214\,
            ce => 'H',
            sr => \N__49528\
        );

    \current_shift_inst.PI_CTRL.prop_term_15_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27955\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50214\,
            ce => 'H',
            sr => \N__49528\
        );

    \current_shift_inst.PI_CTRL.prop_term_28_LC_5_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28048\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50214\,
            ce => 'H',
            sr => \N__49528\
        );

    \current_shift_inst.PI_CTRL.prop_term_23_LC_5_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28201\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50214\,
            ce => 'H',
            sr => \N__49528\
        );

    \current_shift_inst.PI_CTRL.prop_term_24_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28171\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50204\,
            ce => 'H',
            sr => \N__49532\
        );

    \current_shift_inst.PI_CTRL.prop_term_17_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27892\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50204\,
            ce => 'H',
            sr => \N__49532\
        );

    \current_shift_inst.PI_CTRL.prop_term_29_LC_5_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28025\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50204\,
            ce => 'H',
            sr => \N__49532\
        );

    \current_shift_inst.PI_CTRL.prop_term_26_LC_5_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28111\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50204\,
            ce => 'H',
            sr => \N__49532\
        );

    \current_shift_inst.PI_CTRL.prop_term_25_LC_5_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28142\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50195\,
            ce => 'H',
            sr => \N__49535\
        );

    \current_shift_inst.PI_CTRL.prop_term_30_LC_5_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27991\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50195\,
            ce => 'H',
            sr => \N__49535\
        );

    \current_shift_inst.PI_CTRL.prop_term_0_LC_5_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29725\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50189\,
            ce => 'H',
            sr => \N__49538\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24434\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50185\,
            ce => 'H',
            sr => \N__49540\
        );

    \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_5_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24410\,
            in2 => \N__24419\,
            in3 => \N__24710\,
            lcout => \pwm_generator_inst.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_5_23_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_5_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24395\,
            in2 => \N__24404\,
            in3 => \N__24686\,
            lcout => \pwm_generator_inst.counter_i_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_0\,
            carryout => \pwm_generator_inst.un14_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_5_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24380\,
            in2 => \N__24389\,
            in3 => \N__24662\,
            lcout => \pwm_generator_inst.counter_i_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_1\,
            carryout => \pwm_generator_inst.un14_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_5_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24638\,
            in1 => \N__24362\,
            in2 => \N__24371\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_2\,
            carryout => \pwm_generator_inst.un14_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_5_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24356\,
            in2 => \N__24350\,
            in3 => \N__24614\,
            lcout => \pwm_generator_inst.counter_i_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_3\,
            carryout => \pwm_generator_inst.un14_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_5_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24590\,
            in1 => \N__24332\,
            in2 => \N__24341\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_4\,
            carryout => \pwm_generator_inst.un14_counter_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_5_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24533\,
            in2 => \N__24542\,
            in3 => \N__24566\,
            lcout => \pwm_generator_inst.counter_i_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_5\,
            carryout => \pwm_generator_inst.un14_counter_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_5_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24527\,
            in2 => \N__24521\,
            in3 => \N__24854\,
            lcout => \pwm_generator_inst.counter_i_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_6\,
            carryout => \pwm_generator_inst.un14_counter_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_5_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24503\,
            in2 => \N__24512\,
            in3 => \N__24830\,
            lcout => \pwm_generator_inst.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_5_24_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_5_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24485\,
            in2 => \N__24497\,
            in3 => \N__24758\,
            lcout => \pwm_generator_inst.counter_i_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_8\,
            carryout => \pwm_generator_inst.un14_counter_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.pwm_out_LC_5_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24479\,
            lcout => pwm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50180\,
            ce => 'H',
            sr => \N__49544\
        );

    \rgb_drv_RNO_0_LC_5_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__49572\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33553\,
            lcout => \N_38_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIVDL3_9_LC_5_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__24757\,
            in1 => \N__24829\,
            in2 => \_gnd_net_\,
            in3 => \N__24852\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto9_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIFA6C_5_LC_5_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__24565\,
            in1 => \N__24589\,
            in2 => \N__24437\,
            in3 => \N__24716\,
            lcout => \pwm_generator_inst.un1_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNISQD2_0_LC_5_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24705\,
            in2 => \_gnd_net_\,
            in3 => \N__24657\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIBO26_1_LC_5_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__24612\,
            in1 => \N__24684\,
            in2 => \N__24719\,
            in3 => \N__24636\,
            lcout => \pwm_generator_inst.un1_counterlt9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_0_LC_5_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24800\,
            in1 => \N__24709\,
            in2 => \_gnd_net_\,
            in3 => \N__24689\,
            lcout => \pwm_generator_inst.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_5_26_0_\,
            carryout => \pwm_generator_inst.counter_cry_0\,
            clk => \N__50176\,
            ce => 'H',
            sr => \N__49549\
        );

    \pwm_generator_inst.counter_1_LC_5_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24794\,
            in1 => \N__24685\,
            in2 => \_gnd_net_\,
            in3 => \N__24665\,
            lcout => \pwm_generator_inst.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_0\,
            carryout => \pwm_generator_inst.counter_cry_1\,
            clk => \N__50176\,
            ce => 'H',
            sr => \N__49549\
        );

    \pwm_generator_inst.counter_2_LC_5_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24801\,
            in1 => \N__24661\,
            in2 => \_gnd_net_\,
            in3 => \N__24641\,
            lcout => \pwm_generator_inst.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_1\,
            carryout => \pwm_generator_inst.counter_cry_2\,
            clk => \N__50176\,
            ce => 'H',
            sr => \N__49549\
        );

    \pwm_generator_inst.counter_3_LC_5_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24795\,
            in1 => \N__24637\,
            in2 => \_gnd_net_\,
            in3 => \N__24617\,
            lcout => \pwm_generator_inst.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_2\,
            carryout => \pwm_generator_inst.counter_cry_3\,
            clk => \N__50176\,
            ce => 'H',
            sr => \N__49549\
        );

    \pwm_generator_inst.counter_4_LC_5_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24802\,
            in1 => \N__24613\,
            in2 => \_gnd_net_\,
            in3 => \N__24593\,
            lcout => \pwm_generator_inst.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_3\,
            carryout => \pwm_generator_inst.counter_cry_4\,
            clk => \N__50176\,
            ce => 'H',
            sr => \N__49549\
        );

    \pwm_generator_inst.counter_5_LC_5_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24796\,
            in1 => \N__24588\,
            in2 => \_gnd_net_\,
            in3 => \N__24569\,
            lcout => \pwm_generator_inst.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_4\,
            carryout => \pwm_generator_inst.counter_cry_5\,
            clk => \N__50176\,
            ce => 'H',
            sr => \N__49549\
        );

    \pwm_generator_inst.counter_6_LC_5_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24803\,
            in1 => \N__24564\,
            in2 => \_gnd_net_\,
            in3 => \N__24545\,
            lcout => \pwm_generator_inst.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_5\,
            carryout => \pwm_generator_inst.counter_cry_6\,
            clk => \N__50176\,
            ce => 'H',
            sr => \N__49549\
        );

    \pwm_generator_inst.counter_7_LC_5_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24797\,
            in1 => \N__24853\,
            in2 => \_gnd_net_\,
            in3 => \N__24833\,
            lcout => \pwm_generator_inst.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_6\,
            carryout => \pwm_generator_inst.counter_cry_7\,
            clk => \N__50176\,
            ce => 'H',
            sr => \N__49549\
        );

    \pwm_generator_inst.counter_8_LC_5_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24799\,
            in1 => \N__24828\,
            in2 => \_gnd_net_\,
            in3 => \N__24806\,
            lcout => \pwm_generator_inst.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_5_27_0_\,
            carryout => \pwm_generator_inst.counter_cry_8\,
            clk => \N__50173\,
            ce => 'H',
            sr => \N__49552\
        );

    \pwm_generator_inst.counter_9_LC_5_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__24756\,
            in1 => \N__24798\,
            in2 => \_gnd_net_\,
            in3 => \N__24761\,
            lcout => \pwm_generator_inst.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50173\,
            ce => 'H',
            sr => \N__49552\
        );

    \phase_controller_inst2.stoper_tr.target_time_29_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34758\,
            in1 => \N__28907\,
            in2 => \_gnd_net_\,
            in3 => \N__28886\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50319\,
            ce => \N__29760\,
            sr => \N__49460\
        );

    \delay_measurement_inst.delay_tr_timer.counter_0_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25075\,
            in1 => \N__25485\,
            in2 => \_gnd_net_\,
            in3 => \N__24734\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_7_7_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            clk => \N__50314\,
            ce => \N__25160\,
            sr => \N__49468\
        );

    \delay_measurement_inst.delay_tr_timer.counter_1_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25067\,
            in1 => \N__25464\,
            in2 => \_gnd_net_\,
            in3 => \N__24731\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            clk => \N__50314\,
            ce => \N__25160\,
            sr => \N__49468\
        );

    \delay_measurement_inst.delay_tr_timer.counter_2_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25076\,
            in1 => \N__25441\,
            in2 => \_gnd_net_\,
            in3 => \N__24728\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            clk => \N__50314\,
            ce => \N__25160\,
            sr => \N__49468\
        );

    \delay_measurement_inst.delay_tr_timer.counter_3_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25068\,
            in1 => \N__25417\,
            in2 => \_gnd_net_\,
            in3 => \N__24725\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            clk => \N__50314\,
            ce => \N__25160\,
            sr => \N__49468\
        );

    \delay_measurement_inst.delay_tr_timer.counter_4_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25077\,
            in1 => \N__25393\,
            in2 => \_gnd_net_\,
            in3 => \N__24722\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            clk => \N__50314\,
            ce => \N__25160\,
            sr => \N__49468\
        );

    \delay_measurement_inst.delay_tr_timer.counter_5_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25069\,
            in1 => \N__25369\,
            in2 => \_gnd_net_\,
            in3 => \N__24881\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            clk => \N__50314\,
            ce => \N__25160\,
            sr => \N__49468\
        );

    \delay_measurement_inst.delay_tr_timer.counter_6_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25078\,
            in1 => \N__25345\,
            in2 => \_gnd_net_\,
            in3 => \N__24878\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            clk => \N__50314\,
            ce => \N__25160\,
            sr => \N__49468\
        );

    \delay_measurement_inst.delay_tr_timer.counter_7_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25070\,
            in1 => \N__25321\,
            in2 => \_gnd_net_\,
            in3 => \N__24875\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            clk => \N__50314\,
            ce => \N__25160\,
            sr => \N__49468\
        );

    \delay_measurement_inst.delay_tr_timer.counter_8_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25066\,
            in1 => \N__25297\,
            in2 => \_gnd_net_\,
            in3 => \N__24872\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_7_8_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            clk => \N__50306\,
            ce => \N__25149\,
            sr => \N__49475\
        );

    \delay_measurement_inst.delay_tr_timer.counter_9_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25102\,
            in1 => \N__25678\,
            in2 => \_gnd_net_\,
            in3 => \N__24869\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            clk => \N__50306\,
            ce => \N__25149\,
            sr => \N__49475\
        );

    \delay_measurement_inst.delay_tr_timer.counter_10_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25063\,
            in1 => \N__25654\,
            in2 => \_gnd_net_\,
            in3 => \N__24866\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            clk => \N__50306\,
            ce => \N__25149\,
            sr => \N__49475\
        );

    \delay_measurement_inst.delay_tr_timer.counter_11_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25099\,
            in1 => \N__25630\,
            in2 => \_gnd_net_\,
            in3 => \N__24863\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            clk => \N__50306\,
            ce => \N__25149\,
            sr => \N__49475\
        );

    \delay_measurement_inst.delay_tr_timer.counter_12_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25064\,
            in1 => \N__25606\,
            in2 => \_gnd_net_\,
            in3 => \N__24860\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            clk => \N__50306\,
            ce => \N__25149\,
            sr => \N__49475\
        );

    \delay_measurement_inst.delay_tr_timer.counter_13_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25100\,
            in1 => \N__25582\,
            in2 => \_gnd_net_\,
            in3 => \N__24857\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            clk => \N__50306\,
            ce => \N__25149\,
            sr => \N__49475\
        );

    \delay_measurement_inst.delay_tr_timer.counter_14_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25065\,
            in1 => \N__25558\,
            in2 => \_gnd_net_\,
            in3 => \N__24908\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            clk => \N__50306\,
            ce => \N__25149\,
            sr => \N__49475\
        );

    \delay_measurement_inst.delay_tr_timer.counter_15_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25101\,
            in1 => \N__25534\,
            in2 => \_gnd_net_\,
            in3 => \N__24905\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            clk => \N__50306\,
            ce => \N__25149\,
            sr => \N__49475\
        );

    \delay_measurement_inst.delay_tr_timer.counter_16_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25079\,
            in1 => \N__25510\,
            in2 => \_gnd_net_\,
            in3 => \N__24902\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_7_9_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            clk => \N__50297\,
            ce => \N__25156\,
            sr => \N__49482\
        );

    \delay_measurement_inst.delay_tr_timer.counter_17_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25095\,
            in1 => \N__25891\,
            in2 => \_gnd_net_\,
            in3 => \N__24899\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            clk => \N__50297\,
            ce => \N__25156\,
            sr => \N__49482\
        );

    \delay_measurement_inst.delay_tr_timer.counter_18_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25080\,
            in1 => \N__25867\,
            in2 => \_gnd_net_\,
            in3 => \N__24896\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            clk => \N__50297\,
            ce => \N__25156\,
            sr => \N__49482\
        );

    \delay_measurement_inst.delay_tr_timer.counter_19_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25096\,
            in1 => \N__25843\,
            in2 => \_gnd_net_\,
            in3 => \N__24893\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            clk => \N__50297\,
            ce => \N__25156\,
            sr => \N__49482\
        );

    \delay_measurement_inst.delay_tr_timer.counter_20_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25081\,
            in1 => \N__25819\,
            in2 => \_gnd_net_\,
            in3 => \N__24890\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            clk => \N__50297\,
            ce => \N__25156\,
            sr => \N__49482\
        );

    \delay_measurement_inst.delay_tr_timer.counter_21_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25097\,
            in1 => \N__25795\,
            in2 => \_gnd_net_\,
            in3 => \N__24887\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            clk => \N__50297\,
            ce => \N__25156\,
            sr => \N__49482\
        );

    \delay_measurement_inst.delay_tr_timer.counter_22_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25082\,
            in1 => \N__25771\,
            in2 => \_gnd_net_\,
            in3 => \N__24884\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            clk => \N__50297\,
            ce => \N__25156\,
            sr => \N__49482\
        );

    \delay_measurement_inst.delay_tr_timer.counter_23_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25098\,
            in1 => \N__25747\,
            in2 => \_gnd_net_\,
            in3 => \N__24929\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            clk => \N__50297\,
            ce => \N__25156\,
            sr => \N__49482\
        );

    \delay_measurement_inst.delay_tr_timer.counter_24_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25071\,
            in1 => \N__25723\,
            in2 => \_gnd_net_\,
            in3 => \N__24926\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_7_10_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            clk => \N__50284\,
            ce => \N__25148\,
            sr => \N__49488\
        );

    \delay_measurement_inst.delay_tr_timer.counter_25_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25108\,
            in1 => \N__25699\,
            in2 => \_gnd_net_\,
            in3 => \N__24923\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            clk => \N__50284\,
            ce => \N__25148\,
            sr => \N__49488\
        );

    \delay_measurement_inst.delay_tr_timer.counter_26_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25072\,
            in1 => \N__25984\,
            in2 => \_gnd_net_\,
            in3 => \N__24920\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            clk => \N__50284\,
            ce => \N__25148\,
            sr => \N__49488\
        );

    \delay_measurement_inst.delay_tr_timer.counter_27_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25109\,
            in1 => \N__25948\,
            in2 => \_gnd_net_\,
            in3 => \N__24917\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            clk => \N__50284\,
            ce => \N__25148\,
            sr => \N__49488\
        );

    \delay_measurement_inst.delay_tr_timer.counter_28_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25073\,
            in1 => \N__26000\,
            in2 => \_gnd_net_\,
            in3 => \N__24914\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_28\,
            clk => \N__50284\,
            ce => \N__25148\,
            sr => \N__49488\
        );

    \delay_measurement_inst.delay_tr_timer.counter_29_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__25964\,
            in1 => \N__25074\,
            in2 => \_gnd_net_\,
            in3 => \N__24911\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50284\,
            ce => \N__25148\,
            sr => \N__49488\
        );

    \phase_controller_inst2.state_RNIG7JF_2_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24950\,
            in2 => \_gnd_net_\,
            in3 => \N__24976\,
            lcout => \phase_controller_inst2.state_RNIG7JFZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__31255\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31294\,
            lcout => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31389\,
            in2 => \_gnd_net_\,
            in3 => \N__31350\,
            lcout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33870\,
            in1 => \N__33900\,
            in2 => \_gnd_net_\,
            in3 => \N__34742\,
            lcout => \elapsed_time_ns_1_RNI3EPBB_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1_30_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__31390\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31351\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1Z0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_tr_RNO_0_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__24945\,
            in1 => \N__26218\,
            in2 => \N__24977\,
            in3 => \N__25275\,
            lcout => \phase_controller_inst2.start_timer_tr_RNO_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26408\,
            lcout => \delay_measurement_inst.delay_tr_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI54EN_30_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31595\,
            in2 => \_gnd_net_\,
            in3 => \N__27413\,
            lcout => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.time_passed_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010001011100010"
        )
    port map (
            in0 => \N__24974\,
            in1 => \N__35074\,
            in2 => \N__31259\,
            in3 => \N__37661\,
            lcout => \phase_controller_inst2.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50248\,
            ce => 'H',
            sr => \N__49500\
        );

    \phase_controller_inst2.start_timer_tr_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__46926\,
            in1 => \N__24983\,
            in2 => \N__31573\,
            in3 => \N__25121\,
            lcout => \phase_controller_inst2.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50248\,
            ce => 'H',
            sr => \N__49500\
        );

    \phase_controller_inst2.state_2_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__25185\,
            in1 => \N__24949\,
            in2 => \N__26268\,
            in3 => \N__24975\,
            lcout => \phase_controller_inst2.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50248\,
            ce => 'H',
            sr => \N__49500\
        );

    \phase_controller_inst2.stoper_tr.start_latched_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31565\,
            lcout => \phase_controller_inst2.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50248\,
            ce => 'H',
            sr => \N__49500\
        );

    \phase_controller_inst2.state_3_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111011100"
        )
    port map (
            in0 => \N__25186\,
            in1 => \N__25120\,
            in2 => \N__26269\,
            in3 => \N__33581\,
            lcout => \phase_controller_inst2.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50248\,
            ce => 'H',
            sr => \N__49500\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__26137\,
            in1 => \N__26157\,
            in2 => \N__25241\,
            in3 => \N__29162\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__29161\,
            in1 => \N__26136\,
            in2 => \N__26159\,
            in3 => \N__25237\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_27_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31178\,
            in1 => \N__31199\,
            in2 => \_gnd_net_\,
            in3 => \N__34815\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50237\,
            ce => \N__29768\,
            sr => \N__49504\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__25207\,
            in1 => \N__26100\,
            in2 => \N__25229\,
            in3 => \N__26118\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001100"
        )
    port map (
            in0 => \N__26119\,
            in1 => \N__25228\,
            in2 => \N__26102\,
            in3 => \N__25208\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_hc_RNO_0_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25193\,
            in2 => \_gnd_net_\,
            in3 => \N__26264\,
            lcout => \phase_controller_inst2.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26406\,
            in2 => \N__26306\,
            in3 => \N__26330\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_201_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__31604\,
            in1 => \N__26446\,
            in2 => \_gnd_net_\,
            in3 => \N__31569\,
            lcout => \phase_controller_inst2.stoper_tr.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_RNI9M3O_0_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26073\,
            in2 => \_gnd_net_\,
            in3 => \N__25252\,
            lcout => \phase_controller_inst2.state_RNI9M3OZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_1_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__26207\,
            in1 => \N__25277\,
            in2 => \_gnd_net_\,
            in3 => \N__26425\,
            lcout => \phase_controller_inst2.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50215\,
            ce => 'H',
            sr => \N__49512\
        );

    \phase_controller_inst2.state_0_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__26075\,
            in1 => \N__25276\,
            in2 => \N__26217\,
            in3 => \N__25253\,
            lcout => \phase_controller_inst2.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50215\,
            ce => 'H',
            sr => \N__49512\
        );

    \delay_measurement_inst.delay_tr_timer.running_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__26407\,
            in1 => \N__26302\,
            in2 => \_gnd_net_\,
            in3 => \N__26327\,
            lcout => \delay_measurement_inst.delay_tr_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50215\,
            ce => 'H',
            sr => \N__49512\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28966\,
            in1 => \N__28938\,
            in2 => \_gnd_net_\,
            in3 => \N__34709\,
            lcout => \elapsed_time_ns_1_RNI1CPBB_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29189\,
            in1 => \N__34019\,
            in2 => \N__30807\,
            in3 => \N__32168\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25489\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50315\,
            ce => \N__26381\,
            sr => \N__49454\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25468\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50315\,
            ce => \N__26381\,
            sr => \N__49454\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29190\,
            in1 => \N__29217\,
            in2 => \_gnd_net_\,
            in3 => \N__34581\,
            lcout => \elapsed_time_ns_1_RNIFE91B_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30800\,
            in2 => \N__34711\,
            in3 => \N__30831\,
            lcout => \elapsed_time_ns_1_RNIGF91B_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25440\,
            in2 => \N__25490\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\,
            ltout => OPEN,
            carryin => \bfn_8_7_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__50307\,
            ce => \N__26380\,
            sr => \N__49461\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25416\,
            in2 => \N__25469\,
            in3 => \N__25448\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__50307\,
            ce => \N__26380\,
            sr => \N__49461\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25392\,
            in2 => \N__25445\,
            in3 => \N__25424\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__50307\,
            ce => \N__26380\,
            sr => \N__49461\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25368\,
            in2 => \N__25421\,
            in3 => \N__25400\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__50307\,
            ce => \N__26380\,
            sr => \N__49461\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25344\,
            in2 => \N__25397\,
            in3 => \N__25376\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__50307\,
            ce => \N__26380\,
            sr => \N__49461\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25320\,
            in2 => \N__25373\,
            in3 => \N__25352\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__50307\,
            ce => \N__26380\,
            sr => \N__49461\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25296\,
            in2 => \N__25349\,
            in3 => \N__25328\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__50307\,
            ce => \N__26380\,
            sr => \N__49461\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25677\,
            in2 => \N__25325\,
            in3 => \N__25304\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__50307\,
            ce => \N__26380\,
            sr => \N__49461\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25653\,
            in2 => \N__25301\,
            in3 => \N__25280\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__50298\,
            ce => \N__26371\,
            sr => \N__49469\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25629\,
            in2 => \N__25682\,
            in3 => \N__25661\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__50298\,
            ce => \N__26371\,
            sr => \N__49469\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25605\,
            in2 => \N__25658\,
            in3 => \N__25637\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__50298\,
            ce => \N__26371\,
            sr => \N__49469\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25581\,
            in2 => \N__25634\,
            in3 => \N__25613\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__50298\,
            ce => \N__26371\,
            sr => \N__49469\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25557\,
            in2 => \N__25610\,
            in3 => \N__25589\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__50298\,
            ce => \N__26371\,
            sr => \N__49469\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25533\,
            in2 => \N__25586\,
            in3 => \N__25565\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__50298\,
            ce => \N__26371\,
            sr => \N__49469\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25509\,
            in2 => \N__25562\,
            in3 => \N__25541\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__50298\,
            ce => \N__26371\,
            sr => \N__49469\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25890\,
            in2 => \N__25538\,
            in3 => \N__25517\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__50298\,
            ce => \N__26371\,
            sr => \N__49469\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25866\,
            in2 => \N__25514\,
            in3 => \N__25493\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\,
            ltout => OPEN,
            carryin => \bfn_8_9_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__50285\,
            ce => \N__26379\,
            sr => \N__49476\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25842\,
            in2 => \N__25895\,
            in3 => \N__25874\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__50285\,
            ce => \N__26379\,
            sr => \N__49476\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25818\,
            in2 => \N__25871\,
            in3 => \N__25850\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__50285\,
            ce => \N__26379\,
            sr => \N__49476\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25794\,
            in2 => \N__25847\,
            in3 => \N__25826\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__50285\,
            ce => \N__26379\,
            sr => \N__49476\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25770\,
            in2 => \N__25823\,
            in3 => \N__25802\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__50285\,
            ce => \N__26379\,
            sr => \N__49476\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25746\,
            in2 => \N__25799\,
            in3 => \N__25778\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__50285\,
            ce => \N__26379\,
            sr => \N__49476\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25722\,
            in2 => \N__25775\,
            in3 => \N__25754\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__50285\,
            ce => \N__26379\,
            sr => \N__49476\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25698\,
            in2 => \N__25751\,
            in3 => \N__25730\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__50285\,
            ce => \N__26379\,
            sr => \N__49476\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25983\,
            in2 => \N__25727\,
            in3 => \N__25706\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\,
            ltout => OPEN,
            carryin => \bfn_8_10_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__50272\,
            ce => \N__26372\,
            sr => \N__49483\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25947\,
            in2 => \N__25703\,
            in3 => \N__26003\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__50272\,
            ce => \N__26372\,
            sr => \N__49483\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25999\,
            in2 => \N__25988\,
            in3 => \N__25967\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__50272\,
            ce => \N__26372\,
            sr => \N__49483\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25963\,
            in2 => \N__25952\,
            in3 => \N__25931\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__50272\,
            ce => \N__26372\,
            sr => \N__49483\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25928\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50272\,
            ce => \N__26372\,
            sr => \N__49483\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31331\,
            in2 => \N__25925\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_11_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31523\,
            in1 => \N__26852\,
            in2 => \_gnd_net_\,
            in3 => \N__25916\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \N__50261\,
            ce => 'H',
            sr => \N__49489\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__31527\,
            in1 => \N__26831\,
            in2 => \N__25913\,
            in3 => \N__25904\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \N__50261\,
            ce => 'H',
            sr => \N__49489\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31524\,
            in1 => \N__26810\,
            in2 => \_gnd_net_\,
            in3 => \N__25901\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \N__50261\,
            ce => 'H',
            sr => \N__49489\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31528\,
            in1 => \N__26777\,
            in2 => \_gnd_net_\,
            in3 => \N__25898\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \N__50261\,
            ce => 'H',
            sr => \N__49489\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31525\,
            in1 => \N__26756\,
            in2 => \_gnd_net_\,
            in3 => \N__26030\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \N__50261\,
            ce => 'H',
            sr => \N__49489\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31529\,
            in1 => \N__27128\,
            in2 => \_gnd_net_\,
            in3 => \N__26027\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \N__50261\,
            ce => 'H',
            sr => \N__49489\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31526\,
            in1 => \N__27107\,
            in2 => \_gnd_net_\,
            in3 => \N__26024\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \N__50261\,
            ce => 'H',
            sr => \N__49489\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31515\,
            in1 => \N__27089\,
            in2 => \_gnd_net_\,
            in3 => \N__26021\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_8_12_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \N__50249\,
            ce => 'H',
            sr => \N__49493\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31508\,
            in1 => \N__27058\,
            in2 => \_gnd_net_\,
            in3 => \N__26018\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \N__50249\,
            ce => 'H',
            sr => \N__49493\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31512\,
            in1 => \N__27026\,
            in2 => \_gnd_net_\,
            in3 => \N__26015\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \N__50249\,
            ce => 'H',
            sr => \N__49493\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31509\,
            in1 => \N__26993\,
            in2 => \_gnd_net_\,
            in3 => \N__26012\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \N__50249\,
            ce => 'H',
            sr => \N__49493\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31513\,
            in1 => \N__26975\,
            in2 => \_gnd_net_\,
            in3 => \N__26009\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \N__50249\,
            ce => 'H',
            sr => \N__49493\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31510\,
            in1 => \N__26942\,
            in2 => \_gnd_net_\,
            in3 => \N__26006\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \N__50249\,
            ce => 'H',
            sr => \N__49493\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31514\,
            in1 => \N__27248\,
            in2 => \_gnd_net_\,
            in3 => \N__26057\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \N__50249\,
            ce => 'H',
            sr => \N__49493\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31511\,
            in1 => \N__29863\,
            in2 => \_gnd_net_\,
            in3 => \N__26054\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \N__50249\,
            ce => 'H',
            sr => \N__49493\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31519\,
            in1 => \N__29887\,
            in2 => \_gnd_net_\,
            in3 => \N__26051\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_8_13_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \N__50238\,
            ce => 'H',
            sr => \N__49497\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31537\,
            in1 => \N__29362\,
            in2 => \_gnd_net_\,
            in3 => \N__26048\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \N__50238\,
            ce => 'H',
            sr => \N__49497\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31520\,
            in1 => \N__29338\,
            in2 => \_gnd_net_\,
            in3 => \N__26045\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \N__50238\,
            ce => 'H',
            sr => \N__49497\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31538\,
            in1 => \N__29517\,
            in2 => \_gnd_net_\,
            in3 => \N__26042\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \N__50238\,
            ce => 'H',
            sr => \N__49497\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31521\,
            in1 => \N__29496\,
            in2 => \_gnd_net_\,
            in3 => \N__26039\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\,
            clk => \N__50238\,
            ce => 'H',
            sr => \N__49497\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31539\,
            in1 => \N__26485\,
            in2 => \_gnd_net_\,
            in3 => \N__26036\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\,
            clk => \N__50238\,
            ce => 'H',
            sr => \N__49497\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31522\,
            in1 => \N__26506\,
            in2 => \_gnd_net_\,
            in3 => \N__26033\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\,
            clk => \N__50238\,
            ce => 'H',
            sr => \N__49497\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31540\,
            in1 => \N__26628\,
            in2 => \_gnd_net_\,
            in3 => \N__26165\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\,
            clk => \N__50238\,
            ce => 'H',
            sr => \N__49497\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31530\,
            in1 => \N__26649\,
            in2 => \_gnd_net_\,
            in3 => \N__26162\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_8_14_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\,
            clk => \N__50226\,
            ce => 'H',
            sr => \N__49501\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31534\,
            in1 => \N__26158\,
            in2 => \_gnd_net_\,
            in3 => \N__26141\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\,
            clk => \N__50226\,
            ce => 'H',
            sr => \N__49501\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31531\,
            in1 => \N__26138\,
            in2 => \_gnd_net_\,
            in3 => \N__26123\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\,
            clk => \N__50226\,
            ce => 'H',
            sr => \N__49501\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31535\,
            in1 => \N__26120\,
            in2 => \_gnd_net_\,
            in3 => \N__26105\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\,
            clk => \N__50226\,
            ce => 'H',
            sr => \N__49501\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31532\,
            in1 => \N__26101\,
            in2 => \_gnd_net_\,
            in3 => \N__26084\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\,
            clk => \N__50226\,
            ce => 'H',
            sr => \N__49501\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31536\,
            in1 => \N__26922\,
            in2 => \_gnd_net_\,
            in3 => \N__26081\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\,
            clk => \N__50226\,
            ce => 'H',
            sr => \N__49501\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31533\,
            in1 => \N__26884\,
            in2 => \_gnd_net_\,
            in3 => \N__26078\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50226\,
            ce => 'H',
            sr => \N__49501\
        );

    \phase_controller_inst2.stoper_tr.time_passed_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010001011100010"
        )
    port map (
            in0 => \N__26074\,
            in1 => \N__31380\,
            in2 => \N__31615\,
            in3 => \N__27408\,
            lcout => \phase_controller_inst2.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50216\,
            ce => 'H',
            sr => \N__49505\
        );

    \phase_controller_inst2.stoper_tr.running_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000101110"
        )
    port map (
            in0 => \N__26447\,
            in1 => \N__31379\,
            in2 => \N__31616\,
            in3 => \N__27409\,
            lcout => \phase_controller_inst2.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50216\,
            ce => 'H',
            sr => \N__49505\
        );

    \phase_controller_inst2.start_timer_hc_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101110101010"
        )
    port map (
            in0 => \N__26435\,
            in1 => \N__26429\,
            in2 => \N__46931\,
            in3 => \N__31280\,
            lcout => \phase_controller_inst2.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50216\,
            ce => 'H',
            sr => \N__49505\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26405\,
            in2 => \_gnd_net_\,
            in3 => \N__26298\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_200_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.start_timer_tr_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26328\,
            lcout => \delay_measurement_inst.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26282\,
            ce => 'H',
            sr => \N__49513\
        );

    \delay_measurement_inst.stop_timer_tr_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26329\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.stop_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26282\,
            ce => 'H',
            sr => \N__49513\
        );

    \phase_controller_inst2.S1_LC_8_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26273\,
            lcout => s3_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50170\,
            ce => 'H',
            sr => \N__49550\
        );

    \phase_controller_inst2.S2_LC_8_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26225\,
            lcout => s4_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50170\,
            ce => 'H',
            sr => \N__49550\
        );

    \GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_8_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50324\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_clock_output_0_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_23_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34710\,
            in1 => \N__28962\,
            in2 => \_gnd_net_\,
            in3 => \N__28946\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50316\,
            ce => \N__29758\,
            sr => \N__49437\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001100"
        )
    port map (
            in0 => \N__26492\,
            in1 => \N__26528\,
            in2 => \N__26519\,
            in3 => \N__26470\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001010111011"
        )
    port map (
            in0 => \N__26527\,
            in1 => \N__26518\,
            in2 => \N__26471\,
            in3 => \N__26491\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_22_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34613\,
            in1 => \N__28618\,
            in2 => \_gnd_net_\,
            in3 => \N__28639\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50308\,
            ce => \N__29759\,
            sr => \N__49447\
        );

    \phase_controller_inst2.stoper_tr.target_time_12_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28699\,
            in1 => \N__28681\,
            in2 => \_gnd_net_\,
            in3 => \N__34614\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50308\,
            ce => \N__29759\,
            sr => \N__49447\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__29105\,
            in1 => \N__31164\,
            in2 => \_gnd_net_\,
            in3 => \N__26459\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__32253\,
            in1 => \N__26555\,
            in2 => \N__26453\,
            in3 => \N__26564\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3\,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__29025\,
            in1 => \_gnd_net_\,
            in2 => \N__26450\,
            in3 => \N__29005\,
            lcout => \elapsed_time_ns_1_RNIVAQBB_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34364\,
            in2 => \_gnd_net_\,
            in3 => \N__34871\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28721\,
            in1 => \N__28740\,
            in2 => \_gnd_net_\,
            in3 => \N__34612\,
            lcout => \elapsed_time_ns_1_RNIHG91B_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28818\,
            in1 => \N__28770\,
            in2 => \N__28679\,
            in3 => \N__29578\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__29441\,
            in1 => \N__28739\,
            in2 => \N__26573\,
            in3 => \N__26570\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28877\,
            in1 => \N__31104\,
            in2 => \N__29006\,
            in3 => \N__33860\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26537\,
            in1 => \N__26549\,
            in2 => \N__26558\,
            in3 => \N__26543\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29270\,
            in1 => \N__26690\,
            in2 => \N__33399\,
            in3 => \N__29631\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__33022\,
            in1 => \N__29803\,
            in2 => \N__33267\,
            in3 => \N__26722\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28928\,
            in1 => \N__29678\,
            in2 => \N__28607\,
            in3 => \N__34938\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29679\,
            in1 => \N__29656\,
            in2 => \_gnd_net_\,
            in3 => \N__34604\,
            lcout => \elapsed_time_ns_1_RNIV9PBB_0_21\,
            ltout => \elapsed_time_ns_1_RNIV9PBB_0_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_21_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__34605\,
            in1 => \_gnd_net_\,
            in2 => \N__26531\,
            in3 => \N__29680\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50286\,
            ce => \N__34321\,
            sr => \N__49462\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__26597\,
            in1 => \N__32966\,
            in2 => \N__32993\,
            in3 => \N__26585\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__26691\,
            in1 => \N__26671\,
            in2 => \N__34765\,
            in3 => \_gnd_net_\,
            lcout => \elapsed_time_ns_1_RNI5FOBB_0_18\,
            ltout => \elapsed_time_ns_1_RNI5FOBB_0_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_18_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34684\,
            in2 => \N__26600\,
            in3 => \N__26692\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50273\,
            ce => \N__34276\,
            sr => \N__49470\
        );

    \phase_controller_inst1.stoper_tr.target_time_19_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__34685\,
            in1 => \N__29308\,
            in2 => \N__29286\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50273\,
            ce => \N__34276\,
            sr => \N__49470\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__26596\,
            in1 => \N__32965\,
            in2 => \N__32992\,
            in3 => \N__26584\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34679\,
            in1 => \N__26734\,
            in2 => \_gnd_net_\,
            in3 => \N__26717\,
            lcout => \elapsed_time_ns_1_RNI1BOBB_0_14\,
            ltout => \elapsed_time_ns_1_RNI1BOBB_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_14_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__26718\,
            in1 => \_gnd_net_\,
            in2 => \N__26576\,
            in3 => \N__34683\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50273\,
            ce => \N__34276\,
            sr => \N__49470\
        );

    \phase_controller_inst2.stoper_tr.target_time_24_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34948\,
            in1 => \N__33830\,
            in2 => \_gnd_net_\,
            in3 => \N__34772\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50262\,
            ce => \N__29762\,
            sr => \N__49477\
        );

    \phase_controller_inst2.stoper_tr.target_time_30_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__29026\,
            in1 => \N__34767\,
            in2 => \_gnd_net_\,
            in3 => \N__28994\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50262\,
            ce => \N__29762\,
            sr => \N__49477\
        );

    \phase_controller_inst2.stoper_tr.target_time_10_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28799\,
            in1 => \N__28782\,
            in2 => \_gnd_net_\,
            in3 => \N__34770\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50262\,
            ce => \N__29762\,
            sr => \N__49477\
        );

    \phase_controller_inst2.stoper_tr.target_time_5_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34769\,
            in1 => \N__28748\,
            in2 => \_gnd_net_\,
            in3 => \N__28720\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50262\,
            ce => \N__29762\,
            sr => \N__49477\
        );

    \phase_controller_inst2.stoper_tr.target_time_14_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26735\,
            in1 => \N__26723\,
            in2 => \_gnd_net_\,
            in3 => \N__34771\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50262\,
            ce => \N__29762\,
            sr => \N__49477\
        );

    \phase_controller_inst2.stoper_tr.target_time_11_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28829\,
            in1 => \N__34766\,
            in2 => \_gnd_net_\,
            in3 => \N__28844\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50262\,
            ce => \N__29762\,
            sr => \N__49477\
        );

    \phase_controller_inst2.stoper_tr.target_time_7_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34913\,
            in1 => \N__34885\,
            in2 => \_gnd_net_\,
            in3 => \N__34773\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50262\,
            ce => \N__29762\,
            sr => \N__49477\
        );

    \phase_controller_inst2.stoper_tr.target_time_18_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34768\,
            in1 => \N__26696\,
            in2 => \_gnd_net_\,
            in3 => \N__26672\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50262\,
            ce => \N__29762\,
            sr => \N__49477\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__26651\,
            in1 => \N__26629\,
            in2 => \N__26612\,
            in3 => \N__26660\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__26659\,
            in1 => \N__26650\,
            in2 => \N__26633\,
            in3 => \N__26608\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_25_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__33901\,
            in1 => \N__33874\,
            in2 => \_gnd_net_\,
            in3 => \N__34775\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50250\,
            ce => \N__29764\,
            sr => \N__49484\
        );

    \phase_controller_inst2.stoper_tr.target_time_31_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34774\,
            in1 => \N__32243\,
            in2 => \_gnd_net_\,
            in3 => \N__32219\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50250\,
            ce => \N__29764\,
            sr => \N__49484\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010011011101"
        )
    port map (
            in0 => \N__26869\,
            in1 => \N__26893\,
            in2 => \N__26906\,
            in3 => \N__26923\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_30_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__26924\,
            in1 => \N__26905\,
            in2 => \N__26894\,
            in3 => \N__26870\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29543\,
            in2 => \N__26861\,
            in3 => \N__31327\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_9_12_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29237\,
            in2 => \N__26840\,
            in3 => \N__26851\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29174\,
            in2 => \N__26819\,
            in3 => \N__26830\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29168\,
            in2 => \N__26798\,
            in3 => \N__26809\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26765\,
            in2 => \N__26789\,
            in3 => \N__26776\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29399\,
            in2 => \N__26744\,
            in3 => \N__26755\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27137\,
            in2 => \N__27116\,
            in3 => \N__27127\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27095\,
            in2 => \N__29147\,
            in3 => \N__27106\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_7\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27077\,
            in2 => \N__29552\,
            in3 => \N__27088\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_9_13_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27071\,
            in2 => \N__27044\,
            in3 => \N__27062\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27035\,
            in2 => \N__27014\,
            in3 => \N__27025\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26981\,
            in2 => \N__27005\,
            in3 => \N__26992\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26974\,
            in1 => \N__29693\,
            in2 => \N__26963\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26930\,
            in2 => \N__26954\,
            in3 => \N__26941\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27236\,
            in2 => \N__29777\,
            in3 => \N__27247\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29849\,
            in2 => \N__29906\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_15\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29324\,
            in2 => \N__29393\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_14_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29468\,
            in2 => \N__29537\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27230\,
            in2 => \N__27221\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_20\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27209\,
            in2 => \N__27200\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_22\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27185\,
            in2 => \N__27176\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_24\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27164\,
            in2 => \N__27152\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_26\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_30_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27440\,
            in2 => \N__27431\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_28\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27416\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31748\,
            in1 => \N__27392\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axb_0\,
            ltout => OPEN,
            carryin => \bfn_9_15_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_1_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31739\,
            in2 => \_gnd_net_\,
            in3 => \N__27362\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            clk => \N__50205\,
            ce => 'H',
            sr => \N__49502\
        );

    \current_shift_inst.PI_CTRL.error_control_2_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31727\,
            in2 => \_gnd_net_\,
            in3 => \N__27332\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            clk => \N__50205\,
            ce => 'H',
            sr => \N__49502\
        );

    \current_shift_inst.PI_CTRL.error_control_3_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31715\,
            in2 => \_gnd_net_\,
            in3 => \N__27302\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            clk => \N__50205\,
            ce => 'H',
            sr => \N__49502\
        );

    \current_shift_inst.PI_CTRL.error_control_4_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31703\,
            in2 => \_gnd_net_\,
            in3 => \N__27278\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            clk => \N__50205\,
            ce => 'H',
            sr => \N__49502\
        );

    \current_shift_inst.PI_CTRL.error_control_5_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31691\,
            in3 => \N__27251\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            clk => \N__50205\,
            ce => 'H',
            sr => \N__49502\
        );

    \current_shift_inst.PI_CTRL.error_control_6_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31676\,
            in3 => \N__27683\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            clk => \N__50205\,
            ce => 'H',
            sr => \N__49502\
        );

    \current_shift_inst.PI_CTRL.error_control_7_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31661\,
            in3 => \N__27653\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            clk => \N__50205\,
            ce => 'H',
            sr => \N__49502\
        );

    \current_shift_inst.PI_CTRL.error_control_8_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31928\,
            in2 => \_gnd_net_\,
            in3 => \N__27629\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_8\,
            ltout => OPEN,
            carryin => \bfn_9_16_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            clk => \N__50196\,
            ce => 'H',
            sr => \N__49506\
        );

    \current_shift_inst.PI_CTRL.error_control_9_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31910\,
            in2 => \_gnd_net_\,
            in3 => \N__27596\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            clk => \N__50196\,
            ce => 'H',
            sr => \N__49506\
        );

    \current_shift_inst.PI_CTRL.error_control_10_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31889\,
            in2 => \_gnd_net_\,
            in3 => \N__27560\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            clk => \N__50196\,
            ce => 'H',
            sr => \N__49506\
        );

    \current_shift_inst.PI_CTRL.error_control_11_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31874\,
            in2 => \_gnd_net_\,
            in3 => \N__27530\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            clk => \N__50196\,
            ce => 'H',
            sr => \N__49506\
        );

    \current_shift_inst.PI_CTRL.error_control_12_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31862\,
            in3 => \N__27500\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            clk => \N__50196\,
            ce => 'H',
            sr => \N__49506\
        );

    \current_shift_inst.PI_CTRL.error_control_13_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31847\,
            in3 => \N__27473\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_13\,
            clk => \N__50196\,
            ce => 'H',
            sr => \N__49506\
        );

    \current_shift_inst.PI_CTRL.error_control_14_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31832\,
            in3 => \N__27443\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_14\,
            clk => \N__50196\,
            ce => 'H',
            sr => \N__49506\
        );

    \current_shift_inst.PI_CTRL.error_control_15_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31817\,
            in3 => \N__27932\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_15\,
            clk => \N__50196\,
            ce => 'H',
            sr => \N__49506\
        );

    \current_shift_inst.PI_CTRL.error_control_16_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32048\,
            in3 => \N__27902\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_16\,
            ltout => OPEN,
            carryin => \bfn_9_17_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_16\,
            clk => \N__50190\,
            ce => 'H',
            sr => \N__49508\
        );

    \current_shift_inst.PI_CTRL.error_control_17_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32033\,
            in3 => \N__27866\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_17\,
            clk => \N__50190\,
            ce => 'H',
            sr => \N__49508\
        );

    \current_shift_inst.PI_CTRL.error_control_18_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32018\,
            in2 => \_gnd_net_\,
            in3 => \N__27836\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_18\,
            clk => \N__50190\,
            ce => 'H',
            sr => \N__49508\
        );

    \current_shift_inst.PI_CTRL.error_control_19_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31997\,
            in2 => \_gnd_net_\,
            in3 => \N__27803\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_19\,
            clk => \N__50190\,
            ce => 'H',
            sr => \N__49508\
        );

    \current_shift_inst.PI_CTRL.error_control_20_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31985\,
            in2 => \_gnd_net_\,
            in3 => \N__27767\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_20\,
            clk => \N__50190\,
            ce => 'H',
            sr => \N__49508\
        );

    \current_shift_inst.PI_CTRL.error_control_21_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31973\,
            in2 => \_gnd_net_\,
            in3 => \N__27740\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_21\,
            clk => \N__50190\,
            ce => 'H',
            sr => \N__49508\
        );

    \current_shift_inst.PI_CTRL.error_control_22_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31961\,
            in2 => \_gnd_net_\,
            in3 => \N__27707\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_22\,
            clk => \N__50190\,
            ce => 'H',
            sr => \N__49508\
        );

    \current_shift_inst.PI_CTRL.error_control_23_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31949\,
            in3 => \N__28178\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_23\,
            clk => \N__50190\,
            ce => 'H',
            sr => \N__49508\
        );

    \current_shift_inst.PI_CTRL.error_control_24_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32150\,
            in2 => \_gnd_net_\,
            in3 => \N__28145\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_24\,
            ltout => OPEN,
            carryin => \bfn_9_18_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_24\,
            clk => \N__50186\,
            ce => 'H',
            sr => \N__49514\
        );

    \current_shift_inst.PI_CTRL.error_control_25_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32138\,
            in3 => \N__28118\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_25\,
            clk => \N__50186\,
            ce => 'H',
            sr => \N__49514\
        );

    \current_shift_inst.PI_CTRL.error_control_26_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32123\,
            in2 => \_gnd_net_\,
            in3 => \N__28085\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_26\,
            clk => \N__50186\,
            ce => 'H',
            sr => \N__49514\
        );

    \current_shift_inst.PI_CTRL.error_control_27_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32111\,
            in2 => \_gnd_net_\,
            in3 => \N__28058\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_27\,
            clk => \N__50186\,
            ce => 'H',
            sr => \N__49514\
        );

    \current_shift_inst.PI_CTRL.error_control_28_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32099\,
            in3 => \N__28028\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_28\,
            clk => \N__50186\,
            ce => 'H',
            sr => \N__49514\
        );

    \current_shift_inst.PI_CTRL.error_control_29_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32084\,
            in2 => \_gnd_net_\,
            in3 => \N__28001\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_29\,
            clk => \N__50186\,
            ce => 'H',
            sr => \N__49514\
        );

    \current_shift_inst.PI_CTRL.error_control_30_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30107\,
            in2 => \_gnd_net_\,
            in3 => \N__27965\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_30\,
            clk => \N__50186\,
            ce => 'H',
            sr => \N__49514\
        );

    \current_shift_inst.PI_CTRL.error_control_31_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32069\,
            in2 => \_gnd_net_\,
            in3 => \N__28490\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50186\,
            ce => 'H',
            sr => \N__49514\
        );

    \current_shift_inst.PI_CTRL.prop_term_31_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28487\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50181\,
            ce => 'H',
            sr => \N__49521\
        );

    \current_shift_inst.PI_CTRL.control_out_10_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28466\,
            lcout => \N_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50174\,
            ce => 'H',
            sr => \N__49533\
        );

    \pwm_generator_inst.un3_threshold_cry_0_c_LC_9_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28403\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_26_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_9_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28379\,
            in2 => \_gnd_net_\,
            in3 => \N__28337\,
            lcout => \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_0\,
            carryout => \pwm_generator_inst.un3_threshold_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_9_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28334\,
            in2 => \_gnd_net_\,
            in3 => \N__28298\,
            lcout => \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_1\,
            carryout => \pwm_generator_inst.un3_threshold_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_9_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28295\,
            in2 => \_gnd_net_\,
            in3 => \N__28259\,
            lcout => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_2\,
            carryout => \pwm_generator_inst.un3_threshold_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_9_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30062\,
            in2 => \_gnd_net_\,
            in3 => \N__28235\,
            lcout => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_3\,
            carryout => \pwm_generator_inst.un3_threshold_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_9_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48431\,
            in2 => \N__30017\,
            in3 => \N__28211\,
            lcout => \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_4\,
            carryout => \pwm_generator_inst.un3_threshold_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_9_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29966\,
            in2 => \N__48440\,
            in3 => \N__28538\,
            lcout => \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_5\,
            carryout => \pwm_generator_inst.un3_threshold_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_9_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48435\,
            in2 => \N__29921\,
            in3 => \N__28511\,
            lcout => \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_6\,
            carryout => \pwm_generator_inst.un3_threshold_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_9_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30374\,
            in2 => \_gnd_net_\,
            in3 => \N__28493\,
            lcout => \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11\,
            ltout => OPEN,
            carryin => \bfn_9_27_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_9_c_LC_9_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30329\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_8\,
            carryout => \pwm_generator_inst.un3_threshold_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_10_c_LC_9_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30284\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_9\,
            carryout => \pwm_generator_inst.un3_threshold_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_11_c_LC_9_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30242\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_10\,
            carryout => \pwm_generator_inst.un3_threshold_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_12_c_LC_9_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30197\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_11\,
            carryout => \pwm_generator_inst.un3_threshold_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_13_c_LC_9_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30146\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_12\,
            carryout => \pwm_generator_inst.un3_threshold_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_14_c_LC_9_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30116\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_13\,
            carryout => \pwm_generator_inst.un3_threshold_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_15_c_LC_9_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30659\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_14\,
            carryout => \pwm_generator_inst.un3_threshold_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_16_c_LC_9_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30629\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_28_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_17_c_LC_9_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30599\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_16\,
            carryout => \pwm_generator_inst.un3_threshold_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_18_c_LC_9_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30569\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_17\,
            carryout => \pwm_generator_inst.un3_threshold_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_c_LC_9_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30548\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_18\,
            carryout => \pwm_generator_inst.un3_threshold_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_9_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28580\,
            lcout => \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D2_LC_10_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28565\,
            lcout => \il_min_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50309\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D1_LC_10_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28577\,
            lcout => \il_min_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50309\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28640\,
            in1 => \N__28617\,
            in2 => \_gnd_net_\,
            in3 => \N__34603\,
            lcout => \elapsed_time_ns_1_RNI0BPBB_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28906\,
            in1 => \N__28885\,
            in2 => \_gnd_net_\,
            in3 => \N__34601\,
            lcout => \elapsed_time_ns_1_RNI7IPBB_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34599\,
            in1 => \N__29307\,
            in2 => \_gnd_net_\,
            in3 => \N__29287\,
            lcout => \elapsed_time_ns_1_RNI6GOBB_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29419\,
            in1 => \N__29458\,
            in2 => \_gnd_net_\,
            in3 => \N__34600\,
            lcout => \elapsed_time_ns_1_RNIIH91B_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28700\,
            in1 => \N__28680\,
            in2 => \_gnd_net_\,
            in3 => \N__34602\,
            lcout => \elapsed_time_ns_1_RNIV8OBB_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29454\,
            in1 => \N__29415\,
            in2 => \_gnd_net_\,
            in3 => \N__34672\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50274\,
            ce => \N__34312\,
            sr => \N__49438\
        );

    \phase_controller_inst1.stoper_tr.target_time_5_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34669\,
            in1 => \N__28747\,
            in2 => \_gnd_net_\,
            in3 => \N__28719\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50274\,
            ce => \N__34312\,
            sr => \N__49438\
        );

    \phase_controller_inst1.stoper_tr.target_time_12_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28698\,
            in1 => \N__28682\,
            in2 => \_gnd_net_\,
            in3 => \N__34670\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50274\,
            ce => \N__34312\,
            sr => \N__49438\
        );

    \phase_controller_inst1.stoper_tr.target_time_22_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__34666\,
            in1 => \N__28638\,
            in2 => \N__28622\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50274\,
            ce => \N__34312\,
            sr => \N__49438\
        );

    \phase_controller_inst1.stoper_tr.target_time_3_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34668\,
            in1 => \N__29224\,
            in2 => \_gnd_net_\,
            in3 => \N__29197\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50274\,
            ce => \N__34312\,
            sr => \N__49438\
        );

    \phase_controller_inst1.stoper_tr.target_time_23_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28970\,
            in1 => \N__28945\,
            in2 => \_gnd_net_\,
            in3 => \N__34671\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50274\,
            ce => \N__34312\,
            sr => \N__49438\
        );

    \phase_controller_inst1.stoper_tr.target_time_29_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34667\,
            in1 => \N__28902\,
            in2 => \_gnd_net_\,
            in3 => \N__28884\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50274\,
            ce => \N__34312\,
            sr => \N__49438\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34608\,
            in1 => \N__28827\,
            in2 => \_gnd_net_\,
            in3 => \N__28840\,
            lcout => \elapsed_time_ns_1_RNIU7OBB_0_11\,
            ltout => \elapsed_time_ns_1_RNIU7OBB_0_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_11_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__28828\,
            in1 => \_gnd_net_\,
            in2 => \N__28802\,
            in3 => \N__34611\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50263\,
            ce => \N__34316\,
            sr => \N__49448\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34606\,
            in1 => \N__28783\,
            in2 => \_gnd_net_\,
            in3 => \N__28795\,
            lcout => \elapsed_time_ns_1_RNIT6OBB_0_10\,
            ltout => \elapsed_time_ns_1_RNIT6OBB_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_10_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__28784\,
            in1 => \_gnd_net_\,
            in2 => \N__28754\,
            in3 => \N__34610\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50263\,
            ce => \N__34316\,
            sr => \N__49448\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29592\,
            in1 => \N__29563\,
            in2 => \_gnd_net_\,
            in3 => \N__34607\,
            lcout => \elapsed_time_ns_1_RNILK91B_0_9\,
            ltout => \elapsed_time_ns_1_RNILK91B_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_9_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__34609\,
            in1 => \_gnd_net_\,
            in2 => \N__28751\,
            in3 => \N__29593\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50263\,
            ce => \N__34316\,
            sr => \N__49448\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011010100"
        )
    port map (
            in0 => \N__32920\,
            in1 => \N__29132\,
            in2 => \N__29123\,
            in3 => \N__32944\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29640\,
            in1 => \N__29611\,
            in2 => \_gnd_net_\,
            in3 => \N__34733\,
            lcout => \elapsed_time_ns_1_RNIU8PBB_0_20\,
            ltout => \elapsed_time_ns_1_RNIU8PBB_0_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_20_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__34735\,
            in1 => \_gnd_net_\,
            in2 => \N__29138\,
            in3 => \N__29641\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50252\,
            ce => \N__34263\,
            sr => \N__49455\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29817\,
            in1 => \N__29788\,
            in2 => \_gnd_net_\,
            in3 => \N__34732\,
            lcout => \elapsed_time_ns_1_RNI2COBB_0_15\,
            ltout => \elapsed_time_ns_1_RNI2COBB_0_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_15_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__34734\,
            in1 => \_gnd_net_\,
            in2 => \N__29135\,
            in3 => \N__29818\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50252\,
            ce => \N__34263\,
            sr => \N__49455\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__29131\,
            in1 => \N__32921\,
            in2 => \N__32945\,
            in3 => \N__29122\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__29054\,
            in1 => \N__33134\,
            in2 => \N__29045\,
            in3 => \N__33155\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_28_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29107\,
            in1 => \N__29075\,
            in2 => \_gnd_net_\,
            in3 => \N__34839\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50240\,
            ce => \N__34254\,
            sr => \N__49463\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__29053\,
            in1 => \N__33133\,
            in2 => \N__29044\,
            in3 => \N__33154\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_30_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29027\,
            in1 => \N__29001\,
            in2 => \_gnd_net_\,
            in3 => \N__34840\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50240\,
            ce => \N__34254\,
            sr => \N__49463\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011110010"
        )
    port map (
            in0 => \N__31646\,
            in1 => \N__33112\,
            in2 => \N__33083\,
            in3 => \N__31634\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__29368\,
            in1 => \N__29347\,
            in2 => \N__29249\,
            in3 => \N__29378\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__29377\,
            in1 => \N__29369\,
            in2 => \N__29348\,
            in3 => \N__29245\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_19_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29312\,
            in1 => \N__29288\,
            in2 => \_gnd_net_\,
            in3 => \N__34830\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50228\,
            ce => \N__29761\,
            sr => \N__49471\
        );

    \phase_controller_inst2.stoper_tr.target_time_2_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34828\,
            in1 => \N__34001\,
            in2 => \_gnd_net_\,
            in3 => \N__34043\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50228\,
            ce => \N__29761\,
            sr => \N__49471\
        );

    \phase_controller_inst2.stoper_tr.target_time_3_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29231\,
            in1 => \N__29201\,
            in2 => \_gnd_net_\,
            in3 => \N__34831\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50228\,
            ce => \N__29761\,
            sr => \N__49471\
        );

    \phase_controller_inst2.stoper_tr.target_time_4_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34829\,
            in1 => \N__30845\,
            in2 => \_gnd_net_\,
            in3 => \N__30814\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50228\,
            ce => \N__29761\,
            sr => \N__49471\
        );

    \phase_controller_inst2.stoper_tr.target_time_26_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34833\,
            in1 => \N__31121\,
            in2 => \_gnd_net_\,
            in3 => \N__31136\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50218\,
            ce => \N__29763\,
            sr => \N__49478\
        );

    \phase_controller_inst2.stoper_tr.target_time_8_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__34412\,
            in1 => \N__34838\,
            in2 => \_gnd_net_\,
            in3 => \N__34384\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50218\,
            ce => \N__29763\,
            sr => \N__49478\
        );

    \phase_controller_inst2.stoper_tr.target_time_13_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__33041\,
            in1 => \N__34835\,
            in2 => \_gnd_net_\,
            in3 => \N__33059\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50218\,
            ce => \N__29763\,
            sr => \N__49478\
        );

    \phase_controller_inst2.stoper_tr.target_time_21_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34832\,
            in1 => \N__29687\,
            in2 => \_gnd_net_\,
            in3 => \N__29663\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50218\,
            ce => \N__29763\,
            sr => \N__49478\
        );

    \phase_controller_inst2.stoper_tr.target_time_20_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29645\,
            in1 => \N__34837\,
            in2 => \_gnd_net_\,
            in3 => \N__29615\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50218\,
            ce => \N__29763\,
            sr => \N__49478\
        );

    \phase_controller_inst2.stoper_tr.target_time_9_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34834\,
            in1 => \N__29600\,
            in2 => \_gnd_net_\,
            in3 => \N__29567\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50218\,
            ce => \N__29763\,
            sr => \N__49478\
        );

    \phase_controller_inst2.stoper_tr.target_time_1_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__32744\,
            in1 => \N__34836\,
            in2 => \_gnd_net_\,
            in3 => \N__32186\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50218\,
            ce => \N__29763\,
            sr => \N__49478\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__29518\,
            in1 => \N__29528\,
            in2 => \N__29480\,
            in3 => \N__29500\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__29527\,
            in1 => \N__29519\,
            in2 => \N__29501\,
            in3 => \N__29479\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_6_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29462\,
            in1 => \N__29423\,
            in2 => \_gnd_net_\,
            in3 => \N__34844\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50207\,
            ce => \N__29765\,
            sr => \N__49485\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011110010"
        )
    port map (
            in0 => \N__29843\,
            in1 => \N__29869\,
            in2 => \N__29834\,
            in3 => \N__29894\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101000101"
        )
    port map (
            in0 => \N__29893\,
            in1 => \N__29842\,
            in2 => \N__29873\,
            in3 => \N__29830\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_16_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33281\,
            in1 => \N__33299\,
            in2 => \_gnd_net_\,
            in3 => \N__34843\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50197\,
            ce => \N__29766\,
            sr => \N__49490\
        );

    \phase_controller_inst2.stoper_tr.target_time_17_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34841\,
            in1 => \N__33412\,
            in2 => \_gnd_net_\,
            in3 => \N__33434\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50197\,
            ce => \N__29766\,
            sr => \N__49490\
        );

    \phase_controller_inst2.stoper_tr.target_time_15_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29822\,
            in1 => \N__29792\,
            in2 => \_gnd_net_\,
            in3 => \N__34842\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50197\,
            ce => \N__29766\,
            sr => \N__49490\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__36464\,
            in1 => \N__33707\,
            in2 => \_gnd_net_\,
            in3 => \N__43574\,
            lcout => \current_shift_inst.control_input_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__36386\,
            in1 => \N__33653\,
            in2 => \_gnd_net_\,
            in3 => \N__43572\,
            lcout => \current_shift_inst.control_input_axb_0\,
            ltout => \current_shift_inst.control_input_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_0_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29729\,
            in3 => \N__31768\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50191\,
            ce => 'H',
            sr => \N__49494\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43573\,
            lcout => \current_shift_inst.N_1269_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__43575\,
            in1 => \N__36449\,
            in2 => \_gnd_net_\,
            in3 => \N__33692\,
            lcout => \current_shift_inst.control_input_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__33677\,
            in1 => \N__36434\,
            in2 => \_gnd_net_\,
            in3 => \N__43591\,
            lcout => \current_shift_inst.control_input_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__33746\,
            in1 => \N__36530\,
            in2 => \_gnd_net_\,
            in3 => \N__43592\,
            lcout => \current_shift_inst.control_input_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32065\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__32522\,
            in1 => \N__32551\,
            in2 => \_gnd_net_\,
            in3 => \N__32367\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_axb_4_LC_10_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30101\,
            in2 => \N__30083\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un3_threshold_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \bfn_10_26_0_\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_10_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30056\,
            in2 => \N__30038\,
            in3 => \N__30008\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_0\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_10_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30005\,
            in2 => \N__29987\,
            in3 => \N__29960\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_1\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_10_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29957\,
            in2 => \N__29942\,
            in3 => \N__29909\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_2\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_10_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30413\,
            in2 => \N__30395\,
            in3 => \N__30368\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_3\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_10_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30365\,
            in2 => \N__30347\,
            in3 => \N__30323\,
            lcout => \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_4\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_10_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30320\,
            in2 => \N__30302\,
            in3 => \N__30278\,
            lcout => \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_5\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_10_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30275\,
            in2 => \N__30260\,
            in3 => \N__30236\,
            lcout => \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_6\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_10_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30233\,
            in2 => \N__30218\,
            in3 => \N__30191\,
            lcout => \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \bfn_10_27_0_\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_10_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30188\,
            in2 => \N__30170\,
            in3 => \N__30140\,
            lcout => \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_8\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_10_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32501\,
            in2 => \N__30137\,
            in3 => \N__30110\,
            lcout => \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_9\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_10_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32504\,
            in2 => \N__30683\,
            in3 => \N__30653\,
            lcout => \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_10\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_10_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32502\,
            in2 => \N__30650\,
            in3 => \N__30623\,
            lcout => \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_11\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_10_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32505\,
            in2 => \N__30620\,
            in3 => \N__30593\,
            lcout => \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_12\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_10_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32503\,
            in2 => \N__30590\,
            in3 => \N__30563\,
            lcout => \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_13\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_10_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32506\,
            in2 => \N__30560\,
            in3 => \N__30542\,
            lcout => \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_14\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_10_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__30539\,
            in1 => \N__32291\,
            in2 => \_gnd_net_\,
            in3 => \N__30533\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_2_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__33997\,
            in1 => \N__34738\,
            in2 => \_gnd_net_\,
            in3 => \N__34039\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50288\,
            ce => \N__34337\,
            sr => \N__49413\
        );

    \phase_controller_inst1.stoper_tr.target_time_1_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34757\,
            in1 => \N__32733\,
            in2 => \_gnd_net_\,
            in3 => \N__32179\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50275\,
            ce => \N__34280\,
            sr => \N__49418\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100010000"
        )
    port map (
            in0 => \N__32879\,
            in1 => \N__32900\,
            in2 => \N__30868\,
            in3 => \N__30854\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011101010001"
        )
    port map (
            in0 => \N__32878\,
            in1 => \N__32899\,
            in2 => \N__30869\,
            in3 => \N__30853\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30838\,
            in1 => \N__30815\,
            in2 => \_gnd_net_\,
            in3 => \N__34673\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50264\,
            ce => \N__34322\,
            sr => \N__49427\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30770\,
            in2 => \N__30782\,
            in3 => \N__32713\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_11_8_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30764\,
            in2 => \N__30755\,
            in3 => \N__32680\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30746\,
            in2 => \N__30740\,
            in3 => \N__32662\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32647\,
            in1 => \N__30722\,
            in2 => \N__30731\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30716\,
            in2 => \N__30710\,
            in3 => \N__32632\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32617\,
            in1 => \N__30701\,
            in2 => \N__30695\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34853\,
            in2 => \N__30980\,
            in3 => \N__32602\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34346\,
            in2 => \N__30971\,
            in3 => \N__32587\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_7\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30962\,
            in2 => \N__30956\,
            in3 => \N__32851\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30947\,
            in2 => \N__30941\,
            in3 => \N__32836\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30932\,
            in2 => \N__30926\,
            in3 => \N__32821\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32806\,
            in1 => \N__30914\,
            in2 => \N__30905\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30893\,
            in2 => \N__33008\,
            in3 => \N__32791\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32776\,
            in1 => \N__30887\,
            in2 => \N__30878\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32761\,
            in1 => \N__31070\,
            in2 => \N__31079\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33308\,
            in2 => \N__33374\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_15\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31064\,
            in2 => \N__31052\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_10_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31034\,
            in2 => \N__31028\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31019\,
            in2 => \N__31010\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33920\,
            in2 => \N__33971\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31205\,
            in2 => \N__31214\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30998\,
            in2 => \N__30992\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_30_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31622\,
            in2 => \N__31226\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31217\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101110"
        )
    port map (
            in0 => \N__31145\,
            in1 => \N__31088\,
            in2 => \N__33197\,
            in3 => \N__33174\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__31087\,
            in1 => \N__33195\,
            in2 => \N__33176\,
            in3 => \N__31144\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31173\,
            in1 => \N__31192\,
            in2 => \_gnd_net_\,
            in3 => \N__34746\,
            lcout => \elapsed_time_ns_1_RNI5GPBB_0_27\,
            ltout => \elapsed_time_ns_1_RNI5GPBB_0_27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_27_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__34749\,
            in1 => \_gnd_net_\,
            in2 => \N__31181\,
            in3 => \N__31174\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50219\,
            ce => \N__34261\,
            sr => \N__49464\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31119\,
            in1 => \N__31135\,
            in2 => \_gnd_net_\,
            in3 => \N__34747\,
            lcout => \elapsed_time_ns_1_RNI4FPBB_0_26\,
            ltout => \elapsed_time_ns_1_RNI4FPBB_0_26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_26_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__34748\,
            in1 => \_gnd_net_\,
            in2 => \N__31124\,
            in3 => \N__31120\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50219\,
            ce => \N__34261\,
            sr => \N__49464\
        );

    \phase_controller_inst1.stoper_tr.target_time_31_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32257\,
            in1 => \N__32215\,
            in2 => \_gnd_net_\,
            in3 => \N__34750\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50219\,
            ce => \N__34261\,
            sr => \N__49464\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110011101111"
        )
    port map (
            in0 => \N__31645\,
            in1 => \N__33078\,
            in2 => \N__33113\,
            in3 => \N__31633\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31614\,
            in2 => \_gnd_net_\,
            in3 => \N__31574\,
            lcout => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\,
            ltout => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__31391\,
            in1 => \N__31355\,
            in2 => \N__31334\,
            in3 => \N__31326\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50208\,
            ce => 'H',
            sr => \N__49472\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__34141\,
            in1 => \N__33226\,
            in2 => \N__35171\,
            in3 => \N__32712\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50198\,
            ce => 'H',
            sr => \N__49479\
        );

    \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__31242\,
            in1 => \N__31303\,
            in2 => \_gnd_net_\,
            in3 => \N__31290\,
            lcout => \phase_controller_inst2.stoper_hc.un2_start_0\,
            ltout => \phase_controller_inst2.stoper_hc.un2_start_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.running_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101000111010"
        )
    port map (
            in0 => \N__31304\,
            in1 => \N__31243\,
            in2 => \N__31307\,
            in3 => \N__37657\,
            lcout => \phase_controller_inst2.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50198\,
            ce => 'H',
            sr => \N__49479\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIFU8H_30_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31241\,
            in2 => \_gnd_net_\,
            in3 => \N__37656\,
            lcout => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.start_latched_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31295\,
            lcout => \phase_controller_inst2.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50192\,
            ce => 'H',
            sr => \N__49486\
        );

    \phase_controller_inst1.T45_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31786\,
            in2 => \_gnd_net_\,
            in3 => \N__33457\,
            lcout => \T45_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50192\,
            ce => 'H',
            sr => \N__49486\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31775\,
            in2 => \N__31769\,
            in3 => \N__31767\,
            lcout => \current_shift_inst.control_input_1\,
            ltout => OPEN,
            carryin => \bfn_11_15_0_\,
            carryout => \current_shift_inst.control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33506\,
            in2 => \_gnd_net_\,
            in3 => \N__31730\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_0\,
            carryout => \current_shift_inst.control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33500\,
            in2 => \_gnd_net_\,
            in3 => \N__31718\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_1\,
            carryout => \current_shift_inst.control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33494\,
            in2 => \_gnd_net_\,
            in3 => \N__31706\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_2\,
            carryout => \current_shift_inst.control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33488\,
            in2 => \_gnd_net_\,
            in3 => \N__31694\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_3\,
            carryout => \current_shift_inst.control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33482\,
            in2 => \_gnd_net_\,
            in3 => \N__31679\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_4\,
            carryout => \current_shift_inst.control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33476\,
            in2 => \_gnd_net_\,
            in3 => \N__31664\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_5\,
            carryout => \current_shift_inst.control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35201\,
            in2 => \_gnd_net_\,
            in3 => \N__31649\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_6\,
            carryout => \current_shift_inst.control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31934\,
            in2 => \_gnd_net_\,
            in3 => \N__31919\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_11_16_0_\,
            carryout => \current_shift_inst.control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31916\,
            in2 => \_gnd_net_\,
            in3 => \N__31901\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_8\,
            carryout => \current_shift_inst.control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31898\,
            in3 => \N__31877\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_9\,
            carryout => \current_shift_inst.control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35339\,
            in3 => \N__31865\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_10\,
            carryout => \current_shift_inst.control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35321\,
            in2 => \_gnd_net_\,
            in3 => \N__31850\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_11\,
            carryout => \current_shift_inst.control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35303\,
            in2 => \_gnd_net_\,
            in3 => \N__31835\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_12\,
            carryout => \current_shift_inst.control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35285\,
            in2 => \_gnd_net_\,
            in3 => \N__31820\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_13\,
            carryout => \current_shift_inst.control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35267\,
            in2 => \_gnd_net_\,
            in3 => \N__31805\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_14\,
            carryout => \current_shift_inst.control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35393\,
            in2 => \_gnd_net_\,
            in3 => \N__32036\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_11_17_0_\,
            carryout => \current_shift_inst.control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32564\,
            in2 => \_gnd_net_\,
            in3 => \N__32021\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_16\,
            carryout => \current_shift_inst.control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32573\,
            in2 => \_gnd_net_\,
            in3 => \N__32006\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_17\,
            carryout => \current_shift_inst.control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32003\,
            in2 => \_gnd_net_\,
            in3 => \N__31988\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_18\,
            carryout => \current_shift_inst.control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35462\,
            in2 => \_gnd_net_\,
            in3 => \N__31976\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_19\,
            carryout => \current_shift_inst.control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35747\,
            in2 => \_gnd_net_\,
            in3 => \N__31964\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_20\,
            carryout => \current_shift_inst.control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35729\,
            in2 => \_gnd_net_\,
            in3 => \N__31952\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_21\,
            carryout => \current_shift_inst.control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35702\,
            in2 => \_gnd_net_\,
            in3 => \N__31937\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_22\,
            carryout => \current_shift_inst.control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35534\,
            in2 => \_gnd_net_\,
            in3 => \N__32141\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_11_18_0_\,
            carryout => \current_shift_inst.control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35378\,
            in2 => \_gnd_net_\,
            in3 => \N__32126\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_24\,
            carryout => \current_shift_inst.control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35480\,
            in2 => \_gnd_net_\,
            in3 => \N__32114\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_25\,
            carryout => \current_shift_inst.control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32054\,
            in2 => \_gnd_net_\,
            in3 => \N__32102\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_26\,
            carryout => \current_shift_inst.control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33788\,
            in2 => \_gnd_net_\,
            in3 => \N__32087\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_27\,
            carryout => \current_shift_inst.control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33782\,
            in2 => \_gnd_net_\,
            in3 => \N__32075\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_28\,
            carryout => \current_shift_inst.control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__43516\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32072\,
            lcout => \current_shift_inst.control_input_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__36638\,
            in1 => \N__33800\,
            in2 => \_gnd_net_\,
            in3 => \N__43515\,
            lcout => \current_shift_inst.control_input_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45376\,
            in1 => \N__41055\,
            in2 => \N__42785\,
            in3 => \N__41017\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__43560\,
            in1 => \N__33755\,
            in2 => \_gnd_net_\,
            in3 => \N__36554\,
            lcout => \current_shift_inst.control_input_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__33764\,
            in1 => \N__36569\,
            in2 => \_gnd_net_\,
            in3 => \N__43559\,
            lcout => \current_shift_inst.control_input_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__32555\,
            in1 => \N__32521\,
            in2 => \N__32411\,
            in3 => \N__32309\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D2_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32264\,
            lcout => \il_max_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50287\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D1_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32279\,
            lcout => \il_max_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50287\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.start_timer_hc_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35852\,
            lcout => \delay_measurement_inst.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34054\,
            ce => 'H',
            sr => \N__49405\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35170\,
            in2 => \_gnd_net_\,
            in3 => \N__33230\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32258\,
            in1 => \N__32208\,
            in2 => \_gnd_net_\,
            in3 => \N__34737\,
            lcout => \elapsed_time_ns_1_RNI0CQBB_0_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32178\,
            in1 => \N__32737\,
            in2 => \_gnd_net_\,
            in3 => \N__34736\,
            lcout => \elapsed_time_ns_1_RNIDC91B_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32717\,
            in2 => \N__32690\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_7_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34234\,
            in1 => \N__32681\,
            in2 => \_gnd_net_\,
            in3 => \N__32669\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \N__50251\,
            ce => 'H',
            sr => \N__49419\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__34331\,
            in1 => \N__33209\,
            in2 => \N__32666\,
            in3 => \N__32651\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \N__50251\,
            ce => 'H',
            sr => \N__49419\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34235\,
            in1 => \N__32648\,
            in2 => \_gnd_net_\,
            in3 => \N__32636\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \N__50251\,
            ce => 'H',
            sr => \N__49419\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34332\,
            in1 => \N__32633\,
            in2 => \_gnd_net_\,
            in3 => \N__32621\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \N__50251\,
            ce => 'H',
            sr => \N__49419\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34236\,
            in1 => \N__32618\,
            in2 => \_gnd_net_\,
            in3 => \N__32606\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \N__50251\,
            ce => 'H',
            sr => \N__49419\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34333\,
            in1 => \N__32603\,
            in2 => \_gnd_net_\,
            in3 => \N__32591\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \N__50251\,
            ce => 'H',
            sr => \N__49419\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34237\,
            in1 => \N__32588\,
            in2 => \_gnd_net_\,
            in3 => \N__32576\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \N__50251\,
            ce => 'H',
            sr => \N__49419\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34330\,
            in1 => \N__32852\,
            in2 => \_gnd_net_\,
            in3 => \N__32840\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_12_8_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \N__50239\,
            ce => 'H',
            sr => \N__49428\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34317\,
            in1 => \N__32837\,
            in2 => \_gnd_net_\,
            in3 => \N__32825\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \N__50239\,
            ce => 'H',
            sr => \N__49428\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34327\,
            in1 => \N__32822\,
            in2 => \_gnd_net_\,
            in3 => \N__32810\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \N__50239\,
            ce => 'H',
            sr => \N__49428\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34318\,
            in1 => \N__32807\,
            in2 => \_gnd_net_\,
            in3 => \N__32795\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \N__50239\,
            ce => 'H',
            sr => \N__49428\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34328\,
            in1 => \N__32792\,
            in2 => \_gnd_net_\,
            in3 => \N__32780\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \N__50239\,
            ce => 'H',
            sr => \N__49428\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34319\,
            in1 => \N__32777\,
            in2 => \_gnd_net_\,
            in3 => \N__32765\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \N__50239\,
            ce => 'H',
            sr => \N__49428\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34329\,
            in1 => \N__32762\,
            in2 => \_gnd_net_\,
            in3 => \N__32750\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \N__50239\,
            ce => 'H',
            sr => \N__49428\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34320\,
            in1 => \N__33354\,
            in2 => \_gnd_net_\,
            in3 => \N__32747\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \N__50239\,
            ce => 'H',
            sr => \N__49428\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34230\,
            in1 => \N__33324\,
            in2 => \_gnd_net_\,
            in3 => \N__32996\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_12_9_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \N__50227\,
            ce => 'H',
            sr => \N__49439\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34323\,
            in1 => \N__32985\,
            in2 => \_gnd_net_\,
            in3 => \N__32969\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \N__50227\,
            ce => 'H',
            sr => \N__49439\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34231\,
            in1 => \N__32964\,
            in2 => \_gnd_net_\,
            in3 => \N__32948\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \N__50227\,
            ce => 'H',
            sr => \N__49439\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34324\,
            in1 => \N__32940\,
            in2 => \_gnd_net_\,
            in3 => \N__32924\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \N__50227\,
            ce => 'H',
            sr => \N__49439\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34232\,
            in1 => \N__32919\,
            in2 => \_gnd_net_\,
            in3 => \N__32903\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\,
            clk => \N__50227\,
            ce => 'H',
            sr => \N__49439\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34325\,
            in1 => \N__32898\,
            in2 => \_gnd_net_\,
            in3 => \N__32882\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\,
            clk => \N__50227\,
            ce => 'H',
            sr => \N__49439\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34233\,
            in1 => \N__32877\,
            in2 => \_gnd_net_\,
            in3 => \N__32861\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\,
            clk => \N__50227\,
            ce => 'H',
            sr => \N__49439\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34326\,
            in1 => \N__33956\,
            in2 => \_gnd_net_\,
            in3 => \N__32858\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\,
            clk => \N__50227\,
            ce => 'H',
            sr => \N__49439\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34226\,
            in1 => \N__33936\,
            in2 => \_gnd_net_\,
            in3 => \N__32855\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_12_10_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\,
            clk => \N__50217\,
            ce => 'H',
            sr => \N__49449\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34309\,
            in1 => \N__33196\,
            in2 => \_gnd_net_\,
            in3 => \N__33179\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\,
            clk => \N__50217\,
            ce => 'H',
            sr => \N__49449\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34227\,
            in1 => \N__33175\,
            in2 => \_gnd_net_\,
            in3 => \N__33158\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\,
            clk => \N__50217\,
            ce => 'H',
            sr => \N__49449\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34310\,
            in1 => \N__33153\,
            in2 => \_gnd_net_\,
            in3 => \N__33137\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\,
            clk => \N__50217\,
            ce => 'H',
            sr => \N__49449\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34228\,
            in1 => \N__33132\,
            in2 => \_gnd_net_\,
            in3 => \N__33116\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\,
            clk => \N__50217\,
            ce => 'H',
            sr => \N__49449\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34311\,
            in1 => \N__33111\,
            in2 => \_gnd_net_\,
            in3 => \N__33089\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\,
            clk => \N__50217\,
            ce => 'H',
            sr => \N__49449\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34229\,
            in1 => \N__33079\,
            in2 => \_gnd_net_\,
            in3 => \N__33086\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50217\,
            ce => 'H',
            sr => \N__49449\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34752\,
            in1 => \N__33036\,
            in2 => \_gnd_net_\,
            in3 => \N__33055\,
            lcout => \elapsed_time_ns_1_RNI0AOBB_0_13\,
            ltout => \elapsed_time_ns_1_RNI0AOBB_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_13_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011100010111000"
        )
    port map (
            in0 => \N__33037\,
            in1 => \N__34754\,
            in2 => \N__33011\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50206\,
            ce => \N__34202\,
            sr => \N__49456\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__34753\,
            in1 => \_gnd_net_\,
            in2 => \N__33413\,
            in3 => \N__33427\,
            lcout => \elapsed_time_ns_1_RNI4EOBB_0_17\,
            ltout => \elapsed_time_ns_1_RNI4EOBB_0_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_17_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34756\,
            in2 => \N__33416\,
            in3 => \N__33411\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50206\,
            ce => \N__34202\,
            sr => \N__49456\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101000101"
        )
    port map (
            in0 => \N__33325\,
            in1 => \N__33238\,
            in2 => \N__33359\,
            in3 => \N__33334\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011110010"
        )
    port map (
            in0 => \N__33239\,
            in1 => \N__33355\,
            in2 => \N__33338\,
            in3 => \N__33326\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34751\,
            in1 => \N__33276\,
            in2 => \_gnd_net_\,
            in3 => \N__33292\,
            lcout => \elapsed_time_ns_1_RNI3DOBB_0_16\,
            ltout => \elapsed_time_ns_1_RNI3DOBB_0_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_16_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011100010111000"
        )
    port map (
            in0 => \N__33277\,
            in1 => \N__34755\,
            in2 => \N__33242\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50206\,
            ce => \N__34202\,
            sr => \N__49456\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI3C8N_30_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35011\,
            in2 => \_gnd_net_\,
            in3 => \N__35127\,
            lcout => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1_30_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33212\,
            in3 => \N__35164\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1Z0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_tr_RNO_0_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__34986\,
            in1 => \N__39839\,
            in2 => \N__48065\,
            in3 => \N__48013\,
            lcout => \phase_controller_inst1.start_timer_tr_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__35107\,
            in1 => \N__35012\,
            in2 => \_gnd_net_\,
            in3 => \N__35036\,
            lcout => \phase_controller_inst1.stoper_tr.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36885\,
            in1 => \N__38405\,
            in2 => \_gnd_net_\,
            in3 => \N__48910\,
            lcout => \elapsed_time_ns_1_RNIL73T9_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35013\,
            in2 => \_gnd_net_\,
            in3 => \N__35037\,
            lcout => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35066\,
            in2 => \_gnd_net_\,
            in3 => \N__35091\,
            lcout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1_30_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35067\,
            in2 => \_gnd_net_\,
            in3 => \N__35092\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1Z0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_0_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__34988\,
            in1 => \N__33469\,
            in2 => \N__33458\,
            in3 => \N__39846\,
            lcout => \phase_controller_inst1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50187\,
            ce => 'H',
            sr => \N__49480\
        );

    \phase_controller_inst1.stoper_tr.time_passed_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010001011100010"
        )
    port map (
            in0 => \N__33470\,
            in1 => \N__35169\,
            in2 => \N__35020\,
            in3 => \N__35134\,
            lcout => \phase_controller_inst1.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50187\,
            ce => 'H',
            sr => \N__49480\
        );

    \phase_controller_inst1.state_RNI7NN7_0_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33468\,
            in2 => \_gnd_net_\,
            in3 => \N__33453\,
            lcout => \phase_controller_inst1.state_RNI7NN7Z0Z_0\,
            ltout => \phase_controller_inst1.state_RNI7NN7Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_3_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__35602\,
            in1 => \N__35680\,
            in2 => \N__33437\,
            in3 => \N__33571\,
            lcout => state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50187\,
            ce => 'H',
            sr => \N__49480\
        );

    \phase_controller_inst1.start_timer_hc_RNO_0_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35601\,
            in2 => \_gnd_net_\,
            in3 => \N__35676\,
            lcout => \phase_controller_inst1.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_ns_i_a3_1_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33546\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46894\,
            lcout => state_ns_i_a3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_4_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__46895\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33545\,
            lcout => phase_controller_inst1_state_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50187\,
            ce => 'H',
            sr => \N__49480\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45440\,
            in1 => \N__41519\,
            in2 => \N__42882\,
            in3 => \N__41483\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__43576\,
            in1 => \N__33629\,
            in2 => \_gnd_net_\,
            in3 => \N__36374\,
            lcout => \current_shift_inst.control_input_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__43577\,
            in1 => \N__36362\,
            in2 => \_gnd_net_\,
            in3 => \N__33620\,
            lcout => \current_shift_inst.control_input_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__36335\,
            in1 => \N__33611\,
            in2 => \_gnd_net_\,
            in3 => \N__43578\,
            lcout => \current_shift_inst.control_input_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__43579\,
            in1 => \N__36323\,
            in2 => \_gnd_net_\,
            in3 => \N__33602\,
            lcout => \current_shift_inst.control_input_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__36311\,
            in1 => \N__33593\,
            in2 => \_gnd_net_\,
            in3 => \N__43580\,
            lcout => \current_shift_inst.control_input_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__43581\,
            in1 => \N__36296\,
            in2 => \_gnd_net_\,
            in3 => \N__33722\,
            lcout => \current_shift_inst.control_input_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41179\,
            in2 => \N__41552\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_16_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40886\,
            in2 => \N__37877\,
            in3 => \N__45041\,
            lcout => \current_shift_inst.un38_control_input_5_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__45042\,
            in1 => \N__42431\,
            in2 => \N__36767\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un38_control_input_5_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36611\,
            in2 => \N__42605\,
            in3 => \N__33641\,
            lcout => \current_shift_inst.un38_control_input_0_s0_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42435\,
            in2 => \N__33638\,
            in3 => \N__33623\,
            lcout => \current_shift_inst.un38_control_input_0_s0_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35369\,
            in2 => \N__42606\,
            in3 => \N__33614\,
            lcout => \current_shift_inst.un38_control_input_0_s0_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42439\,
            in2 => \N__35192\,
            in3 => \N__33605\,
            lcout => \current_shift_inst.un38_control_input_0_s0_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35363\,
            in2 => \N__42607\,
            in3 => \N__33596\,
            lcout => \current_shift_inst.un38_control_input_0_s0_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42482\,
            in2 => \N__35432\,
            in3 => \N__33584\,
            lcout => \current_shift_inst.un38_control_input_0_s0_8\,
            ltout => OPEN,
            carryin => \bfn_12_17_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40793\,
            in2 => \N__42716\,
            in3 => \N__33713\,
            lcout => \current_shift_inst.un38_control_input_0_s0_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42486\,
            in2 => \N__35450\,
            in3 => \N__33710\,
            lcout => \current_shift_inst.un38_control_input_0_s0_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35546\,
            in2 => \N__42717\,
            in3 => \N__33695\,
            lcout => \current_shift_inst.un38_control_input_0_s0_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42490\,
            in2 => \N__35357\,
            in3 => \N__33680\,
            lcout => \current_shift_inst.un38_control_input_0_s0_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37760\,
            in2 => \N__42718\,
            in3 => \N__33665\,
            lcout => \current_shift_inst.un38_control_input_0_s0_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42494\,
            in2 => \N__35420\,
            in3 => \N__33662\,
            lcout => \current_shift_inst.un38_control_input_0_s0_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35258\,
            in2 => \N__42719\,
            in3 => \N__33659\,
            lcout => \current_shift_inst.un38_control_input_0_s0_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42563\,
            in2 => \N__35510\,
            in3 => \N__33656\,
            lcout => \current_shift_inst.un38_control_input_0_s0_16\,
            ltout => OPEN,
            carryin => \bfn_12_18_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35411\,
            in2 => \N__42778\,
            in3 => \N__33773\,
            lcout => \current_shift_inst.un38_control_input_0_s0_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42567\,
            in2 => \N__35519\,
            in3 => \N__33770\,
            lcout => \current_shift_inst.un38_control_input_0_s0_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35405\,
            in2 => \N__42779\,
            in3 => \N__33767\,
            lcout => \current_shift_inst.un38_control_input_0_s0_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42571\,
            in2 => \N__37796\,
            in3 => \N__33758\,
            lcout => \current_shift_inst.un38_control_input_0_s0_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37832\,
            in2 => \N__42780\,
            in3 => \N__33749\,
            lcout => \current_shift_inst.un38_control_input_0_s0_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42575\,
            in2 => \N__35441\,
            in3 => \N__33734\,
            lcout => \current_shift_inst.un38_control_input_0_s0_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35525\,
            in2 => \N__42781\,
            in3 => \N__33731\,
            lcout => \current_shift_inst.un38_control_input_0_s0_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42579\,
            in2 => \N__35495\,
            in3 => \N__33728\,
            lcout => \current_shift_inst.un38_control_input_0_s0_24\,
            ltout => OPEN,
            carryin => \bfn_12_19_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42224\,
            in2 => \N__42782\,
            in3 => \N__33725\,
            lcout => \current_shift_inst.un38_control_input_0_s0_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42583\,
            in2 => \N__35717\,
            in3 => \N__33812\,
            lcout => \current_shift_inst.un38_control_input_0_s0_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37859\,
            in2 => \N__42783\,
            in3 => \N__33809\,
            lcout => \current_shift_inst.un38_control_input_0_s0_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42587\,
            in2 => \N__37889\,
            in3 => \N__33806\,
            lcout => \current_shift_inst.un38_control_input_0_s0_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35501\,
            in2 => \N__42784\,
            in3 => \N__33803\,
            lcout => \current_shift_inst.un38_control_input_0_s0_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42591\,
            in2 => \N__41321\,
            in3 => \N__33794\,
            lcout => \current_shift_inst.un38_control_input_0_s0_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001101010011"
        )
    port map (
            in0 => \N__40766\,
            in1 => \N__36623\,
            in2 => \N__43590\,
            in3 => \N__33791\,
            lcout => \current_shift_inst.control_input_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43571\,
            lcout => \current_shift_inst.control_input_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.start_timer_s1_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__35574\,
            in1 => \N__36749\,
            in2 => \_gnd_net_\,
            in3 => \N__35628\,
            lcout => \current_shift_inst.start_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50171\,
            ce => 'H',
            sr => \N__49509\
        );

    \phase_controller_inst1.S1_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35629\,
            lcout => s1_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50171\,
            ce => 'H',
            sr => \N__49509\
        );

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49571\,
            lcout => \pll_inst.red_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_hc_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35853\,
            lcout => \delay_measurement_inst.stop_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34055\,
            ce => 'H',
            sr => \N__49406\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34739\,
            in1 => \N__34404\,
            in2 => \_gnd_net_\,
            in3 => \N__34374\,
            lcout => \elapsed_time_ns_1_RNIKJ91B_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__33996\,
            in1 => \N__34038\,
            in2 => \_gnd_net_\,
            in3 => \N__34740\,
            lcout => \elapsed_time_ns_1_RNIED91B_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34741\,
            in1 => \N__34909\,
            in2 => \_gnd_net_\,
            in3 => \N__34881\,
            lcout => \elapsed_time_ns_1_RNIJI91B_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__33954\,
            in1 => \N__33937\,
            in2 => \N__33842\,
            in3 => \N__34922\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__34921\,
            in1 => \N__33955\,
            in2 => \N__33941\,
            in3 => \N__33838\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_25_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34778\,
            in1 => \N__33908\,
            in2 => \_gnd_net_\,
            in3 => \N__33878\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50253\,
            ce => \N__34262\,
            sr => \N__49420\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34954\,
            in1 => \N__33823\,
            in2 => \_gnd_net_\,
            in3 => \N__34776\,
            lcout => \elapsed_time_ns_1_RNI2DPBB_0_24\,
            ltout => \elapsed_time_ns_1_RNI2DPBB_0_24_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_24_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__34777\,
            in1 => \_gnd_net_\,
            in2 => \N__34958\,
            in3 => \N__34955\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50253\,
            ce => \N__34262\,
            sr => \N__49420\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34905\,
            in1 => \N__34889\,
            in2 => \_gnd_net_\,
            in3 => \N__34780\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50253\,
            ce => \N__34262\,
            sr => \N__49420\
        );

    \phase_controller_inst1.stoper_tr.target_time_8_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34779\,
            in1 => \N__34408\,
            in2 => \_gnd_net_\,
            in3 => \N__34385\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50253\,
            ce => \N__34262\,
            sr => \N__49420\
        );

    \phase_controller_inst1.stoper_hc.target_time_31_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40277\,
            in1 => \N__36685\,
            in2 => \_gnd_net_\,
            in3 => \N__48856\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50241\,
            ce => \N__49832\,
            sr => \N__49429\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__46988\,
            in1 => \N__43991\,
            in2 => \N__44296\,
            in3 => \N__49833\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50229\,
            ce => 'H',
            sr => \N__49440\
        );

    \phase_controller_inst2.stoper_hc.target_time_10_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38345\,
            in1 => \N__48921\,
            in2 => \_gnd_net_\,
            in3 => \N__36788\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50220\,
            ce => \N__47862\,
            sr => \N__49450\
        );

    \phase_controller_inst2.stoper_hc.target_time_22_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48920\,
            in1 => \N__47756\,
            in2 => \_gnd_net_\,
            in3 => \N__47727\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50220\,
            ce => \N__47862\,
            sr => \N__49450\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101110"
        )
    port map (
            in0 => \N__35180\,
            in1 => \N__34076\,
            in2 => \N__36023\,
            in3 => \N__36000\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__34075\,
            in1 => \N__36021\,
            in2 => \N__36002\,
            in3 => \N__35179\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_23_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__47655\,
            in1 => \N__48922\,
            in2 => \_gnd_net_\,
            in3 => \N__47675\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50209\,
            ce => \N__47861\,
            sr => \N__49457\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36987\,
            in1 => \N__38285\,
            in2 => \_gnd_net_\,
            in3 => \N__48880\,
            lcout => \elapsed_time_ns_1_RNIUVBN9_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.running_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000101110"
        )
    port map (
            in0 => \N__35108\,
            in1 => \N__35168\,
            in2 => \N__35021\,
            in3 => \N__35135\,
            lcout => \phase_controller_inst1.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50199\,
            ce => 'H',
            sr => \N__49465\
        );

    \delay_measurement_inst.delay_hc_timer.running_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__35817\,
            in1 => \N__35801\,
            in2 => \_gnd_net_\,
            in3 => \N__35864\,
            lcout => \delay_measurement_inst.delay_hc_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50199\,
            ce => 'H',
            sr => \N__49465\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__36169\,
            in1 => \N__35096\,
            in2 => \N__35078\,
            in3 => \N__37116\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50199\,
            ce => 'H',
            sr => \N__49465\
        );

    \phase_controller_inst1.start_timer_tr_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110111001100"
        )
    port map (
            in0 => \N__35051\,
            in1 => \N__35045\,
            in2 => \N__46916\,
            in3 => \N__35038\,
            lcout => \phase_controller_inst1.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50199\,
            ce => 'H',
            sr => \N__49465\
        );

    \phase_controller_inst1.stoper_tr.start_latched_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__35039\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50199\,
            ce => 'H',
            sr => \N__49465\
        );

    \phase_controller_inst1.state_1_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__34987\,
            in1 => \N__39845\,
            in2 => \_gnd_net_\,
            in3 => \N__47969\,
            lcout => \phase_controller_inst1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50199\,
            ce => 'H',
            sr => \N__49465\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__36277\,
            in1 => \N__35976\,
            in2 => \N__35243\,
            in3 => \N__35252\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__35251\,
            in1 => \N__36276\,
            in2 => \N__35981\,
            in3 => \N__35239\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_24_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__40586\,
            in1 => \N__40628\,
            in2 => \_gnd_net_\,
            in3 => \N__48935\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50193\,
            ce => \N__47860\,
            sr => \N__49473\
        );

    \phase_controller_inst2.stoper_hc.target_time_25_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48931\,
            in1 => \N__40678\,
            in2 => \_gnd_net_\,
            in3 => \N__40697\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50193\,
            ce => \N__47860\,
            sr => \N__49473\
        );

    \phase_controller_inst2.stoper_hc.target_time_31_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40276\,
            in1 => \N__36692\,
            in2 => \_gnd_net_\,
            in3 => \N__48936\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50193\,
            ce => \N__47860\,
            sr => \N__49473\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011111011"
        )
    port map (
            in0 => \N__35218\,
            in1 => \N__36247\,
            in2 => \N__36062\,
            in3 => \N__35227\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_30_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001100"
        )
    port map (
            in0 => \N__36246\,
            in1 => \N__36057\,
            in2 => \N__35231\,
            in3 => \N__35219\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_30_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__35777\,
            in1 => \_gnd_net_\,
            in2 => \N__48938\,
            in3 => \N__39175\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50193\,
            ce => \N__47860\,
            sr => \N__49473\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__36473\,
            in1 => \N__35210\,
            in2 => \_gnd_net_\,
            in3 => \N__43582\,
            lcout => \current_shift_inst.control_input_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001010101"
        )
    port map (
            in0 => \N__41060\,
            in1 => \N__42771\,
            in2 => \N__41018\,
            in3 => \N__45442\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45441\,
            in1 => \N__41141\,
            in2 => \N__42883\,
            in3 => \N__41108\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__43073\,
            in1 => \N__45443\,
            in2 => \N__43034\,
            in3 => \N__42772\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__41377\,
            in1 => \N__45438\,
            in2 => \N__42720\,
            in3 => \N__41345\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100011011"
        )
    port map (
            in0 => \N__43551\,
            in1 => \N__36422\,
            in2 => \N__35348\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.control_input_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__36413\,
            in1 => \N__35327\,
            in2 => \_gnd_net_\,
            in3 => \N__43552\,
            lcout => \current_shift_inst.control_input_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__43553\,
            in1 => \N__35312\,
            in2 => \_gnd_net_\,
            in3 => \N__36404\,
            lcout => \current_shift_inst.control_input_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__35294\,
            in1 => \N__43554\,
            in2 => \_gnd_net_\,
            in3 => \N__36395\,
            lcout => \current_shift_inst.control_input_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__43555\,
            in1 => \N__36587\,
            in2 => \_gnd_net_\,
            in3 => \N__35276\,
            lcout => \current_shift_inst.control_input_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__42502\,
            in1 => \N__45439\,
            in2 => \N__41440\,
            in3 => \N__41405\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__45437\,
            in1 => \N__42498\,
            in2 => \N__40949\,
            in3 => \N__40984\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__45435\,
            in1 => \N__42504\,
            in2 => \N__39980\,
            in3 => \N__40009\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__42503\,
            in1 => \N__45431\,
            in2 => \N__41615\,
            in3 => \N__41573\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45432\,
            in1 => \N__42511\,
            in2 => \N__41974\,
            in3 => \N__41927\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__40010\,
            in1 => \N__45436\,
            in2 => \N__42721\,
            in3 => \N__39978\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__45433\,
            in1 => \N__41897\,
            in2 => \N__41087\,
            in3 => \N__42512\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__41857\,
            in1 => \N__45434\,
            in2 => \N__42722\,
            in3 => \N__41813\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__35399\,
            in1 => \N__36578\,
            in2 => \_gnd_net_\,
            in3 => \N__43556\,
            lcout => \current_shift_inst.control_input_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__36656\,
            in1 => \N__35384\,
            in2 => \_gnd_net_\,
            in3 => \N__43558\,
            lcout => \current_shift_inst.control_input_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45277\,
            in1 => \N__44777\,
            in2 => \N__42861\,
            in3 => \N__44816\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__36665\,
            in1 => \N__35540\,
            in2 => \_gnd_net_\,
            in3 => \N__43557\,
            lcout => \current_shift_inst.control_input_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45279\,
            in1 => \N__43138\,
            in2 => \N__42862\,
            in3 => \N__43097\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45280\,
            in1 => \N__42723\,
            in2 => \N__41792\,
            in3 => \N__41753\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45278\,
            in1 => \N__41252\,
            in2 => \N__42863\,
            in3 => \N__41210\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__42730\,
            in1 => \N__45281\,
            in2 => \N__42209\,
            in3 => \N__42170\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45282\,
            in1 => \N__39949\,
            in2 => \N__42864\,
            in3 => \N__39908\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__35486\,
            in1 => \N__36647\,
            in2 => \_gnd_net_\,
            in3 => \N__43567\,
            lcout => \current_shift_inst.control_input_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__43561\,
            in1 => \N__35468\,
            in2 => \_gnd_net_\,
            in3 => \N__36518\,
            lcout => \current_shift_inst.control_input_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__35753\,
            in1 => \N__36506\,
            in2 => \_gnd_net_\,
            in3 => \N__43562\,
            lcout => \current_shift_inst.control_input_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010100110101"
        )
    port map (
            in0 => \N__36491\,
            in1 => \N__35735\,
            in2 => \N__43589\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.control_input_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45283\,
            in1 => \N__41303\,
            in2 => \N__42865\,
            in3 => \N__39599\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__35708\,
            in1 => \N__36482\,
            in2 => \_gnd_net_\,
            in3 => \N__43566\,
            lcout => \current_shift_inst.control_input_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_2_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__35623\,
            in1 => \N__48047\,
            in2 => \N__35690\,
            in3 => \N__48020\,
            lcout => \phase_controller_inst1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50175\,
            ce => 'H',
            sr => \N__49503\
        );

    \phase_controller_inst1.T01_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35641\,
            in2 => \_gnd_net_\,
            in3 => \N__35624\,
            lcout => \T01_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50175\,
            ce => 'H',
            sr => \N__49503\
        );

    \current_shift_inst.timer_s1.running_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__36727\,
            in1 => \N__36752\,
            in2 => \_gnd_net_\,
            in3 => \N__37948\,
            lcout => \current_shift_inst.timer_s1.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50172\,
            ce => 'H',
            sr => \N__49507\
        );

    \current_shift_inst.stop_timer_s1_LC_13_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101100"
        )
    port map (
            in0 => \N__36751\,
            in1 => \N__36728\,
            in2 => \N__35630\,
            in3 => \N__35575\,
            lcout => \current_shift_inst.stop_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50172\,
            ce => 'H',
            sr => \N__49507\
        );

    \current_shift_inst.timer_s1.running_RNII51H_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37943\,
            in2 => \_gnd_net_\,
            in3 => \N__36725\,
            lcout => \current_shift_inst.timer_s1.N_162_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.S2_LC_13_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39856\,
            lcout => s2_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50165\,
            ce => 'H',
            sr => \N__49539\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__35796\,
            in1 => \N__35831\,
            in2 => \_gnd_net_\,
            in3 => \N__35860\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_199_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_30_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__35769\,
            in1 => \N__39179\,
            in2 => \_gnd_net_\,
            in3 => \N__48908\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50276\,
            ce => \N__49806\,
            sr => \N__49407\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35826\,
            lcout => \delay_measurement_inst.delay_hc_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__47448\,
            in1 => \N__50354\,
            in2 => \N__40679\,
            in3 => \N__39173\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__35932\,
            in1 => \N__38814\,
            in2 => \_gnd_net_\,
            in3 => \N__48877\,
            lcout => \elapsed_time_ns_1_RNI02CN9_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__35827\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35797\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_198_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48876\,
            in1 => \N__35773\,
            in2 => \_gnd_net_\,
            in3 => \N__39174\,
            lcout => \elapsed_time_ns_1_RNIV2EN9_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48855\,
            in1 => \N__38512\,
            in2 => \_gnd_net_\,
            in3 => \N__37152\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50254\,
            ce => \N__49805\,
            sr => \N__49421\
        );

    \phase_controller_inst1.stoper_hc.target_time_13_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48854\,
            in1 => \N__35928\,
            in2 => \_gnd_net_\,
            in3 => \N__38816\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50254\,
            ce => \N__49805\,
            sr => \N__49421\
        );

    \phase_controller_inst2.stoper_hc.target_time_13_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48888\,
            in1 => \N__35933\,
            in2 => \_gnd_net_\,
            in3 => \N__38815\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50242\,
            ce => \N__47866\,
            sr => \N__49430\
        );

    \phase_controller_inst2.stoper_hc.target_time_11_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36991\,
            in1 => \N__38284\,
            in2 => \_gnd_net_\,
            in3 => \N__48890\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50242\,
            ce => \N__47866\,
            sr => \N__49430\
        );

    \phase_controller_inst2.stoper_hc.target_time_15_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48889\,
            in1 => \N__44055\,
            in2 => \_gnd_net_\,
            in3 => \N__44035\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50242\,
            ce => \N__47866\,
            sr => \N__49430\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35912\,
            in2 => \N__37124\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_11_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36223\,
            in1 => \N__37087\,
            in2 => \_gnd_net_\,
            in3 => \N__35900\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \N__50230\,
            ce => 'H',
            sr => \N__49441\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__36227\,
            in1 => \N__37054\,
            in2 => \N__35897\,
            in3 => \N__35882\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \N__50230\,
            ce => 'H',
            sr => \N__49441\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36224\,
            in1 => \N__37027\,
            in2 => \_gnd_net_\,
            in3 => \N__35879\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \N__50230\,
            ce => 'H',
            sr => \N__49441\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36228\,
            in1 => \N__37399\,
            in2 => \_gnd_net_\,
            in3 => \N__35876\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \N__50230\,
            ce => 'H',
            sr => \N__49441\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36225\,
            in1 => \N__37369\,
            in2 => \_gnd_net_\,
            in3 => \N__35873\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \N__50230\,
            ce => 'H',
            sr => \N__49441\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36229\,
            in1 => \N__37327\,
            in2 => \_gnd_net_\,
            in3 => \N__35960\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \N__50230\,
            ce => 'H',
            sr => \N__49441\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36226\,
            in1 => \N__37306\,
            in2 => \_gnd_net_\,
            in3 => \N__35957\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \N__50230\,
            ce => 'H',
            sr => \N__49441\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36196\,
            in1 => \N__37258\,
            in2 => \_gnd_net_\,
            in3 => \N__35954\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_14_12_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \N__50221\,
            ce => 'H',
            sr => \N__49451\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36173\,
            in1 => \N__37219\,
            in2 => \_gnd_net_\,
            in3 => \N__35951\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \N__50221\,
            ce => 'H',
            sr => \N__49451\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36193\,
            in1 => \N__37180\,
            in2 => \_gnd_net_\,
            in3 => \N__35948\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \N__50221\,
            ce => 'H',
            sr => \N__49451\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36174\,
            in1 => \N__37594\,
            in2 => \_gnd_net_\,
            in3 => \N__35945\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \N__50221\,
            ce => 'H',
            sr => \N__49451\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36194\,
            in1 => \N__37570\,
            in2 => \_gnd_net_\,
            in3 => \N__35942\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \N__50221\,
            ce => 'H',
            sr => \N__49451\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36175\,
            in1 => \N__37534\,
            in2 => \_gnd_net_\,
            in3 => \N__35939\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \N__50221\,
            ce => 'H',
            sr => \N__49451\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36195\,
            in1 => \N__37495\,
            in2 => \_gnd_net_\,
            in3 => \N__35936\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \N__50221\,
            ce => 'H',
            sr => \N__49451\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36176\,
            in1 => \N__39115\,
            in2 => \_gnd_net_\,
            in3 => \N__36041\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \N__50221\,
            ce => 'H',
            sr => \N__49451\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36161\,
            in1 => \N__39100\,
            in2 => \_gnd_net_\,
            in3 => \N__36038\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_14_13_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \N__50210\,
            ce => 'H',
            sr => \N__49458\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36165\,
            in1 => \N__36833\,
            in2 => \_gnd_net_\,
            in3 => \N__36035\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \N__50210\,
            ce => 'H',
            sr => \N__49458\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36162\,
            in1 => \N__36850\,
            in2 => \_gnd_net_\,
            in3 => \N__36032\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \N__50210\,
            ce => 'H',
            sr => \N__49458\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36166\,
            in1 => \N__36933\,
            in2 => \_gnd_net_\,
            in3 => \N__36029\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \N__50210\,
            ce => 'H',
            sr => \N__49458\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36163\,
            in1 => \N__36960\,
            in2 => \_gnd_net_\,
            in3 => \N__36026\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\,
            clk => \N__50210\,
            ce => 'H',
            sr => \N__49458\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36167\,
            in1 => \N__36022\,
            in2 => \_gnd_net_\,
            in3 => \N__36005\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\,
            clk => \N__50210\,
            ce => 'H',
            sr => \N__49458\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36164\,
            in1 => \N__36001\,
            in2 => \_gnd_net_\,
            in3 => \N__35984\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\,
            clk => \N__50210\,
            ce => 'H',
            sr => \N__49458\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36168\,
            in1 => \N__35980\,
            in2 => \_gnd_net_\,
            in3 => \N__35963\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\,
            clk => \N__50210\,
            ce => 'H',
            sr => \N__49458\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36220\,
            in1 => \N__36278\,
            in2 => \_gnd_net_\,
            in3 => \N__36263\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_14_14_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\,
            clk => \N__50200\,
            ce => 'H',
            sr => \N__49466\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36216\,
            in1 => \N__44614\,
            in2 => \_gnd_net_\,
            in3 => \N__36260\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\,
            clk => \N__50200\,
            ce => 'H',
            sr => \N__49466\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36221\,
            in1 => \N__44589\,
            in2 => \_gnd_net_\,
            in3 => \N__36257\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\,
            clk => \N__50200\,
            ce => 'H',
            sr => \N__49466\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36217\,
            in1 => \N__45526\,
            in2 => \_gnd_net_\,
            in3 => \N__36254\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\,
            clk => \N__50200\,
            ce => 'H',
            sr => \N__49466\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36222\,
            in1 => \N__45505\,
            in2 => \_gnd_net_\,
            in3 => \N__36251\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\,
            clk => \N__50200\,
            ce => 'H',
            sr => \N__49466\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36218\,
            in1 => \N__36248\,
            in2 => \_gnd_net_\,
            in3 => \N__36233\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\,
            clk => \N__50200\,
            ce => 'H',
            sr => \N__49466\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__36061\,
            in1 => \N__36219\,
            in2 => \_gnd_net_\,
            in3 => \N__36065\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50200\,
            ce => 'H',
            sr => \N__49466\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45083\,
            in2 => \N__41180\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_15_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40899\,
            in2 => \N__40862\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42745\,
            in2 => \N__36707\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36599\,
            in2 => \N__42876\,
            in3 => \N__36377\,
            lcout => \current_shift_inst.un38_control_input_0_s1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42749\,
            in2 => \N__41456\,
            in3 => \N__36365\,
            lcout => \current_shift_inst.un38_control_input_0_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39245\,
            in2 => \N__42877\,
            in3 => \N__36353\,
            lcout => \current_shift_inst.un38_control_input_0_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42753\,
            in2 => \N__36350\,
            in3 => \N__36326\,
            lcout => \current_shift_inst.un38_control_input_0_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37781\,
            in2 => \N__42878\,
            in3 => \N__36314\,
            lcout => \current_shift_inst.un38_control_input_0_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42608\,
            in2 => \N__41156\,
            in3 => \N__36299\,
            lcout => \current_shift_inst.un38_control_input_0_s1_8\,
            ltout => OPEN,
            carryin => \bfn_14_16_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40778\,
            in2 => \N__42792\,
            in3 => \N__36281\,
            lcout => \current_shift_inst.un38_control_input_0_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42612\,
            in2 => \N__37628\,
            in3 => \N__36467\,
            lcout => \current_shift_inst.un38_control_input_0_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37766\,
            in2 => \N__42793\,
            in3 => \N__36452\,
            lcout => \current_shift_inst.un38_control_input_0_s1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42616\,
            in2 => \N__37775\,
            in3 => \N__36437\,
            lcout => \current_shift_inst.un38_control_input_0_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37634\,
            in2 => \N__42794\,
            in3 => \N__36425\,
            lcout => \current_shift_inst.un38_control_input_0_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42620\,
            in2 => \N__37619\,
            in3 => \N__36416\,
            lcout => \current_shift_inst.un38_control_input_0_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37610\,
            in2 => \N__42795\,
            in3 => \N__36407\,
            lcout => \current_shift_inst.un38_control_input_0_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42796\,
            in2 => \N__39881\,
            in3 => \N__36398\,
            lcout => \current_shift_inst.un38_control_input_0_s1_16\,
            ltout => OPEN,
            carryin => \bfn_14_17_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37850\,
            in2 => \N__42889\,
            in3 => \N__36389\,
            lcout => \current_shift_inst.un38_control_input_0_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42800\,
            in2 => \N__37739\,
            in3 => \N__36581\,
            lcout => \current_shift_inst.un38_control_input_0_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37745\,
            in2 => \N__42890\,
            in3 => \N__36572\,
            lcout => \current_shift_inst.un38_control_input_0_s1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42804\,
            in2 => \N__37805\,
            in3 => \N__36557\,
            lcout => \current_shift_inst.un38_control_input_0_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37751\,
            in2 => \N__42891\,
            in3 => \N__36542\,
            lcout => \current_shift_inst.un38_control_input_0_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42808\,
            in2 => \N__36539\,
            in3 => \N__36521\,
            lcout => \current_shift_inst.un38_control_input_0_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37724\,
            in2 => \N__42892\,
            in3 => \N__36509\,
            lcout => \current_shift_inst.un38_control_input_0_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39260\,
            in2 => \N__42893\,
            in3 => \N__36494\,
            lcout => \current_shift_inst.un38_control_input_0_s1_24\,
            ltout => OPEN,
            carryin => \bfn_14_18_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42815\,
            in2 => \N__37907\,
            in3 => \N__36485\,
            lcout => \current_shift_inst.un38_control_input_0_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37895\,
            in2 => \N__42894\,
            in3 => \N__36476\,
            lcout => \current_shift_inst.un38_control_input_0_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42819\,
            in2 => \N__37823\,
            in3 => \N__36659\,
            lcout => \current_shift_inst.un38_control_input_0_s1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37811\,
            in2 => \N__42895\,
            in3 => \N__36650\,
            lcout => \current_shift_inst.un38_control_input_0_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42823\,
            in2 => \N__37844\,
            in3 => \N__36641\,
            lcout => \current_shift_inst.un38_control_input_0_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42825\,
            in2 => \N__42968\,
            in3 => \N__36629\,
            lcout => \current_shift_inst.un38_control_input_0_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__45284\,
            in1 => \N__42824\,
            in2 => \_gnd_net_\,
            in3 => \N__36626\,
            lcout => \current_shift_inst.un38_control_input_0_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__42786\,
            in1 => \N__45223\,
            in2 => \N__42034\,
            in3 => \N__41998\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44997\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50178\,
            ce => \N__44954\,
            sr => \N__49495\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__42787\,
            in1 => \N__45224\,
            in2 => \N__42035\,
            in3 => \N__41999\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI00M61_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45222\,
            in1 => \N__42788\,
            in2 => \N__42146\,
            in3 => \N__42109\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIEOIK_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__36750\,
            in1 => \N__37947\,
            in2 => \_gnd_net_\,
            in3 => \N__36726\,
            lcout => \current_shift_inst.timer_s1.N_163_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45335\,
            in1 => \N__42145\,
            in2 => \N__42910\,
            in3 => \N__42113\,
            lcout => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_19_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44105\,
            in1 => \N__48906\,
            in2 => \_gnd_net_\,
            in3 => \N__44126\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50299\,
            ce => \N__47872\,
            sr => \N__49398\
        );

    \phase_controller_inst2.stoper_hc.target_time_1_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__46487\,
            in1 => \N__46340\,
            in2 => \_gnd_net_\,
            in3 => \N__48907\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50289\,
            ce => \N__47871\,
            sr => \N__49402\
        );

    \phase_controller_inst2.stoper_hc.target_time_21_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39770\,
            in1 => \N__39799\,
            in2 => \_gnd_net_\,
            in3 => \N__48879\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50277\,
            ce => \N__47869\,
            sr => \N__49408\
        );

    \phase_controller_inst2.stoper_hc.target_time_12_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__40043\,
            in1 => \N__40073\,
            in2 => \_gnd_net_\,
            in3 => \N__48878\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50277\,
            ce => \N__47869\,
            sr => \N__49408\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40275\,
            in1 => \N__36684\,
            in2 => \_gnd_net_\,
            in3 => \N__48776\,
            lcout => \elapsed_time_ns_1_RNI04EN9_0_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__38796\,
            in1 => \N__44027\,
            in2 => \N__47792\,
            in3 => \N__47079\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__47720\,
            in1 => \N__47643\,
            in2 => \N__40627\,
            in3 => \N__39767\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__36818\,
            in1 => \N__36803\,
            in2 => \N__36812\,
            in3 => \N__36809\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__44094\,
            in1 => \N__47907\,
            in2 => \N__43938\,
            in3 => \N__47199\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44059\,
            in1 => \N__44028\,
            in2 => \_gnd_net_\,
            in3 => \N__48777\,
            lcout => \elapsed_time_ns_1_RNI24CN9_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48778\,
            in1 => \N__38505\,
            in2 => \_gnd_net_\,
            in3 => \N__37156\,
            lcout => \elapsed_time_ns_1_RNII43T9_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__38273\,
            in1 => \N__38336\,
            in2 => \N__38400\,
            in3 => \N__40064\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__40322\,
            in1 => \N__38504\,
            in2 => \N__36797\,
            in3 => \N__36794\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__47508\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40118\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38337\,
            in1 => \N__48884\,
            in2 => \_gnd_net_\,
            in3 => \N__36781\,
            lcout => \elapsed_time_ns_1_RNITUBN9_0_10\,
            ltout => \elapsed_time_ns_1_RNITUBN9_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_10_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__48885\,
            in1 => \_gnd_net_\,
            in2 => \N__36770\,
            in3 => \N__38338\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50255\,
            ce => \N__49791\,
            sr => \N__49422\
        );

    \phase_controller_inst1.stoper_hc.target_time_9_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36893\,
            in1 => \N__38399\,
            in2 => \_gnd_net_\,
            in3 => \N__48887\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50255\,
            ce => \N__49791\,
            sr => \N__49422\
        );

    \phase_controller_inst1.stoper_hc.target_time_11_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__48886\,
            in1 => \_gnd_net_\,
            in2 => \N__36995\,
            in3 => \N__38274\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50255\,
            ce => \N__49791\,
            sr => \N__49422\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001100"
        )
    port map (
            in0 => \N__36940\,
            in1 => \N__36917\,
            in2 => \N__36965\,
            in3 => \N__36902\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__36901\,
            in1 => \N__36964\,
            in2 => \N__36944\,
            in3 => \N__36916\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_20_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43889\,
            in1 => \N__43919\,
            in2 => \_gnd_net_\,
            in3 => \N__48905\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50243\,
            ce => \N__47867\,
            sr => \N__49431\
        );

    \phase_controller_inst2.stoper_hc.target_time_8_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__40124\,
            in1 => \N__48891\,
            in2 => \_gnd_net_\,
            in3 => \N__40097\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50243\,
            ce => \N__47867\,
            sr => \N__49431\
        );

    \phase_controller_inst2.stoper_hc.target_time_7_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48893\,
            in1 => \N__47520\,
            in2 => \_gnd_net_\,
            in3 => \N__47543\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50243\,
            ce => \N__47867\,
            sr => \N__49431\
        );

    \phase_controller_inst2.stoper_hc.target_time_9_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38404\,
            in1 => \N__48892\,
            in2 => \_gnd_net_\,
            in3 => \N__36892\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50243\,
            ce => \N__47867\,
            sr => \N__49431\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__36832\,
            in1 => \N__47891\,
            in2 => \N__36869\,
            in3 => \N__36849\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011001111"
        )
    port map (
            in0 => \N__47890\,
            in1 => \N__36868\,
            in2 => \N__36851\,
            in3 => \N__36831\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_3_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43724\,
            in1 => \N__46460\,
            in2 => \_gnd_net_\,
            in3 => \N__48903\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50231\,
            ce => \N__47863\,
            sr => \N__49442\
        );

    \phase_controller_inst2.stoper_hc.target_time_4_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48901\,
            in1 => \N__43700\,
            in2 => \_gnd_net_\,
            in3 => \N__46384\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50231\,
            ce => \N__47863\,
            sr => \N__49442\
        );

    \phase_controller_inst2.stoper_hc.target_time_5_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40331\,
            in1 => \N__40301\,
            in2 => \_gnd_net_\,
            in3 => \N__48904\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50231\,
            ce => \N__47863\,
            sr => \N__49442\
        );

    \phase_controller_inst2.stoper_hc.target_time_6_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48902\,
            in1 => \N__38516\,
            in2 => \_gnd_net_\,
            in3 => \N__37157\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50231\,
            ce => \N__47863\,
            sr => \N__49442\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37094\,
            in2 => \N__37136\,
            in3 => \N__37117\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_15_13_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39056\,
            in2 => \N__37073\,
            in3 => \N__37088\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37064\,
            in2 => \N__37040\,
            in3 => \N__37058\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37031\,
            in1 => \N__37013\,
            in2 => \N__37007\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37400\,
            in1 => \N__37376\,
            in2 => \N__37385\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37370\,
            in1 => \N__37355\,
            in2 => \N__37349\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37313\,
            in2 => \N__37340\,
            in3 => \N__37328\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37307\,
            in1 => \N__37292\,
            in2 => \N__37283\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_7\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37274\,
            in2 => \N__37244\,
            in3 => \N__37262\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_15_14_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37232\,
            in2 => \N__37205\,
            in3 => \N__37220\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37196\,
            in2 => \N__37166\,
            in3 => \N__37184\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37604\,
            in2 => \N__37580\,
            in3 => \N__37595\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37571\,
            in1 => \N__37556\,
            in2 => \N__37544\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37535\,
            in1 => \N__39062\,
            in2 => \N__37520\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37508\,
            in2 => \N__37481\,
            in3 => \N__37496\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39131\,
            in2 => \N__39080\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_15\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37472\,
            in2 => \N__37463\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_15_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37451\,
            in2 => \N__37442\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37427\,
            in2 => \N__37415\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_20\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37718\,
            in2 => \N__37706\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_22\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44573\,
            in2 => \N__44639\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_24\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45491\,
            in2 => \N__44564\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_26\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_30_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37691\,
            in2 => \N__37679\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_28\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37664\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__41537\,
            in1 => \N__42857\,
            in2 => \N__42083\,
            in3 => \N__45383\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45378\,
            in1 => \N__40985\,
            in2 => \N__42902\,
            in3 => \N__40948\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__41926\,
            in1 => \N__42858\,
            in2 => \N__41975\,
            in3 => \N__45384\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45385\,
            in1 => \N__42859\,
            in2 => \N__41441\,
            in3 => \N__41401\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__43069\,
            in1 => \N__45377\,
            in2 => \N__43029\,
            in3 => \N__42854\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41048\,
            lcout => \current_shift_inst.un4_control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__41344\,
            in1 => \N__42856\,
            in2 => \N__41381\,
            in3 => \N__45382\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \N__42855\,
            in1 => \N__44776\,
            in2 => \N__45447\,
            in3 => \N__44812\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__42076\,
            in1 => \N__45407\,
            in2 => \N__42896\,
            in3 => \N__41536\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010101111"
        )
    port map (
            in0 => \N__41638\,
            in1 => \N__42827\,
            in2 => \N__45451\,
            in3 => \N__41675\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001111"
        )
    port map (
            in0 => \N__42831\,
            in1 => \N__41809\,
            in2 => \N__41858\,
            in3 => \N__45410\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__45409\,
            in1 => \N__42826\,
            in2 => \N__41752\,
            in3 => \N__41791\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI25021_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001111"
        )
    port map (
            in0 => \N__42832\,
            in1 => \N__43090\,
            in2 => \N__43139\,
            in3 => \N__45414\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41369\,
            lcout => \current_shift_inst.un4_control_input_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__41896\,
            in1 => \N__45408\,
            in2 => \N__42897\,
            in3 => \N__41079\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__45415\,
            in1 => \N__42833\,
            in2 => \N__42169\,
            in3 => \N__42208\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__41671\,
            in1 => \N__45390\,
            in2 => \N__41639\,
            in3 => \N__42839\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \N__42837\,
            in1 => \N__39656\,
            in2 => \N__45449\,
            in3 => \N__39619\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__39443\,
            in1 => \N__42838\,
            in2 => \N__39710\,
            in3 => \N__45396\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001111"
        )
    port map (
            in0 => \N__42841\,
            in1 => \N__41725\,
            in2 => \N__45448\,
            in3 => \N__41708\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__41707\,
            in1 => \N__45386\,
            in2 => \N__41726\,
            in3 => \N__42840\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40002\,
            lcout => \current_shift_inst.un4_control_input_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__42285\,
            in1 => \N__42842\,
            in2 => \N__42263\,
            in3 => \N__45391\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45392\,
            in1 => \N__41302\,
            in2 => \N__42898\,
            in3 => \N__39597\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41948\,
            lcout => \current_shift_inst.un4_control_input_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__45221\,
            in1 => \N__42847\,
            in2 => \N__39442\,
            in3 => \N__39700\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__39699\,
            in1 => \N__45219\,
            in2 => \_gnd_net_\,
            in3 => \N__39435\,
            lcout => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__45218\,
            in1 => \N__40817\,
            in2 => \N__40909\,
            in3 => \N__40847\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40964\,
            lcout => \current_shift_inst.un4_control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45220\,
            in1 => \N__42846\,
            in2 => \N__39655\,
            in3 => \N__39618\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41418\,
            lcout => \current_shift_inst.un4_control_input_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41231\,
            lcout => \current_shift_inst.un4_control_input_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42245\,
            lcout => \current_shift_inst.un4_control_input_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41771\,
            lcout => \current_shift_inst.un4_control_input_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIUKI8_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37949\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.timer_s1.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41660\,
            lcout => \current_shift_inst.un4_control_input_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.counter_0_LC_16_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38178\,
            in1 => \N__43854\,
            in2 => \_gnd_net_\,
            in3 => \N__37922\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_16_5_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            clk => \N__50317\,
            ce => \N__38055\,
            sr => \N__49394\
        );

    \delay_measurement_inst.delay_hc_timer.counter_1_LC_16_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38162\,
            in1 => \N__43824\,
            in2 => \_gnd_net_\,
            in3 => \N__37919\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            clk => \N__50317\,
            ce => \N__38055\,
            sr => \N__49394\
        );

    \delay_measurement_inst.delay_hc_timer.counter_2_LC_16_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38179\,
            in1 => \N__38559\,
            in2 => \_gnd_net_\,
            in3 => \N__37916\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            clk => \N__50317\,
            ce => \N__38055\,
            sr => \N__49394\
        );

    \delay_measurement_inst.delay_hc_timer.counter_3_LC_16_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38163\,
            in1 => \N__38530\,
            in2 => \_gnd_net_\,
            in3 => \N__37913\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            clk => \N__50317\,
            ce => \N__38055\,
            sr => \N__49394\
        );

    \delay_measurement_inst.delay_hc_timer.counter_4_LC_16_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38180\,
            in1 => \N__38472\,
            in2 => \_gnd_net_\,
            in3 => \N__37910\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            clk => \N__50317\,
            ce => \N__38055\,
            sr => \N__49394\
        );

    \delay_measurement_inst.delay_hc_timer.counter_5_LC_16_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38164\,
            in1 => \N__38445\,
            in2 => \_gnd_net_\,
            in3 => \N__37976\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            clk => \N__50317\,
            ce => \N__38055\,
            sr => \N__49394\
        );

    \delay_measurement_inst.delay_hc_timer.counter_6_LC_16_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38181\,
            in1 => \N__38419\,
            in2 => \_gnd_net_\,
            in3 => \N__37973\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            clk => \N__50317\,
            ce => \N__38055\,
            sr => \N__49394\
        );

    \delay_measurement_inst.delay_hc_timer.counter_7_LC_16_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38165\,
            in1 => \N__38359\,
            in2 => \_gnd_net_\,
            in3 => \N__37970\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            clk => \N__50317\,
            ce => \N__38055\,
            sr => \N__49394\
        );

    \delay_measurement_inst.delay_hc_timer.counter_8_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38161\,
            in1 => \N__38301\,
            in2 => \_gnd_net_\,
            in3 => \N__37967\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_16_6_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            clk => \N__50310\,
            ce => \N__38054\,
            sr => \N__49395\
        );

    \delay_measurement_inst.delay_hc_timer.counter_9_LC_16_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38173\,
            in1 => \N__38238\,
            in2 => \_gnd_net_\,
            in3 => \N__37964\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            clk => \N__50310\,
            ce => \N__38054\,
            sr => \N__49395\
        );

    \delay_measurement_inst.delay_hc_timer.counter_10_LC_16_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38158\,
            in1 => \N__38212\,
            in2 => \_gnd_net_\,
            in3 => \N__37961\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            clk => \N__50310\,
            ce => \N__38054\,
            sr => \N__49395\
        );

    \delay_measurement_inst.delay_hc_timer.counter_11_LC_16_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38170\,
            in1 => \N__38773\,
            in2 => \_gnd_net_\,
            in3 => \N__37958\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            clk => \N__50310\,
            ce => \N__38054\,
            sr => \N__49395\
        );

    \delay_measurement_inst.delay_hc_timer.counter_12_LC_16_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38159\,
            in1 => \N__38748\,
            in2 => \_gnd_net_\,
            in3 => \N__37955\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            clk => \N__50310\,
            ce => \N__38054\,
            sr => \N__49395\
        );

    \delay_measurement_inst.delay_hc_timer.counter_13_LC_16_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38171\,
            in1 => \N__38721\,
            in2 => \_gnd_net_\,
            in3 => \N__37952\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            clk => \N__50310\,
            ce => \N__38054\,
            sr => \N__49395\
        );

    \delay_measurement_inst.delay_hc_timer.counter_14_LC_16_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38160\,
            in1 => \N__38695\,
            in2 => \_gnd_net_\,
            in3 => \N__38006\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            clk => \N__50310\,
            ce => \N__38054\,
            sr => \N__49395\
        );

    \delay_measurement_inst.delay_hc_timer.counter_15_LC_16_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38172\,
            in1 => \N__38673\,
            in2 => \_gnd_net_\,
            in3 => \N__38003\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            clk => \N__50310\,
            ce => \N__38054\,
            sr => \N__49395\
        );

    \delay_measurement_inst.delay_hc_timer.counter_16_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38154\,
            in1 => \N__38640\,
            in2 => \_gnd_net_\,
            in3 => \N__38000\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_16_7_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            clk => \N__50300\,
            ce => \N__38056\,
            sr => \N__49399\
        );

    \delay_measurement_inst.delay_hc_timer.counter_17_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38166\,
            in1 => \N__38616\,
            in2 => \_gnd_net_\,
            in3 => \N__37997\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            clk => \N__50300\,
            ce => \N__38056\,
            sr => \N__49399\
        );

    \delay_measurement_inst.delay_hc_timer.counter_18_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38155\,
            in1 => \N__38586\,
            in2 => \_gnd_net_\,
            in3 => \N__37994\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            clk => \N__50300\,
            ce => \N__38056\,
            sr => \N__49399\
        );

    \delay_measurement_inst.delay_hc_timer.counter_19_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38167\,
            in1 => \N__39048\,
            in2 => \_gnd_net_\,
            in3 => \N__37991\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            clk => \N__50300\,
            ce => \N__38056\,
            sr => \N__49399\
        );

    \delay_measurement_inst.delay_hc_timer.counter_20_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38156\,
            in1 => \N__39024\,
            in2 => \_gnd_net_\,
            in3 => \N__37988\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            clk => \N__50300\,
            ce => \N__38056\,
            sr => \N__49399\
        );

    \delay_measurement_inst.delay_hc_timer.counter_21_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38168\,
            in1 => \N__38991\,
            in2 => \_gnd_net_\,
            in3 => \N__37985\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            clk => \N__50300\,
            ce => \N__38056\,
            sr => \N__49399\
        );

    \delay_measurement_inst.delay_hc_timer.counter_22_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38157\,
            in1 => \N__38962\,
            in2 => \_gnd_net_\,
            in3 => \N__37982\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            clk => \N__50300\,
            ce => \N__38056\,
            sr => \N__49399\
        );

    \delay_measurement_inst.delay_hc_timer.counter_23_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38169\,
            in1 => \N__38932\,
            in2 => \_gnd_net_\,
            in3 => \N__37979\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            clk => \N__50300\,
            ce => \N__38056\,
            sr => \N__49399\
        );

    \delay_measurement_inst.delay_hc_timer.counter_24_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38174\,
            in1 => \N__38901\,
            in2 => \_gnd_net_\,
            in3 => \N__38198\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_16_8_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            clk => \N__50290\,
            ce => \N__38057\,
            sr => \N__49403\
        );

    \delay_measurement_inst.delay_hc_timer.counter_25_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38182\,
            in1 => \N__38877\,
            in2 => \_gnd_net_\,
            in3 => \N__38195\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            clk => \N__50290\,
            ce => \N__38057\,
            sr => \N__49403\
        );

    \delay_measurement_inst.delay_hc_timer.counter_26_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38175\,
            in1 => \N__38853\,
            in2 => \_gnd_net_\,
            in3 => \N__38192\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            clk => \N__50290\,
            ce => \N__38057\,
            sr => \N__49403\
        );

    \delay_measurement_inst.delay_hc_timer.counter_27_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38183\,
            in1 => \N__39198\,
            in2 => \_gnd_net_\,
            in3 => \N__38189\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            clk => \N__50290\,
            ce => \N__38057\,
            sr => \N__49403\
        );

    \delay_measurement_inst.delay_hc_timer.counter_28_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38176\,
            in1 => \N__38833\,
            in2 => \_gnd_net_\,
            in3 => \N__38186\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_28\,
            clk => \N__50290\,
            ce => \N__38057\,
            sr => \N__49403\
        );

    \delay_measurement_inst.delay_hc_timer.counter_29_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__39217\,
            in1 => \N__38177\,
            in2 => \_gnd_net_\,
            in3 => \N__38060\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50290\,
            ce => \N__38057\,
            sr => \N__49403\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43861\,
            in2 => \N__38566\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\,
            ltout => OPEN,
            carryin => \bfn_16_9_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__50278\,
            ce => \N__43792\,
            sr => \N__49409\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38536\,
            in2 => \N__43838\,
            in3 => \N__38009\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__50278\,
            ce => \N__43792\,
            sr => \N__49409\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38567\,
            in2 => \N__38479\,
            in3 => \N__38540\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__50278\,
            ce => \N__43792\,
            sr => \N__49409\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38537\,
            in2 => \N__38452\,
            in3 => \N__38483\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__50278\,
            ce => \N__43792\,
            sr => \N__49409\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38425\,
            in2 => \N__38480\,
            in3 => \N__38456\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__50278\,
            ce => \N__43792\,
            sr => \N__49409\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38365\,
            in2 => \N__38453\,
            in3 => \N__38429\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__50278\,
            ce => \N__43792\,
            sr => \N__49409\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38426\,
            in2 => \N__38314\,
            in3 => \N__38369\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__50278\,
            ce => \N__43792\,
            sr => \N__49409\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38366\,
            in2 => \N__38251\,
            in3 => \N__38318\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__50278\,
            ce => \N__43792\,
            sr => \N__49409\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38218\,
            in2 => \N__38315\,
            in3 => \N__38255\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\,
            ltout => OPEN,
            carryin => \bfn_16_10_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__50265\,
            ce => \N__43801\,
            sr => \N__49414\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38779\,
            in2 => \N__38252\,
            in3 => \N__38222\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__50265\,
            ce => \N__43801\,
            sr => \N__49414\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38219\,
            in2 => \N__38755\,
            in3 => \N__38783\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__50265\,
            ce => \N__43801\,
            sr => \N__49414\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38780\,
            in2 => \N__38728\,
            in3 => \N__38759\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__50265\,
            ce => \N__43801\,
            sr => \N__49414\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38701\,
            in2 => \N__38756\,
            in3 => \N__38732\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__50265\,
            ce => \N__43801\,
            sr => \N__49414\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38674\,
            in2 => \N__38729\,
            in3 => \N__38705\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__50265\,
            ce => \N__43801\,
            sr => \N__49414\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38702\,
            in2 => \N__38651\,
            in3 => \N__38681\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__50265\,
            ce => \N__43801\,
            sr => \N__49414\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38617\,
            in2 => \N__38678\,
            in3 => \N__38654\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__50265\,
            ce => \N__43801\,
            sr => \N__49414\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38650\,
            in2 => \N__38593\,
            in3 => \N__38624\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\,
            ltout => OPEN,
            carryin => \bfn_16_11_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__50256\,
            ce => \N__43800\,
            sr => \N__49423\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39049\,
            in2 => \N__38621\,
            in3 => \N__38597\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__50256\,
            ce => \N__43800\,
            sr => \N__49423\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39025\,
            in2 => \N__38594\,
            in3 => \N__38570\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__50256\,
            ce => \N__43800\,
            sr => \N__49423\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39050\,
            in2 => \N__39002\,
            in3 => \N__39032\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__50256\,
            ce => \N__43800\,
            sr => \N__49423\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38968\,
            in2 => \N__39029\,
            in3 => \N__39005\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__50256\,
            ce => \N__43800\,
            sr => \N__49423\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39001\,
            in2 => \N__38944\,
            in3 => \N__38972\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__50256\,
            ce => \N__43800\,
            sr => \N__49423\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38969\,
            in2 => \N__38914\,
            in3 => \N__38948\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__50256\,
            ce => \N__43800\,
            sr => \N__49423\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38878\,
            in2 => \N__38945\,
            in3 => \N__38918\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__50256\,
            ce => \N__43800\,
            sr => \N__49423\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38854\,
            in2 => \N__38915\,
            in3 => \N__38885\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\,
            ltout => OPEN,
            carryin => \bfn_16_12_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__50244\,
            ce => \N__43805\,
            sr => \N__49432\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39199\,
            in2 => \N__38882\,
            in3 => \N__38858\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__50244\,
            ce => \N__43805\,
            sr => \N__49432\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38855\,
            in2 => \N__38837\,
            in3 => \N__38819\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__50244\,
            ce => \N__43805\,
            sr => \N__49432\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39221\,
            in2 => \N__39203\,
            in3 => \N__39137\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__50244\,
            ce => \N__43805\,
            sr => \N__49432\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39134\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50244\,
            ce => \N__43805\,
            sr => \N__49432\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101110"
        )
    port map (
            in0 => \N__39071\,
            in1 => \N__47048\,
            in2 => \N__39125\,
            in3 => \N__39099\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__47047\,
            in1 => \N__39124\,
            in2 => \N__39101\,
            in3 => \N__39070\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_17_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48926\,
            in1 => \N__47209\,
            in2 => \_gnd_net_\,
            in3 => \N__47234\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50232\,
            ce => \N__47864\,
            sr => \N__49443\
        );

    \phase_controller_inst2.stoper_hc.target_time_14_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47111\,
            in1 => \N__47091\,
            in2 => \_gnd_net_\,
            in3 => \N__48930\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50232\,
            ce => \N__47864\,
            sr => \N__49443\
        );

    \phase_controller_inst2.stoper_hc.target_time_2_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__43748\,
            in1 => \_gnd_net_\,
            in2 => \N__48937\,
            in3 => \N__46421\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50232\,
            ce => \N__47864\,
            sr => \N__49443\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43068\,
            lcout => \current_shift_inst.un4_control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41598\,
            lcout => \current_shift_inst.un4_control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001111"
        )
    port map (
            in0 => \N__42887\,
            in1 => \N__39904\,
            in2 => \N__39953\,
            in3 => \N__45455\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42021\,
            lcout => \current_shift_inst.un4_control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__41518\,
            in1 => \N__44898\,
            in2 => \_gnd_net_\,
            in3 => \N__41472\,
            lcout => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41517\,
            lcout => \current_shift_inst.un4_control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__41133\,
            in1 => \N__45454\,
            in2 => \N__42909\,
            in3 => \N__41104\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI68O61_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41132\,
            lcout => \current_shift_inst.un4_control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40916\,
            in2 => \N__45482\,
            in3 => \N__45480\,
            lcout => \current_shift_inst.un4_control_input1_2\,
            ltout => OPEN,
            carryin => \bfn_16_15_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39509\,
            in2 => \_gnd_net_\,
            in3 => \N__39233\,
            lcout => \current_shift_inst.un4_control_input1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_1\,
            carryout => \current_shift_inst.un4_control_input_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39230\,
            in2 => \_gnd_net_\,
            in3 => \N__39224\,
            lcout => \current_shift_inst.un4_control_input1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_2\,
            carryout => \current_shift_inst.un4_control_input_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39335\,
            in2 => \_gnd_net_\,
            in3 => \N__39329\,
            lcout => \current_shift_inst.un4_control_input1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_3\,
            carryout => \current_shift_inst.un4_control_input_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39326\,
            in2 => \_gnd_net_\,
            in3 => \N__39320\,
            lcout => \current_shift_inst.un4_control_input1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_4\,
            carryout => \current_shift_inst.un4_control_input_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39317\,
            in2 => \_gnd_net_\,
            in3 => \N__39311\,
            lcout => \current_shift_inst.un4_control_input1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_5\,
            carryout => \current_shift_inst.un4_control_input_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39308\,
            in2 => \_gnd_net_\,
            in3 => \N__39302\,
            lcout => \current_shift_inst.un4_control_input1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_6\,
            carryout => \current_shift_inst.un4_control_input_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39299\,
            in2 => \_gnd_net_\,
            in3 => \N__39293\,
            lcout => \current_shift_inst.un4_control_input1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_7\,
            carryout => \current_shift_inst.un4_control_input_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42923\,
            in3 => \N__39290\,
            lcout => \current_shift_inst.un4_control_input1_10\,
            ltout => OPEN,
            carryin => \bfn_16_16_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39287\,
            in2 => \_gnd_net_\,
            in3 => \N__39275\,
            lcout => \current_shift_inst.un4_control_input1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_9\,
            carryout => \current_shift_inst.un4_control_input_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44741\,
            in2 => \_gnd_net_\,
            in3 => \N__39272\,
            lcout => \current_shift_inst.un4_control_input1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_10\,
            carryout => \current_shift_inst.un4_control_input_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39269\,
            in2 => \_gnd_net_\,
            in3 => \N__39263\,
            lcout => \current_shift_inst.un4_control_input1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_11\,
            carryout => \current_shift_inst.un4_control_input_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42047\,
            in2 => \_gnd_net_\,
            in3 => \N__39416\,
            lcout => \current_shift_inst.un4_control_input1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_12\,
            carryout => \current_shift_inst.un4_control_input_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39413\,
            in2 => \_gnd_net_\,
            in3 => \N__39404\,
            lcout => \current_shift_inst.un4_control_input1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_13\,
            carryout => \current_shift_inst.un4_control_input_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39401\,
            in2 => \_gnd_net_\,
            in3 => \N__39389\,
            lcout => \current_shift_inst.un4_control_input1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_14\,
            carryout => \current_shift_inst.un4_control_input_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39386\,
            in2 => \_gnd_net_\,
            in3 => \N__39374\,
            lcout => \current_shift_inst.un4_control_input1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_15\,
            carryout => \current_shift_inst.un4_control_input_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41864\,
            in2 => \_gnd_net_\,
            in3 => \N__39371\,
            lcout => \current_shift_inst.un4_control_input1_18\,
            ltout => OPEN,
            carryin => \bfn_16_17_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39368\,
            in2 => \_gnd_net_\,
            in3 => \N__39359\,
            lcout => \current_shift_inst.un4_control_input1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_17\,
            carryout => \current_shift_inst.un4_control_input_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40019\,
            in2 => \_gnd_net_\,
            in3 => \N__39356\,
            lcout => \current_shift_inst.un4_control_input1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_18\,
            carryout => \current_shift_inst.un4_control_input_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41684\,
            in3 => \N__39353\,
            lcout => \current_shift_inst.un4_control_input1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_19\,
            carryout => \current_shift_inst.un4_control_input_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39350\,
            in2 => \_gnd_net_\,
            in3 => \N__39338\,
            lcout => \current_shift_inst.un4_control_input1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_20\,
            carryout => \current_shift_inst.un4_control_input_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39476\,
            in2 => \_gnd_net_\,
            in3 => \N__39470\,
            lcout => \current_shift_inst.un4_control_input1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_21\,
            carryout => \current_shift_inst.un4_control_input_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41903\,
            in2 => \_gnd_net_\,
            in3 => \N__39467\,
            lcout => \current_shift_inst.un4_control_input1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_22\,
            carryout => \current_shift_inst.un4_control_input_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39500\,
            in2 => \_gnd_net_\,
            in3 => \N__39464\,
            lcout => \current_shift_inst.un4_control_input1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_23\,
            carryout => \current_shift_inst.un4_control_input_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39461\,
            in2 => \_gnd_net_\,
            in3 => \N__39452\,
            lcout => \current_shift_inst.un4_control_input1_26\,
            ltout => OPEN,
            carryin => \bfn_16_18_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41258\,
            in2 => \_gnd_net_\,
            in3 => \N__39449\,
            lcout => \current_shift_inst.un4_control_input1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_25\,
            carryout => \current_shift_inst.un4_control_input_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39719\,
            in2 => \_gnd_net_\,
            in3 => \N__39446\,
            lcout => \current_shift_inst.un4_control_input1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_26\,
            carryout => \current_shift_inst.un4_control_input_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39674\,
            in2 => \_gnd_net_\,
            in3 => \N__39422\,
            lcout => \current_shift_inst.un4_control_input1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_27\,
            carryout => \current_shift_inst.un4_control_input_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39665\,
            in2 => \_gnd_net_\,
            in3 => \N__39419\,
            lcout => \current_shift_inst.un4_control_input1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_28\,
            carryout => \current_shift_inst.un4_control_input1_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39512\,
            lcout => \current_shift_inst.un4_control_input1_31_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42131\,
            lcout => \current_shift_inst.un4_control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39938\,
            lcout => \current_shift_inst.un4_control_input_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44732\,
            in2 => \N__45760\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_3\,
            ltout => OPEN,
            carryin => \bfn_16_19_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            clk => \N__50184\,
            ce => \N__44957\,
            sr => \N__49487\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45791\,
            in2 => \N__45730\,
            in3 => \N__39494\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            clk => \N__50184\,
            ce => \N__44957\,
            sr => \N__49487\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45697\,
            in2 => \N__45761\,
            in3 => \N__39491\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            clk => \N__50184\,
            ce => \N__44957\,
            sr => \N__49487\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45667\,
            in2 => \N__45731\,
            in3 => \N__39488\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            clk => \N__50184\,
            ce => \N__44957\,
            sr => \N__49487\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45637\,
            in2 => \N__45701\,
            in3 => \N__39485\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            clk => \N__50184\,
            ce => \N__44957\,
            sr => \N__49487\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45607\,
            in2 => \N__45671\,
            in3 => \N__39482\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            clk => \N__50184\,
            ce => \N__44957\,
            sr => \N__49487\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45577\,
            in2 => \N__45641\,
            in3 => \N__39479\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            clk => \N__50184\,
            ce => \N__44957\,
            sr => \N__49487\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46057\,
            in2 => \N__45611\,
            in3 => \N__39539\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            clk => \N__50184\,
            ce => \N__44957\,
            sr => \N__49487\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46024\,
            in2 => \N__45581\,
            in3 => \N__39536\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_11\,
            ltout => OPEN,
            carryin => \bfn_16_20_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            clk => \N__50182\,
            ce => \N__44956\,
            sr => \N__49491\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46000\,
            in2 => \N__46061\,
            in3 => \N__39533\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            clk => \N__50182\,
            ce => \N__44956\,
            sr => \N__49491\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46025\,
            in2 => \N__45976\,
            in3 => \N__39530\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            clk => \N__50182\,
            ce => \N__44956\,
            sr => \N__49491\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46001\,
            in2 => \N__45946\,
            in3 => \N__39527\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            clk => \N__50182\,
            ce => \N__44956\,
            sr => \N__49491\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45916\,
            in2 => \N__45977\,
            in3 => \N__39524\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            clk => \N__50182\,
            ce => \N__44956\,
            sr => \N__49491\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45889\,
            in2 => \N__45947\,
            in3 => \N__39521\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            clk => \N__50182\,
            ce => \N__44956\,
            sr => \N__49491\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45917\,
            in2 => \N__45862\,
            in3 => \N__39518\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            clk => \N__50182\,
            ce => \N__44956\,
            sr => \N__49491\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45820\,
            in2 => \N__45893\,
            in3 => \N__39515\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            clk => \N__50182\,
            ce => \N__44956\,
            sr => \N__49491\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46297\,
            in2 => \N__45863\,
            in3 => \N__39566\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_19\,
            ltout => OPEN,
            carryin => \bfn_16_21_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            clk => \N__50179\,
            ce => \N__44955\,
            sr => \N__49496\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46270\,
            in2 => \N__45824\,
            in3 => \N__39563\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            clk => \N__50179\,
            ce => \N__44955\,
            sr => \N__49496\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46243\,
            in2 => \N__46301\,
            in3 => \N__39560\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            clk => \N__50179\,
            ce => \N__44955\,
            sr => \N__49496\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46271\,
            in2 => \N__46216\,
            in3 => \N__39557\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            clk => \N__50179\,
            ce => \N__44955\,
            sr => \N__49496\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46186\,
            in2 => \N__46247\,
            in3 => \N__39554\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            clk => \N__50179\,
            ce => \N__44955\,
            sr => \N__49496\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46162\,
            in2 => \N__46217\,
            in3 => \N__39551\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            clk => \N__50179\,
            ce => \N__44955\,
            sr => \N__49496\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46187\,
            in2 => \N__46138\,
            in3 => \N__39548\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            clk => \N__50179\,
            ce => \N__44955\,
            sr => \N__49496\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46163\,
            in2 => \N__46099\,
            in3 => \N__39545\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            clk => \N__50179\,
            ce => \N__44955\,
            sr => \N__49496\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46777\,
            in2 => \N__46139\,
            in3 => \N__39542\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_27\,
            ltout => OPEN,
            carryin => \bfn_16_22_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            clk => \N__50177\,
            ce => \N__44953\,
            sr => \N__49498\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46747\,
            in2 => \N__46100\,
            in3 => \N__39731\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            clk => \N__50177\,
            ce => \N__44953\,
            sr => \N__49498\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46721\,
            in2 => \N__46781\,
            in3 => \N__39728\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            clk => \N__50177\,
            ce => \N__44953\,
            sr => \N__49498\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46571\,
            in2 => \N__46751\,
            in3 => \N__39725\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\,
            clk => \N__50177\,
            ce => \N__44953\,
            sr => \N__49498\
        );

    \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39722\,
            lcout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39641\,
            lcout => \current_shift_inst.un4_control_input_1_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39690\,
            lcout => \current_shift_inst.un4_control_input_1_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_16_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42188\,
            lcout => \current_shift_inst.un4_control_input_1_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__39642\,
            in1 => \N__45399\,
            in2 => \_gnd_net_\,
            in3 => \N__39623\,
            lcout => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__41274\,
            in1 => \N__45398\,
            in2 => \_gnd_net_\,
            in3 => \N__39598\,
            lcout => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41843\,
            lcout => \current_shift_inst.un4_control_input_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44929\,
            in1 => \N__40008\,
            in2 => \_gnd_net_\,
            in3 => \N__39979\,
            lcout => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__39939\,
            in1 => \N__44930\,
            in2 => \_gnd_net_\,
            in3 => \N__39903\,
            lcout => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__41209\,
            in1 => \N__42888\,
            in2 => \N__41251\,
            in3 => \N__45400\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISST11_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45397\,
            in1 => \N__42255\,
            in2 => \_gnd_net_\,
            in3 => \N__42286\,
            lcout => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.T23_LC_16_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39811\,
            in2 => \_gnd_net_\,
            in3 => \N__39863\,
            lcout => \T23_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50169\,
            ce => 'H',
            sr => \N__49529\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_17_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__39792\,
            in1 => \N__39768\,
            in2 => \_gnd_net_\,
            in3 => \N__48689\,
            lcout => \elapsed_time_ns_1_RNIV1DN9_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_21_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__39800\,
            in1 => \N__39769\,
            in2 => \_gnd_net_\,
            in3 => \N__48827\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50311\,
            ce => \N__49834\,
            sr => \N__49396\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46379\,
            in1 => \N__43692\,
            in2 => \_gnd_net_\,
            in3 => \N__48828\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50311\,
            ce => \N__49834\,
            sr => \N__49396\
        );

    \phase_controller_inst1.stoper_hc.target_time_12_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__40035\,
            in1 => \N__40072\,
            in2 => \_gnd_net_\,
            in3 => \N__48674\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50301\,
            ce => \N__49792\,
            sr => \N__49400\
        );

    \phase_controller_inst1.stoper_hc.target_time_8_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48673\,
            in1 => \N__40089\,
            in2 => \_gnd_net_\,
            in3 => \N__40120\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50301\,
            ce => \N__49792\,
            sr => \N__49400\
        );

    \phase_controller_inst1.stoper_hc.target_time_5_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40324\,
            in1 => \N__40293\,
            in2 => \_gnd_net_\,
            in3 => \N__48677\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50301\,
            ce => \N__49792\,
            sr => \N__49400\
        );

    \phase_controller_inst1.stoper_hc.target_time_1_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48672\,
            in1 => \N__46483\,
            in2 => \_gnd_net_\,
            in3 => \N__46335\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50301\,
            ce => \N__49792\,
            sr => \N__49400\
        );

    \phase_controller_inst1.stoper_hc.target_time_3_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43716\,
            in1 => \N__46448\,
            in2 => \_gnd_net_\,
            in3 => \N__48676\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50301\,
            ce => \N__49792\,
            sr => \N__49400\
        );

    \phase_controller_inst1.stoper_hc.target_time_2_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46413\,
            in1 => \N__43740\,
            in2 => \_gnd_net_\,
            in3 => \N__48675\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50301\,
            ce => \N__49792\,
            sr => \N__49400\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__40093\,
            in1 => \N__40119\,
            in2 => \_gnd_net_\,
            in3 => \N__48667\,
            lcout => \elapsed_time_ns_1_RNIK63T9_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_30_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100011001110"
        )
    port map (
            in0 => \N__40358\,
            in1 => \N__44660\,
            in2 => \N__44692\,
            in3 => \N__40343\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__40039\,
            in1 => \N__40065\,
            in2 => \_gnd_net_\,
            in3 => \N__48665\,
            lcout => \elapsed_time_ns_1_RNIV0CN9_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110011101111"
        )
    port map (
            in0 => \N__40357\,
            in1 => \N__44659\,
            in2 => \N__44693\,
            in3 => \N__40342\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__40297\,
            in1 => \N__40323\,
            in2 => \_gnd_net_\,
            in3 => \N__48666\,
            lcout => \elapsed_time_ns_1_RNIH33T9_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__40265\,
            in1 => \N__40232\,
            in2 => \N__40220\,
            in3 => \N__47012\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__40578\,
            in1 => \_gnd_net_\,
            in2 => \N__40208\,
            in3 => \N__40622\,
            lcout => \elapsed_time_ns_1_RNI25DN9_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40193\,
            in2 => \N__40205\,
            in3 => \N__44292\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_17_10_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44266\,
            in1 => \N__40187\,
            in2 => \N__40178\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44242\,
            in1 => \N__40169\,
            in2 => \N__40160\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40139\,
            in2 => \N__40151\,
            in3 => \N__44227\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44212\,
            in1 => \N__40133\,
            in2 => \N__40508\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44197\,
            in1 => \N__40496\,
            in2 => \N__40484\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47489\,
            in2 => \N__40472\,
            in3 => \N__44182\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44167\,
            in1 => \N__40463\,
            in2 => \N__40451\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_7\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40439\,
            in2 => \N__40427\,
            in3 => \N__44152\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_17_11_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44407\,
            in1 => \N__40418\,
            in2 => \N__40406\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40397\,
            in2 => \N__40385\,
            in3 => \N__44392\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40376\,
            in2 => \N__40367\,
            in3 => \N__44378\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44356\,
            in1 => \N__40532\,
            in2 => \N__40547\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47060\,
            in2 => \N__40526\,
            in3 => \N__44341\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44012\,
            in2 => \N__40517\,
            in3 => \N__44326\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47123\,
            in2 => \N__46802\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_15\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44138\,
            in2 => \N__43676\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_12_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43952\,
            in2 => \N__43412\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47552\,
            in2 => \N__47690\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40712\,
            in2 => \N__40706\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48995\,
            in2 => \N__49070\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47408\,
            in2 => \N__47345\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_30_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40736\,
            in2 => \N__40727\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40715\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__44449\,
            in1 => \N__40556\,
            in2 => \N__40640\,
            in3 => \N__44430\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011001111"
        )
    port map (
            in0 => \N__40555\,
            in1 => \N__40639\,
            in2 => \N__44432\,
            in3 => \N__44448\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48690\,
            in1 => \N__40670\,
            in2 => \_gnd_net_\,
            in3 => \N__40690\,
            lcout => \elapsed_time_ns_1_RNI36DN9_0_25\,
            ltout => \elapsed_time_ns_1_RNI36DN9_0_25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_25_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__40671\,
            in1 => \_gnd_net_\,
            in2 => \N__40643\,
            in3 => \N__48692\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50245\,
            ce => \N__49799\,
            sr => \N__49433\
        );

    \phase_controller_inst1.stoper_hc.target_time_24_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40626\,
            in1 => \N__40582\,
            in2 => \_gnd_net_\,
            in3 => \N__48691\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50245\,
            ce => \N__49799\,
            sr => \N__49433\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__45790\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50233\,
            ce => \N__44960\,
            sr => \N__49444\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40835\,
            lcout => \current_shift_inst.un4_control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__40836\,
            in1 => \N__45452\,
            in2 => \N__40910\,
            in3 => \N__40810\,
            lcout => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__40837\,
            in1 => \N__40809\,
            in2 => \_gnd_net_\,
            in3 => \N__44865\,
            lcout => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45453\,
            in2 => \_gnd_net_\,
            in3 => \N__43000\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__42952\,
            in1 => \N__45444\,
            in2 => \N__40751\,
            in3 => \N__42880\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45445\,
            in1 => \N__42881\,
            in2 => \N__42953\,
            in3 => \N__40750\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45446\,
            in2 => \_gnd_net_\,
            in3 => \N__42879\,
            lcout => \current_shift_inst.un38_control_input_axb_31_s0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__42948\,
            in1 => \N__44864\,
            in2 => \_gnd_net_\,
            in3 => \N__40746\,
            lcout => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45101\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_1\,
            ltout => \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__45102\,
            in1 => \_gnd_net_\,
            in2 => \N__41183\,
            in3 => \N__44863\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45001\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50222\,
            ce => \N__44958\,
            sr => \N__49452\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44731\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50222\,
            ce => \N__44958\,
            sr => \N__49452\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \N__48150\,
            in1 => \N__45033\,
            in2 => \_gnd_net_\,
            in3 => \N__45076\,
            lcout => \current_shift_inst.un38_control_input_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__41566\,
            in1 => \N__45417\,
            in2 => \N__41614\,
            in3 => \N__42860\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44899\,
            in1 => \N__41134\,
            in2 => \_gnd_net_\,
            in3 => \N__41103\,
            lcout => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__41895\,
            in1 => \N__44903\,
            in2 => \_gnd_net_\,
            in3 => \N__41080\,
            lcout => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__44900\,
            in1 => \_gnd_net_\,
            in2 => \N__41059\,
            in3 => \N__40998\,
            lcout => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__40983\,
            in1 => \N__44902\,
            in2 => \_gnd_net_\,
            in3 => \N__40932\,
            lcout => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44901\,
            in1 => \N__41607\,
            in2 => \_gnd_net_\,
            in3 => \N__41565\,
            lcout => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__45461\,
            in1 => \N__45416\,
            in2 => \_gnd_net_\,
            in3 => \N__45103\,
            lcout => \current_shift_inst.un38_control_input_cry_0_s0_sf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__42075\,
            in1 => \N__44909\,
            in2 => \_gnd_net_\,
            in3 => \N__41535\,
            lcout => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__41513\,
            in1 => \N__45424\,
            in2 => \N__42911\,
            in3 => \N__41479\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI34N61_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__41427\,
            in1 => \N__44911\,
            in2 => \_gnd_net_\,
            in3 => \N__41397\,
            lcout => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44908\,
            in1 => \N__41376\,
            in2 => \_gnd_net_\,
            in3 => \N__41337\,
            lcout => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__45425\,
            in1 => \N__42906\,
            in2 => \N__43001\,
            in3 => \N__45034\,
            lcout => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41301\,
            lcout => \current_shift_inst.un4_control_input_1_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__41250\,
            in1 => \N__44912\,
            in2 => \_gnd_net_\,
            in3 => \N__41199\,
            lcout => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44910\,
            in1 => \N__41958\,
            in2 => \_gnd_net_\,
            in3 => \N__41916\,
            lcout => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43136\,
            lcout => \current_shift_inst.un4_control_input_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41885\,
            lcout => \current_shift_inst.un4_control_input_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__41856\,
            in1 => \N__44914\,
            in2 => \_gnd_net_\,
            in3 => \N__41808\,
            lcout => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44913\,
            in1 => \N__41781\,
            in2 => \_gnd_net_\,
            in3 => \N__41742\,
            lcout => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__41706\,
            in1 => \N__44915\,
            in2 => \_gnd_net_\,
            in3 => \N__41721\,
            lcout => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41705\,
            lcout => \current_shift_inst.un4_control_input_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__41670\,
            in1 => \N__44916\,
            in2 => \_gnd_net_\,
            in3 => \N__41631\,
            lcout => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__43137\,
            in1 => \N__44928\,
            in2 => \_gnd_net_\,
            in3 => \N__43089\,
            lcout => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44907\,
            in1 => \N__43055\,
            in2 => \_gnd_net_\,
            in3 => \N__43033\,
            lcout => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110011"
        )
    port map (
            in0 => \N__42908\,
            in1 => \N__45406\,
            in2 => \N__42996\,
            in3 => \N__45044\,
            lcout => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42934\,
            lcout => \current_shift_inst.un4_control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__42907\,
            in1 => \N__45405\,
            in2 => \N__42287\,
            in3 => \N__42256\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45404\,
            in1 => \N__42198\,
            in2 => \_gnd_net_\,
            in3 => \N__42162\,
            lcout => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__42132\,
            in1 => \N__44905\,
            in2 => \_gnd_net_\,
            in3 => \N__42108\,
            lcout => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42065\,
            lcout => \current_shift_inst.un4_control_input_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__42022\,
            in1 => \N__44906\,
            in2 => \_gnd_net_\,
            in3 => \N__41992\,
            lcout => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_0_c_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45043\,
            in2 => \N__45062\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_20_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48151\,
            in2 => \N__43211\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_0\,
            carryout => \current_shift_inst.un10_control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43196\,
            in2 => \N__48248\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_1\,
            carryout => \current_shift_inst.un10_control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48155\,
            in2 => \N__43190\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_2\,
            carryout => \current_shift_inst.un10_control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43181\,
            in2 => \N__48249\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_3\,
            carryout => \current_shift_inst.un10_control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48159\,
            in2 => \N__43169\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_4\,
            carryout => \current_shift_inst.un10_control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43157\,
            in2 => \N__48250\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_5\,
            carryout => \current_shift_inst.un10_control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48163\,
            in2 => \N__43148\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_6\,
            carryout => \current_shift_inst.un10_control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48263\,
            in2 => \N__43307\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_21_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43292\,
            in2 => \N__48337\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_8\,
            carryout => \current_shift_inst.un10_control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48251\,
            in2 => \N__43283\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_9\,
            carryout => \current_shift_inst.un10_control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44789\,
            in2 => \N__48334\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_10\,
            carryout => \current_shift_inst.un10_control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48255\,
            in2 => \N__43268\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_11\,
            carryout => \current_shift_inst.un10_control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43253\,
            in2 => \N__48335\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_12\,
            carryout => \current_shift_inst.un10_control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_LC_17_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48259\,
            in2 => \N__43244\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_13\,
            carryout => \current_shift_inst.un10_control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_LC_17_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43232\,
            in2 => \N__48336\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_14\,
            carryout => \current_shift_inst.un10_control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_LC_17_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48267\,
            in2 => \N__43223\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_22_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_LC_17_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43397\,
            in2 => \N__48338\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_16\,
            carryout => \current_shift_inst.un10_control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_LC_17_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48271\,
            in2 => \N__43388\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_17\,
            carryout => \current_shift_inst.un10_control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_LC_17_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43373\,
            in2 => \N__48339\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_18\,
            carryout => \current_shift_inst.un10_control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_LC_17_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48275\,
            in2 => \N__43361\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_19\,
            carryout => \current_shift_inst.un10_control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_LC_17_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43346\,
            in2 => \N__48340\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_20\,
            carryout => \current_shift_inst.un10_control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_LC_17_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48279\,
            in2 => \N__43337\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_21\,
            carryout => \current_shift_inst.un10_control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_LC_17_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43325\,
            in2 => \N__48341\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_22\,
            carryout => \current_shift_inst.un10_control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_LC_17_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48283\,
            in2 => \N__43316\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_23_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_LC_17_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43661\,
            in2 => \N__48342\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_24\,
            carryout => \current_shift_inst.un10_control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_LC_17_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48287\,
            in2 => \N__43655\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_25\,
            carryout => \current_shift_inst.un10_control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_LC_17_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43646\,
            in2 => \N__48343\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_26\,
            carryout => \current_shift_inst.un10_control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_LC_17_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48291\,
            in2 => \N__43640\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_27\,
            carryout => \current_shift_inst.un10_control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_LC_17_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43622\,
            in2 => \N__48344\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_28\,
            carryout => \current_shift_inst.un10_control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_LC_17_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48295\,
            in2 => \N__43610\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_29\,
            carryout => \current_shift_inst.un10_control_input_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_17_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45450\,
            in2 => \_gnd_net_\,
            in3 => \N__43595\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_20_LC_18_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43881\,
            in1 => \N__43940\,
            in2 => \_gnd_net_\,
            in3 => \N__48829\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50320\,
            ce => \N__49807\,
            sr => \N__49393\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_18_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110101000100"
        )
    port map (
            in0 => \N__44479\,
            in1 => \N__43964\,
            in2 => \N__44507\,
            in3 => \N__43973\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_18_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011001111"
        )
    port map (
            in0 => \N__43972\,
            in1 => \N__43963\,
            in2 => \N__44483\,
            in3 => \N__44506\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_18_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43885\,
            in1 => \N__43939\,
            in2 => \_gnd_net_\,
            in3 => \N__48826\,
            lcout => \elapsed_time_ns_1_RNIU0DN9_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_18_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43865\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50312\,
            ce => \N__43793\,
            sr => \N__49397\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43837\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50312\,
            ce => \N__43793\,
            sr => \N__49397\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_18_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43744\,
            in1 => \N__46409\,
            in2 => \_gnd_net_\,
            in3 => \N__48651\,
            lcout => \elapsed_time_ns_1_RNIE03T9_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_18_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48652\,
            in1 => \N__43720\,
            in2 => \_gnd_net_\,
            in3 => \N__46459\,
            lcout => \elapsed_time_ns_1_RNIF13T9_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_18_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43696\,
            in1 => \N__46383\,
            in2 => \_gnd_net_\,
            in3 => \N__48653\,
            lcout => \elapsed_time_ns_1_RNIG23T9_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110101000100"
        )
    port map (
            in0 => \N__44528\,
            in1 => \N__44071\,
            in2 => \N__44552\,
            in3 => \N__44003\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__44002\,
            in1 => \N__44527\,
            in2 => \N__44072\,
            in3 => \N__44548\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44103\,
            in1 => \N__48668\,
            in2 => \_gnd_net_\,
            in3 => \N__44119\,
            lcout => \elapsed_time_ns_1_RNI68CN9_0_19\,
            ltout => \elapsed_time_ns_1_RNI68CN9_0_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_19_LC_18_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__48670\,
            in1 => \_gnd_net_\,
            in2 => \N__44108\,
            in3 => \N__44104\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50302\,
            ce => \N__49835\,
            sr => \N__49401\
        );

    \phase_controller_inst1.stoper_hc.target_time_15_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44060\,
            in1 => \N__44039\,
            in2 => \_gnd_net_\,
            in3 => \N__48671\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50302\,
            ce => \N__49835\,
            sr => \N__49401\
        );

    \phase_controller_inst1.stoper_hc.target_time_18_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48669\,
            in1 => \N__47945\,
            in2 => \_gnd_net_\,
            in3 => \N__47924\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50302\,
            ce => \N__49835\,
            sr => \N__49401\
        );

    \phase_controller_inst1.stoper_hc.running_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111001100"
        )
    port map (
            in0 => \N__46835\,
            in1 => \N__47002\,
            in2 => \N__46957\,
            in3 => \N__46987\,
            lcout => \phase_controller_inst1.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50291\,
            ce => 'H',
            sr => \N__49404\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNID63H_30_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46834\,
            in2 => \_gnd_net_\,
            in3 => \N__46950\,
            lcout => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43994\,
            in3 => \N__46985\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1_30_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46986\,
            in2 => \_gnd_net_\,
            in3 => \N__43984\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1Z0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44306\,
            in2 => \N__44300\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_11_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49744\,
            in1 => \N__44267\,
            in2 => \_gnd_net_\,
            in3 => \N__44255\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \N__50279\,
            ce => 'H',
            sr => \N__49410\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__49788\,
            in1 => \N__44243\,
            in2 => \N__44252\,
            in3 => \N__44231\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \N__50279\,
            ce => 'H',
            sr => \N__49410\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49745\,
            in1 => \N__44228\,
            in2 => \_gnd_net_\,
            in3 => \N__44216\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \N__50279\,
            ce => 'H',
            sr => \N__49410\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49789\,
            in1 => \N__44213\,
            in2 => \_gnd_net_\,
            in3 => \N__44201\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \N__50279\,
            ce => 'H',
            sr => \N__49410\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49746\,
            in1 => \N__44198\,
            in2 => \_gnd_net_\,
            in3 => \N__44186\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \N__50279\,
            ce => 'H',
            sr => \N__49410\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49790\,
            in1 => \N__44183\,
            in2 => \_gnd_net_\,
            in3 => \N__44171\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \N__50279\,
            ce => 'H',
            sr => \N__49410\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49747\,
            in1 => \N__44168\,
            in2 => \_gnd_net_\,
            in3 => \N__44156\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \N__50279\,
            ce => 'H',
            sr => \N__49410\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49850\,
            in1 => \N__44153\,
            in2 => \_gnd_net_\,
            in3 => \N__44141\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_18_12_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \N__50266\,
            ce => 'H',
            sr => \N__49415\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49774\,
            in1 => \N__44408\,
            in2 => \_gnd_net_\,
            in3 => \N__44396\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \N__50266\,
            ce => 'H',
            sr => \N__49415\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49847\,
            in1 => \N__44393\,
            in2 => \_gnd_net_\,
            in3 => \N__44381\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \N__50266\,
            ce => 'H',
            sr => \N__49415\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49775\,
            in1 => \N__44374\,
            in2 => \_gnd_net_\,
            in3 => \N__44360\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \N__50266\,
            ce => 'H',
            sr => \N__49415\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49848\,
            in1 => \N__44357\,
            in2 => \_gnd_net_\,
            in3 => \N__44345\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \N__50266\,
            ce => 'H',
            sr => \N__49415\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49776\,
            in1 => \N__44342\,
            in2 => \_gnd_net_\,
            in3 => \N__44330\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \N__50266\,
            ce => 'H',
            sr => \N__49415\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49849\,
            in1 => \N__44327\,
            in2 => \_gnd_net_\,
            in3 => \N__44315\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \N__50266\,
            ce => 'H',
            sr => \N__49415\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_18_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49777\,
            in1 => \N__47180\,
            in2 => \_gnd_net_\,
            in3 => \N__44312\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \N__50266\,
            ce => 'H',
            sr => \N__49415\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49766\,
            in1 => \N__47149\,
            in2 => \_gnd_net_\,
            in3 => \N__44309\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_18_13_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \N__50257\,
            ce => 'H',
            sr => \N__49424\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49836\,
            in1 => \N__44547\,
            in2 => \_gnd_net_\,
            in3 => \N__44531\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \N__50257\,
            ce => 'H',
            sr => \N__49424\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49767\,
            in1 => \N__44526\,
            in2 => \_gnd_net_\,
            in3 => \N__44510\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \N__50257\,
            ce => 'H',
            sr => \N__49424\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49837\,
            in1 => \N__44502\,
            in2 => \_gnd_net_\,
            in3 => \N__44486\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \N__50257\,
            ce => 'H',
            sr => \N__49424\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49768\,
            in1 => \N__44478\,
            in2 => \_gnd_net_\,
            in3 => \N__44459\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\,
            clk => \N__50257\,
            ce => 'H',
            sr => \N__49424\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49838\,
            in1 => \N__47575\,
            in2 => \_gnd_net_\,
            in3 => \N__44456\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\,
            clk => \N__50257\,
            ce => 'H',
            sr => \N__49424\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49769\,
            in1 => \N__47602\,
            in2 => \_gnd_net_\,
            in3 => \N__44453\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\,
            clk => \N__50257\,
            ce => 'H',
            sr => \N__49424\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49839\,
            in1 => \N__44450\,
            in2 => \_gnd_net_\,
            in3 => \N__44435\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\,
            clk => \N__50257\,
            ce => 'H',
            sr => \N__49424\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49770\,
            in1 => \N__44431\,
            in2 => \_gnd_net_\,
            in3 => \N__44414\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_18_14_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\,
            clk => \N__50246\,
            ce => 'H',
            sr => \N__49434\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49851\,
            in1 => \N__49020\,
            in2 => \_gnd_net_\,
            in3 => \N__44411\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\,
            clk => \N__50246\,
            ce => 'H',
            sr => \N__49434\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49771\,
            in1 => \N__49044\,
            in2 => \_gnd_net_\,
            in3 => \N__44702\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\,
            clk => \N__50246\,
            ce => 'H',
            sr => \N__49434\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49852\,
            in1 => \N__47373\,
            in2 => \_gnd_net_\,
            in3 => \N__44699\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\,
            clk => \N__50246\,
            ce => 'H',
            sr => \N__49434\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49772\,
            in1 => \N__47394\,
            in2 => \_gnd_net_\,
            in3 => \N__44696\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\,
            clk => \N__50246\,
            ce => 'H',
            sr => \N__49434\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49853\,
            in1 => \N__44680\,
            in2 => \_gnd_net_\,
            in3 => \N__44666\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\,
            clk => \N__50246\,
            ce => 'H',
            sr => \N__49434\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49773\,
            in1 => \N__44653\,
            in2 => \_gnd_net_\,
            in3 => \N__44663\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50246\,
            ce => 'H',
            sr => \N__49434\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110101000100"
        )
    port map (
            in0 => \N__44596\,
            in1 => \N__47249\,
            in2 => \N__44624\,
            in3 => \N__47261\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__47260\,
            in1 => \N__44623\,
            in2 => \N__44600\,
            in3 => \N__47248\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_28_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48839\,
            in1 => \N__47305\,
            in2 => \_gnd_net_\,
            in3 => \N__47330\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50234\,
            ce => \N__47865\,
            sr => \N__49445\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101000101"
        )
    port map (
            in0 => \N__45511\,
            in1 => \N__45544\,
            in2 => \N__45536\,
            in3 => \N__47032\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011110010"
        )
    port map (
            in0 => \N__45545\,
            in1 => \N__45532\,
            in2 => \N__47036\,
            in3 => \N__45512\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__45481\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input1_1\,
            ltout => \current_shift_inst.un4_control_input1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45418\,
            in2 => \N__45107\,
            in3 => \N__45104\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_0_c_inv_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \N__48333\,
            in1 => \N__44966\,
            in2 => \_gnd_net_\,
            in3 => \N__45058\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45002\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_fast_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50223\,
            ce => \N__44959\,
            sr => \N__49453\
        );

    \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__44775\,
            in1 => \N__44904\,
            in2 => \_gnd_net_\,
            in3 => \N__44811\,
            lcout => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_18_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44774\,
            lcout => \current_shift_inst.un4_control_input_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.counter_0_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46693\,
            in1 => \N__44724\,
            in2 => \_gnd_net_\,
            in3 => \N__44705\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_18_17_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_0\,
            clk => \N__50211\,
            ce => \N__46551\,
            sr => \N__49459\
        );

    \current_shift_inst.timer_s1.counter_1_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46697\,
            in1 => \N__45783\,
            in2 => \_gnd_net_\,
            in3 => \N__45764\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_0\,
            carryout => \current_shift_inst.timer_s1.counter_cry_1\,
            clk => \N__50211\,
            ce => \N__46551\,
            sr => \N__49459\
        );

    \current_shift_inst.timer_s1.counter_2_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46694\,
            in1 => \N__45753\,
            in2 => \_gnd_net_\,
            in3 => \N__45734\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_1\,
            carryout => \current_shift_inst.timer_s1.counter_cry_2\,
            clk => \N__50211\,
            ce => \N__46551\,
            sr => \N__49459\
        );

    \current_shift_inst.timer_s1.counter_3_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46698\,
            in1 => \N__45718\,
            in2 => \_gnd_net_\,
            in3 => \N__45704\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_2\,
            carryout => \current_shift_inst.timer_s1.counter_cry_3\,
            clk => \N__50211\,
            ce => \N__46551\,
            sr => \N__49459\
        );

    \current_shift_inst.timer_s1.counter_4_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46695\,
            in1 => \N__45690\,
            in2 => \_gnd_net_\,
            in3 => \N__45674\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_3\,
            carryout => \current_shift_inst.timer_s1.counter_cry_4\,
            clk => \N__50211\,
            ce => \N__46551\,
            sr => \N__49459\
        );

    \current_shift_inst.timer_s1.counter_5_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46699\,
            in1 => \N__45660\,
            in2 => \_gnd_net_\,
            in3 => \N__45644\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_4\,
            carryout => \current_shift_inst.timer_s1.counter_cry_5\,
            clk => \N__50211\,
            ce => \N__46551\,
            sr => \N__49459\
        );

    \current_shift_inst.timer_s1.counter_6_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46696\,
            in1 => \N__45630\,
            in2 => \_gnd_net_\,
            in3 => \N__45614\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_5\,
            carryout => \current_shift_inst.timer_s1.counter_cry_6\,
            clk => \N__50211\,
            ce => \N__46551\,
            sr => \N__49459\
        );

    \current_shift_inst.timer_s1.counter_7_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46700\,
            in1 => \N__45600\,
            in2 => \_gnd_net_\,
            in3 => \N__45584\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_6\,
            carryout => \current_shift_inst.timer_s1.counter_cry_7\,
            clk => \N__50211\,
            ce => \N__46551\,
            sr => \N__49459\
        );

    \current_shift_inst.timer_s1.counter_8_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46664\,
            in1 => \N__45570\,
            in2 => \_gnd_net_\,
            in3 => \N__45548\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_18_18_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_8\,
            clk => \N__50201\,
            ce => \N__46552\,
            sr => \N__49467\
        );

    \current_shift_inst.timer_s1.counter_9_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46674\,
            in1 => \N__46050\,
            in2 => \_gnd_net_\,
            in3 => \N__46028\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_8\,
            carryout => \current_shift_inst.timer_s1.counter_cry_9\,
            clk => \N__50201\,
            ce => \N__46552\,
            sr => \N__49467\
        );

    \current_shift_inst.timer_s1.counter_10_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46661\,
            in1 => \N__46023\,
            in2 => \_gnd_net_\,
            in3 => \N__46004\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_9\,
            carryout => \current_shift_inst.timer_s1.counter_cry_10\,
            clk => \N__50201\,
            ce => \N__46552\,
            sr => \N__49467\
        );

    \current_shift_inst.timer_s1.counter_11_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46671\,
            in1 => \N__45994\,
            in2 => \_gnd_net_\,
            in3 => \N__45980\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_10\,
            carryout => \current_shift_inst.timer_s1.counter_cry_11\,
            clk => \N__50201\,
            ce => \N__46552\,
            sr => \N__49467\
        );

    \current_shift_inst.timer_s1.counter_12_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46662\,
            in1 => \N__45964\,
            in2 => \_gnd_net_\,
            in3 => \N__45950\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_11\,
            carryout => \current_shift_inst.timer_s1.counter_cry_12\,
            clk => \N__50201\,
            ce => \N__46552\,
            sr => \N__49467\
        );

    \current_shift_inst.timer_s1.counter_13_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46672\,
            in1 => \N__45934\,
            in2 => \_gnd_net_\,
            in3 => \N__45920\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_12\,
            carryout => \current_shift_inst.timer_s1.counter_cry_13\,
            clk => \N__50201\,
            ce => \N__46552\,
            sr => \N__49467\
        );

    \current_shift_inst.timer_s1.counter_14_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46663\,
            in1 => \N__45910\,
            in2 => \_gnd_net_\,
            in3 => \N__45896\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_13\,
            carryout => \current_shift_inst.timer_s1.counter_cry_14\,
            clk => \N__50201\,
            ce => \N__46552\,
            sr => \N__49467\
        );

    \current_shift_inst.timer_s1.counter_15_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46673\,
            in1 => \N__45882\,
            in2 => \_gnd_net_\,
            in3 => \N__45866\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_14\,
            carryout => \current_shift_inst.timer_s1.counter_cry_15\,
            clk => \N__50201\,
            ce => \N__46552\,
            sr => \N__49467\
        );

    \current_shift_inst.timer_s1.counter_16_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46657\,
            in1 => \N__45849\,
            in2 => \_gnd_net_\,
            in3 => \N__45827\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_18_19_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_16\,
            clk => \N__50194\,
            ce => \N__46553\,
            sr => \N__49474\
        );

    \current_shift_inst.timer_s1.counter_17_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46665\,
            in1 => \N__45813\,
            in2 => \_gnd_net_\,
            in3 => \N__46304\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_16\,
            carryout => \current_shift_inst.timer_s1.counter_cry_17\,
            clk => \N__50194\,
            ce => \N__46553\,
            sr => \N__49474\
        );

    \current_shift_inst.timer_s1.counter_18_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46658\,
            in1 => \N__46296\,
            in2 => \_gnd_net_\,
            in3 => \N__46274\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_17\,
            carryout => \current_shift_inst.timer_s1.counter_cry_18\,
            clk => \N__50194\,
            ce => \N__46553\,
            sr => \N__49474\
        );

    \current_shift_inst.timer_s1.counter_19_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46666\,
            in1 => \N__46264\,
            in2 => \_gnd_net_\,
            in3 => \N__46250\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_18\,
            carryout => \current_shift_inst.timer_s1.counter_cry_19\,
            clk => \N__50194\,
            ce => \N__46553\,
            sr => \N__49474\
        );

    \current_shift_inst.timer_s1.counter_20_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46659\,
            in1 => \N__46236\,
            in2 => \_gnd_net_\,
            in3 => \N__46220\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_19\,
            carryout => \current_shift_inst.timer_s1.counter_cry_20\,
            clk => \N__50194\,
            ce => \N__46553\,
            sr => \N__49474\
        );

    \current_shift_inst.timer_s1.counter_21_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46667\,
            in1 => \N__46204\,
            in2 => \_gnd_net_\,
            in3 => \N__46190\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_20\,
            carryout => \current_shift_inst.timer_s1.counter_cry_21\,
            clk => \N__50194\,
            ce => \N__46553\,
            sr => \N__49474\
        );

    \current_shift_inst.timer_s1.counter_22_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46660\,
            in1 => \N__46180\,
            in2 => \_gnd_net_\,
            in3 => \N__46166\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_21\,
            carryout => \current_shift_inst.timer_s1.counter_cry_22\,
            clk => \N__50194\,
            ce => \N__46553\,
            sr => \N__49474\
        );

    \current_shift_inst.timer_s1.counter_23_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46668\,
            in1 => \N__46156\,
            in2 => \_gnd_net_\,
            in3 => \N__46142\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_22\,
            carryout => \current_shift_inst.timer_s1.counter_cry_23\,
            clk => \N__50194\,
            ce => \N__46553\,
            sr => \N__49474\
        );

    \current_shift_inst.timer_s1.counter_24_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46653\,
            in1 => \N__46125\,
            in2 => \_gnd_net_\,
            in3 => \N__46103\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_18_20_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_24\,
            clk => \N__50188\,
            ce => \N__46544\,
            sr => \N__49481\
        );

    \current_shift_inst.timer_s1.counter_25_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46669\,
            in1 => \N__46086\,
            in2 => \_gnd_net_\,
            in3 => \N__46064\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_24\,
            carryout => \current_shift_inst.timer_s1.counter_cry_25\,
            clk => \N__50188\,
            ce => \N__46544\,
            sr => \N__49481\
        );

    \current_shift_inst.timer_s1.counter_26_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46654\,
            in1 => \N__46776\,
            in2 => \_gnd_net_\,
            in3 => \N__46754\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_25\,
            carryout => \current_shift_inst.timer_s1.counter_cry_26\,
            clk => \N__50188\,
            ce => \N__46544\,
            sr => \N__49481\
        );

    \current_shift_inst.timer_s1.counter_27_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46670\,
            in1 => \N__46740\,
            in2 => \_gnd_net_\,
            in3 => \N__46724\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_26\,
            carryout => \current_shift_inst.timer_s1.counter_cry_27\,
            clk => \N__50188\,
            ce => \N__46544\,
            sr => \N__49481\
        );

    \current_shift_inst.timer_s1.counter_28_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46655\,
            in1 => \N__46717\,
            in2 => \_gnd_net_\,
            in3 => \N__46703\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_27\,
            carryout => \current_shift_inst.timer_s1.counter_cry_28\,
            clk => \N__50188\,
            ce => \N__46544\,
            sr => \N__49481\
        );

    \current_shift_inst.timer_s1.counter_29_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__46567\,
            in1 => \N__46656\,
            in2 => \_gnd_net_\,
            in3 => \N__46574\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50188\,
            ce => \N__46544\,
            sr => \N__49481\
        );

    \phase_controller_inst1.T12_LC_18_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46498\,
            in2 => \_gnd_net_\,
            in3 => \N__48063\,
            lcout => \T12_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50183\,
            ce => 'H',
            sr => \N__49492\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_20_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__46476\,
            in1 => \N__46339\,
            in2 => \_gnd_net_\,
            in3 => \N__48835\,
            lcout => \elapsed_time_ns_1_RNIDV2T9_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_20_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__46458\,
            in1 => \N__46414\,
            in2 => \N__46385\,
            in3 => \N__46331\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_20_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47944\,
            in1 => \N__47923\,
            in2 => \_gnd_net_\,
            in3 => \N__48759\,
            lcout => \elapsed_time_ns_1_RNI57CN9_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_20_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__47301\,
            in1 => \N__48968\,
            in2 => \_gnd_net_\,
            in3 => \N__47018\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_20_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47748\,
            in1 => \N__47728\,
            in2 => \_gnd_net_\,
            in3 => \N__48757\,
            lcout => \elapsed_time_ns_1_RNI03DN9_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_20_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48758\,
            in1 => \N__47475\,
            in2 => \_gnd_net_\,
            in3 => \N__47447\,
            lcout => \elapsed_time_ns_1_RNI7ADN9_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_20_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__46821\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46851\,
            lcout => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_20_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48859\,
            in1 => \N__50385\,
            in2 => \_gnd_net_\,
            in3 => \N__50355\,
            lcout => \elapsed_time_ns_1_RNI47DN9_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_20_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__46820\,
            in1 => \N__47003\,
            in2 => \_gnd_net_\,
            in3 => \N__46850\,
            lcout => \phase_controller_inst1.stoper_hc.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_LC_20_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010001011100010"
        )
    port map (
            in0 => \N__47996\,
            in1 => \N__46981\,
            in2 => \N__46833\,
            in3 => \N__46958\,
            lcout => \phase_controller_inst1.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50303\,
            ce => 'H',
            sr => \N__49411\
        );

    \phase_controller_inst1.start_timer_hc_LC_20_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__46930\,
            in1 => \N__47962\,
            in2 => \N__46856\,
            in3 => \N__46871\,
            lcout => \phase_controller_inst1.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50303\,
            ce => 'H',
            sr => \N__49411\
        );

    \phase_controller_inst1.stoper_hc.start_latched_LC_20_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46852\,
            lcout => \phase_controller_inst1.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50303\,
            ce => 'H',
            sr => \N__49411\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_20_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100000010"
        )
    port map (
            in0 => \N__47765\,
            in1 => \N__47178\,
            in2 => \N__47161\,
            in3 => \N__47132\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_20_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47825\,
            in1 => \N__47802\,
            in2 => \_gnd_net_\,
            in3 => \N__48862\,
            lcout => \elapsed_time_ns_1_RNI35CN9_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_20_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48861\,
            in1 => \N__47215\,
            in2 => \_gnd_net_\,
            in3 => \N__47227\,
            lcout => \elapsed_time_ns_1_RNI46CN9_0_17\,
            ltout => \elapsed_time_ns_1_RNI46CN9_0_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_17_LC_20_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__47216\,
            in1 => \_gnd_net_\,
            in2 => \N__47183\,
            in3 => \N__48863\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50292\,
            ce => \N__49735\,
            sr => \N__49416\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_20_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__47764\,
            in1 => \N__47179\,
            in2 => \N__47162\,
            in3 => \N__47131\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_20_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__47107\,
            in1 => \N__48860\,
            in2 => \_gnd_net_\,
            in3 => \N__47092\,
            lcout => \elapsed_time_ns_1_RNI13CN9_0_14\,
            ltout => \elapsed_time_ns_1_RNI13CN9_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_14_LC_20_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__47093\,
            in1 => \_gnd_net_\,
            in2 => \N__47063\,
            in3 => \N__48925\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50292\,
            ce => \N__49735\,
            sr => \N__49416\
        );

    \phase_controller_inst2.stoper_hc.target_time_16_LC_20_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47823\,
            in1 => \N__47803\,
            in2 => \_gnd_net_\,
            in3 => \N__48870\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50280\,
            ce => \N__47870\,
            sr => \N__49425\
        );

    \phase_controller_inst2.stoper_hc.target_time_29_LC_20_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48869\,
            in1 => \N__47476\,
            in2 => \_gnd_net_\,
            in3 => \N__47456\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50280\,
            ce => \N__47870\,
            sr => \N__49425\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_20_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48830\,
            in1 => \N__47521\,
            in2 => \_gnd_net_\,
            in3 => \N__47533\,
            lcout => \elapsed_time_ns_1_RNIJ53T9_0_7\,
            ltout => \elapsed_time_ns_1_RNIJ53T9_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_LC_20_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__47522\,
            in1 => \_gnd_net_\,
            in2 => \N__47492\,
            in3 => \N__48834\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50268\,
            ce => \N__49734\,
            sr => \N__49435\
        );

    \phase_controller_inst1.stoper_hc.target_time_29_LC_20_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47477\,
            in1 => \N__47455\,
            in2 => \_gnd_net_\,
            in3 => \N__48833\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50268\,
            ce => \N__49734\,
            sr => \N__49435\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_20_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__47269\,
            in1 => \N__47395\,
            in2 => \N__47378\,
            in3 => \N__47353\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_20_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__47396\,
            in1 => \N__47374\,
            in2 => \N__47357\,
            in3 => \N__47270\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_20_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48831\,
            in1 => \N__47311\,
            in2 => \_gnd_net_\,
            in3 => \N__47323\,
            lcout => \elapsed_time_ns_1_RNI69DN9_0_28\,
            ltout => \elapsed_time_ns_1_RNI69DN9_0_28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_28_LC_20_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__47312\,
            in1 => \_gnd_net_\,
            in2 => \N__47273\,
            in3 => \N__48832\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50268\,
            ce => \N__49734\,
            sr => \N__49435\
        );

    \phase_controller_inst2.stoper_hc.target_time_26_LC_20_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__50390\,
            in1 => \N__50366\,
            in2 => \_gnd_net_\,
            in3 => \N__48924\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50258\,
            ce => \N__47868\,
            sr => \N__49446\
        );

    \phase_controller_inst2.stoper_hc.target_time_27_LC_20_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48923\,
            in1 => \N__48983\,
            in2 => \_gnd_net_\,
            in3 => \N__48467\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50258\,
            ce => \N__47868\,
            sr => \N__49446\
        );

    \phase_controller_inst1.state_RNIE87F_2_LC_20_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48064\,
            in2 => \_gnd_net_\,
            in3 => \N__48000\,
            lcout => \phase_controller_inst1.state_RNIE87FZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_18_LC_21_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47943\,
            in1 => \N__47922\,
            in2 => \_gnd_net_\,
            in3 => \N__48873\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50318\,
            ce => \N__47873\,
            sr => \N__49412\
        );

    \phase_controller_inst1.stoper_hc.target_time_16_LC_21_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47824\,
            in1 => \N__47807\,
            in2 => \_gnd_net_\,
            in3 => \N__48874\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50313\,
            ce => \N__49803\,
            sr => \N__49417\
        );

    \phase_controller_inst1.stoper_hc.target_time_22_LC_21_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47749\,
            in1 => \N__47729\,
            in2 => \_gnd_net_\,
            in3 => \N__48875\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50313\,
            ce => \N__49803\,
            sr => \N__49417\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_21_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__47618\,
            in1 => \N__47609\,
            in2 => \N__47588\,
            in3 => \N__47561\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_21_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48857\,
            in1 => \N__47656\,
            in2 => \_gnd_net_\,
            in3 => \N__47668\,
            lcout => \elapsed_time_ns_1_RNI14DN9_0_23\,
            ltout => \elapsed_time_ns_1_RNI14DN9_0_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_23_LC_21_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__47657\,
            in1 => \_gnd_net_\,
            in2 => \N__47621\,
            in3 => \N__48858\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50304\,
            ce => \N__49733\,
            sr => \N__49426\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_21_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__47617\,
            in1 => \N__47608\,
            in2 => \N__47587\,
            in3 => \N__47560\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_27_LC_21_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48871\,
            in1 => \N__48978\,
            in2 => \_gnd_net_\,
            in3 => \N__48463\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50293\,
            ce => \N__49804\,
            sr => \N__49436\
        );

    \phase_controller_inst1.stoper_hc.target_time_26_LC_21_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__50386\,
            in1 => \N__50362\,
            in2 => \_gnd_net_\,
            in3 => \N__48872\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50293\,
            ce => \N__49804\,
            sr => \N__49436\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_21_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__49055\,
            in1 => \N__49046\,
            in2 => \N__49028\,
            in3 => \N__49004\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_21_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__49054\,
            in1 => \N__49045\,
            in2 => \N__49027\,
            in3 => \N__49003\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_22_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__48462\,
            in1 => \N__48982\,
            in2 => \_gnd_net_\,
            in3 => \N__48909\,
            lcout => \elapsed_time_ns_1_RNI58DN9_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_24_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
