-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Oct 16 2025 00:42:38

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MAIN" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MAIN
entity MAIN is
port (
    s3_phy : out std_logic;
    il_min_comp2 : in std_logic;
    il_max_comp1 : in std_logic;
    s1_phy : out std_logic;
    reset : in std_logic;
    il_min_comp1 : in std_logic;
    delay_tr_input : in std_logic;
    s4_phy : out std_logic;
    rgb_g : out std_logic;
    start_stop : in std_logic;
    s2_phy : out std_logic;
    rgb_r : out std_logic;
    rgb_b : out std_logic;
    pwm_output : out std_logic;
    il_max_comp2 : in std_logic;
    delay_hc_input : in std_logic);
end MAIN;

-- Architecture of MAIN
-- View name is \INTERFACE\
architecture \INTERFACE\ of MAIN is

signal \N__21137\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21124\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21081\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21052\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21027\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21025\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21004\ : std_logic;
signal \N__21003\ : std_logic;
signal \N__21000\ : std_logic;
signal \N__20997\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20982\ : std_logic;
signal \N__20979\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20973\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20965\ : std_logic;
signal \N__20964\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20955\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20941\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20938\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20926\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20923\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20919\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20916\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20908\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20905\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20902\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20899\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20896\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20887\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20884\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20881\ : std_logic;
signal \N__20880\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20878\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20875\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20871\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20613\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20592\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20589\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20529\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20526\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20523\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20511\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20466\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20463\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20421\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20400\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20397\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20383\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20376\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20373\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20368\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20353\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20347\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20172\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20070\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20010\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19986\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19968\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19911\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19893\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19825\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19795\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19735\ : std_logic;
signal \N__19734\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19725\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19707\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19683\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19662\ : std_logic;
signal \N__19659\ : std_logic;
signal \N__19656\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19639\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19633\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19570\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19560\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19557\ : std_logic;
signal \N__19554\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19546\ : std_logic;
signal \N__19543\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19524\ : std_logic;
signal \N__19521\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19449\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19428\ : std_logic;
signal \N__19425\ : std_logic;
signal \N__19422\ : std_logic;
signal \N__19419\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19405\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19374\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19368\ : std_logic;
signal \N__19365\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19347\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19326\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19320\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19309\ : std_logic;
signal \N__19308\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19299\ : std_logic;
signal \N__19296\ : std_logic;
signal \N__19293\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19276\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19269\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19231\ : std_logic;
signal \N__19230\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19188\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19170\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19131\ : std_logic;
signal \N__19128\ : std_logic;
signal \N__19125\ : std_logic;
signal \N__19122\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19104\ : std_logic;
signal \N__19101\ : std_logic;
signal \N__19098\ : std_logic;
signal \N__19095\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19062\ : std_logic;
signal \N__19059\ : std_logic;
signal \N__19056\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19045\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19028\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19023\ : std_logic;
signal \N__19020\ : std_logic;
signal \N__19017\ : std_logic;
signal \N__19014\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__19003\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18985\ : std_logic;
signal \N__18984\ : std_logic;
signal \N__18981\ : std_logic;
signal \N__18978\ : std_logic;
signal \N__18975\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18949\ : std_logic;
signal \N__18946\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18936\ : std_logic;
signal \N__18933\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18916\ : std_logic;
signal \N__18915\ : std_logic;
signal \N__18912\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18885\ : std_logic;
signal \N__18882\ : std_logic;
signal \N__18877\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18868\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18864\ : std_logic;
signal \N__18859\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18852\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18846\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18840\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18838\ : std_logic;
signal \N__18837\ : std_logic;
signal \N__18834\ : std_logic;
signal \N__18831\ : std_logic;
signal \N__18828\ : std_logic;
signal \N__18825\ : std_logic;
signal \N__18820\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18799\ : std_logic;
signal \N__18796\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18775\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18742\ : std_logic;
signal \N__18741\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18728\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18722\ : std_logic;
signal \N__18721\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18714\ : std_logic;
signal \N__18711\ : std_logic;
signal \N__18708\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18699\ : std_logic;
signal \N__18696\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18687\ : std_logic;
signal \N__18684\ : std_logic;
signal \N__18683\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18680\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18648\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18616\ : std_logic;
signal \N__18613\ : std_logic;
signal \N__18612\ : std_logic;
signal \N__18609\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18600\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18591\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18583\ : std_logic;
signal \N__18580\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18577\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18558\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18546\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18540\ : std_logic;
signal \N__18537\ : std_logic;
signal \N__18534\ : std_logic;
signal \N__18531\ : std_logic;
signal \N__18528\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18520\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18514\ : std_logic;
signal \N__18511\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18505\ : std_logic;
signal \N__18502\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18498\ : std_logic;
signal \N__18495\ : std_logic;
signal \N__18492\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18483\ : std_logic;
signal \N__18480\ : std_logic;
signal \N__18477\ : std_logic;
signal \N__18474\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18462\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18442\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18438\ : std_logic;
signal \N__18435\ : std_logic;
signal \N__18432\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18415\ : std_logic;
signal \N__18412\ : std_logic;
signal \N__18409\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18397\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18390\ : std_logic;
signal \N__18387\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18373\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18367\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18354\ : std_logic;
signal \N__18351\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18345\ : std_logic;
signal \N__18340\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18330\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18321\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18315\ : std_logic;
signal \N__18312\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18304\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18295\ : std_logic;
signal \N__18294\ : std_logic;
signal \N__18291\ : std_logic;
signal \N__18286\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18277\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18271\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18265\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18259\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18250\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18246\ : std_logic;
signal \N__18241\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18235\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18229\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18214\ : std_logic;
signal \N__18211\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18196\ : std_logic;
signal \N__18195\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18164\ : std_logic;
signal \N__18161\ : std_logic;
signal \N__18158\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18151\ : std_logic;
signal \N__18150\ : std_logic;
signal \N__18149\ : std_logic;
signal \N__18148\ : std_logic;
signal \N__18147\ : std_logic;
signal \N__18136\ : std_logic;
signal \N__18133\ : std_logic;
signal \N__18128\ : std_logic;
signal \N__18127\ : std_logic;
signal \N__18126\ : std_logic;
signal \N__18123\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18112\ : std_logic;
signal \N__18107\ : std_logic;
signal \N__18106\ : std_logic;
signal \N__18105\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18099\ : std_logic;
signal \N__18096\ : std_logic;
signal \N__18093\ : std_logic;
signal \N__18090\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18086\ : std_logic;
signal \N__18081\ : std_logic;
signal \N__18078\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18069\ : std_logic;
signal \N__18066\ : std_logic;
signal \N__18059\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18043\ : std_logic;
signal \N__18040\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18030\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18022\ : std_logic;
signal \N__18019\ : std_logic;
signal \N__18018\ : std_logic;
signal \N__18015\ : std_logic;
signal \N__18012\ : std_logic;
signal \N__18009\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__18005\ : std_logic;
signal \N__18002\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17984\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17977\ : std_logic;
signal \N__17974\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17970\ : std_logic;
signal \N__17967\ : std_logic;
signal \N__17964\ : std_logic;
signal \N__17961\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17957\ : std_logic;
signal \N__17952\ : std_logic;
signal \N__17949\ : std_logic;
signal \N__17942\ : std_logic;
signal \N__17941\ : std_logic;
signal \N__17940\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17937\ : std_logic;
signal \N__17932\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17922\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17913\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17902\ : std_logic;
signal \N__17901\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17899\ : std_logic;
signal \N__17896\ : std_logic;
signal \N__17893\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17878\ : std_logic;
signal \N__17875\ : std_logic;
signal \N__17872\ : std_logic;
signal \N__17871\ : std_logic;
signal \N__17866\ : std_logic;
signal \N__17863\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17852\ : std_logic;
signal \N__17851\ : std_logic;
signal \N__17850\ : std_logic;
signal \N__17849\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17843\ : std_logic;
signal \N__17840\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17820\ : std_logic;
signal \N__17817\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17809\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17788\ : std_logic;
signal \N__17787\ : std_logic;
signal \N__17784\ : std_logic;
signal \N__17779\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17770\ : std_logic;
signal \N__17769\ : std_logic;
signal \N__17766\ : std_logic;
signal \N__17763\ : std_logic;
signal \N__17760\ : std_logic;
signal \N__17757\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17745\ : std_logic;
signal \N__17742\ : std_logic;
signal \N__17739\ : std_logic;
signal \N__17736\ : std_logic;
signal \N__17729\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17707\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17701\ : std_logic;
signal \N__17696\ : std_logic;
signal \N__17695\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17689\ : std_logic;
signal \N__17686\ : std_logic;
signal \N__17683\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17671\ : std_logic;
signal \N__17668\ : std_logic;
signal \N__17665\ : std_logic;
signal \N__17662\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17644\ : std_logic;
signal \N__17641\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17627\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17612\ : std_logic;
signal \N__17609\ : std_logic;
signal \N__17606\ : std_logic;
signal \N__17603\ : std_logic;
signal \N__17600\ : std_logic;
signal \N__17597\ : std_logic;
signal \N__17594\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17582\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17565\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17563\ : std_logic;
signal \N__17562\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17559\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17556\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17554\ : std_logic;
signal \N__17553\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17551\ : std_logic;
signal \N__17550\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17548\ : std_logic;
signal \N__17547\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17545\ : std_logic;
signal \N__17544\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17533\ : std_logic;
signal \N__17532\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17530\ : std_logic;
signal \N__17529\ : std_logic;
signal \N__17524\ : std_logic;
signal \N__17515\ : std_logic;
signal \N__17506\ : std_logic;
signal \N__17497\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17479\ : std_logic;
signal \N__17476\ : std_logic;
signal \N__17467\ : std_logic;
signal \N__17464\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17452\ : std_logic;
signal \N__17441\ : std_logic;
signal \N__17438\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17428\ : std_logic;
signal \N__17425\ : std_logic;
signal \N__17422\ : std_logic;
signal \N__17417\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17413\ : std_logic;
signal \N__17410\ : std_logic;
signal \N__17407\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17392\ : std_logic;
signal \N__17389\ : std_logic;
signal \N__17388\ : std_logic;
signal \N__17383\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17365\ : std_logic;
signal \N__17362\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17348\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17344\ : std_logic;
signal \N__17341\ : std_logic;
signal \N__17338\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17332\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17324\ : std_logic;
signal \N__17321\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17315\ : std_logic;
signal \N__17312\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17297\ : std_logic;
signal \N__17294\ : std_logic;
signal \N__17291\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17276\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17265\ : std_logic;
signal \N__17264\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17258\ : std_logic;
signal \N__17255\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17243\ : std_logic;
signal \N__17240\ : std_logic;
signal \N__17237\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17233\ : std_logic;
signal \N__17232\ : std_logic;
signal \N__17229\ : std_logic;
signal \N__17226\ : std_logic;
signal \N__17223\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17212\ : std_logic;
signal \N__17211\ : std_logic;
signal \N__17208\ : std_logic;
signal \N__17205\ : std_logic;
signal \N__17202\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17194\ : std_logic;
signal \N__17193\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17177\ : std_logic;
signal \N__17174\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17168\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17162\ : std_logic;
signal \N__17159\ : std_logic;
signal \N__17156\ : std_logic;
signal \N__17153\ : std_logic;
signal \N__17150\ : std_logic;
signal \N__17147\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17141\ : std_logic;
signal \N__17138\ : std_logic;
signal \N__17135\ : std_logic;
signal \N__17132\ : std_logic;
signal \N__17129\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17123\ : std_logic;
signal \N__17120\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17114\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17107\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17099\ : std_logic;
signal \N__17096\ : std_logic;
signal \N__17093\ : std_logic;
signal \N__17092\ : std_logic;
signal \N__17089\ : std_logic;
signal \N__17086\ : std_logic;
signal \N__17085\ : std_logic;
signal \N__17082\ : std_logic;
signal \N__17079\ : std_logic;
signal \N__17076\ : std_logic;
signal \N__17069\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17065\ : std_logic;
signal \N__17062\ : std_logic;
signal \N__17061\ : std_logic;
signal \N__17058\ : std_logic;
signal \N__17055\ : std_logic;
signal \N__17052\ : std_logic;
signal \N__17049\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17039\ : std_logic;
signal \N__17038\ : std_logic;
signal \N__17035\ : std_logic;
signal \N__17032\ : std_logic;
signal \N__17031\ : std_logic;
signal \N__17026\ : std_logic;
signal \N__17023\ : std_logic;
signal \N__17022\ : std_logic;
signal \N__17017\ : std_logic;
signal \N__17016\ : std_logic;
signal \N__17013\ : std_logic;
signal \N__17010\ : std_logic;
signal \N__17007\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16999\ : std_logic;
signal \N__16998\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16996\ : std_logic;
signal \N__16995\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16987\ : std_logic;
signal \N__16984\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16966\ : std_logic;
signal \N__16965\ : std_logic;
signal \N__16964\ : std_logic;
signal \N__16963\ : std_logic;
signal \N__16960\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16952\ : std_logic;
signal \N__16949\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16934\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16927\ : std_logic;
signal \N__16924\ : std_logic;
signal \N__16921\ : std_logic;
signal \N__16920\ : std_logic;
signal \N__16915\ : std_logic;
signal \N__16912\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16901\ : std_logic;
signal \N__16898\ : std_logic;
signal \N__16895\ : std_logic;
signal \N__16892\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16890\ : std_logic;
signal \N__16889\ : std_logic;
signal \N__16886\ : std_logic;
signal \N__16883\ : std_logic;
signal \N__16880\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16869\ : std_logic;
signal \N__16866\ : std_logic;
signal \N__16859\ : std_logic;
signal \N__16856\ : std_logic;
signal \N__16853\ : std_logic;
signal \N__16850\ : std_logic;
signal \N__16847\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16832\ : std_logic;
signal \N__16829\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16820\ : std_logic;
signal \N__16819\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16813\ : std_logic;
signal \N__16808\ : std_logic;
signal \N__16807\ : std_logic;
signal \N__16804\ : std_logic;
signal \N__16801\ : std_logic;
signal \N__16796\ : std_logic;
signal \N__16793\ : std_logic;
signal \N__16792\ : std_logic;
signal \N__16789\ : std_logic;
signal \N__16786\ : std_logic;
signal \N__16783\ : std_logic;
signal \N__16782\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16766\ : std_logic;
signal \N__16761\ : std_logic;
signal \N__16754\ : std_logic;
signal \N__16751\ : std_logic;
signal \N__16750\ : std_logic;
signal \N__16747\ : std_logic;
signal \N__16744\ : std_logic;
signal \N__16741\ : std_logic;
signal \N__16738\ : std_logic;
signal \N__16737\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16730\ : std_logic;
signal \N__16727\ : std_logic;
signal \N__16724\ : std_logic;
signal \N__16715\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16711\ : std_logic;
signal \N__16708\ : std_logic;
signal \N__16705\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16699\ : std_logic;
signal \N__16698\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16688\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16672\ : std_logic;
signal \N__16669\ : std_logic;
signal \N__16666\ : std_logic;
signal \N__16665\ : std_logic;
signal \N__16660\ : std_logic;
signal \N__16657\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16645\ : std_logic;
signal \N__16642\ : std_logic;
signal \N__16639\ : std_logic;
signal \N__16638\ : std_logic;
signal \N__16635\ : std_logic;
signal \N__16632\ : std_logic;
signal \N__16629\ : std_logic;
signal \N__16622\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16618\ : std_logic;
signal \N__16615\ : std_logic;
signal \N__16612\ : std_logic;
signal \N__16611\ : std_logic;
signal \N__16606\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16600\ : std_logic;
signal \N__16597\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16589\ : std_logic;
signal \N__16588\ : std_logic;
signal \N__16585\ : std_logic;
signal \N__16582\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16576\ : std_logic;
signal \N__16573\ : std_logic;
signal \N__16570\ : std_logic;
signal \N__16565\ : std_logic;
signal \N__16564\ : std_logic;
signal \N__16561\ : std_logic;
signal \N__16558\ : std_logic;
signal \N__16555\ : std_logic;
signal \N__16552\ : std_logic;
signal \N__16549\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16543\ : std_logic;
signal \N__16540\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16531\ : std_logic;
signal \N__16528\ : std_logic;
signal \N__16525\ : std_logic;
signal \N__16522\ : std_logic;
signal \N__16519\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16515\ : std_logic;
signal \N__16510\ : std_logic;
signal \N__16507\ : std_logic;
signal \N__16504\ : std_logic;
signal \N__16501\ : std_logic;
signal \N__16496\ : std_logic;
signal \N__16493\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16487\ : std_logic;
signal \N__16484\ : std_logic;
signal \N__16483\ : std_logic;
signal \N__16480\ : std_logic;
signal \N__16477\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16471\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16456\ : std_logic;
signal \N__16453\ : std_logic;
signal \N__16450\ : std_logic;
signal \N__16449\ : std_logic;
signal \N__16446\ : std_logic;
signal \N__16443\ : std_logic;
signal \N__16440\ : std_logic;
signal \N__16437\ : std_logic;
signal \N__16432\ : std_logic;
signal \N__16429\ : std_logic;
signal \N__16426\ : std_logic;
signal \N__16421\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16411\ : std_logic;
signal \N__16408\ : std_logic;
signal \N__16405\ : std_logic;
signal \N__16402\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16395\ : std_logic;
signal \N__16392\ : std_logic;
signal \N__16389\ : std_logic;
signal \N__16386\ : std_logic;
signal \N__16383\ : std_logic;
signal \N__16376\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16374\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16365\ : std_logic;
signal \N__16360\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16352\ : std_logic;
signal \N__16351\ : std_logic;
signal \N__16350\ : std_logic;
signal \N__16347\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16336\ : std_logic;
signal \N__16331\ : std_logic;
signal \N__16328\ : std_logic;
signal \N__16327\ : std_logic;
signal \N__16326\ : std_logic;
signal \N__16323\ : std_logic;
signal \N__16320\ : std_logic;
signal \N__16317\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16307\ : std_logic;
signal \N__16306\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16302\ : std_logic;
signal \N__16299\ : std_logic;
signal \N__16296\ : std_logic;
signal \N__16289\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16282\ : std_logic;
signal \N__16279\ : std_logic;
signal \N__16274\ : std_logic;
signal \N__16273\ : std_logic;
signal \N__16272\ : std_logic;
signal \N__16269\ : std_logic;
signal \N__16266\ : std_logic;
signal \N__16263\ : std_logic;
signal \N__16258\ : std_logic;
signal \N__16253\ : std_logic;
signal \N__16250\ : std_logic;
signal \N__16249\ : std_logic;
signal \N__16246\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16238\ : std_logic;
signal \N__16237\ : std_logic;
signal \N__16236\ : std_logic;
signal \N__16233\ : std_logic;
signal \N__16230\ : std_logic;
signal \N__16227\ : std_logic;
signal \N__16222\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16214\ : std_logic;
signal \N__16211\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16209\ : std_logic;
signal \N__16206\ : std_logic;
signal \N__16203\ : std_logic;
signal \N__16200\ : std_logic;
signal \N__16195\ : std_logic;
signal \N__16190\ : std_logic;
signal \N__16187\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16182\ : std_logic;
signal \N__16179\ : std_logic;
signal \N__16176\ : std_logic;
signal \N__16171\ : std_logic;
signal \N__16166\ : std_logic;
signal \N__16163\ : std_logic;
signal \N__16162\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16158\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16145\ : std_logic;
signal \N__16142\ : std_logic;
signal \N__16141\ : std_logic;
signal \N__16140\ : std_logic;
signal \N__16137\ : std_logic;
signal \N__16134\ : std_logic;
signal \N__16131\ : std_logic;
signal \N__16124\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16119\ : std_logic;
signal \N__16116\ : std_logic;
signal \N__16113\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16105\ : std_logic;
signal \N__16100\ : std_logic;
signal \N__16097\ : std_logic;
signal \N__16096\ : std_logic;
signal \N__16095\ : std_logic;
signal \N__16092\ : std_logic;
signal \N__16089\ : std_logic;
signal \N__16086\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16076\ : std_logic;
signal \N__16073\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16071\ : std_logic;
signal \N__16068\ : std_logic;
signal \N__16063\ : std_logic;
signal \N__16058\ : std_logic;
signal \N__16055\ : std_logic;
signal \N__16054\ : std_logic;
signal \N__16053\ : std_logic;
signal \N__16050\ : std_logic;
signal \N__16045\ : std_logic;
signal \N__16040\ : std_logic;
signal \N__16037\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16035\ : std_logic;
signal \N__16032\ : std_logic;
signal \N__16027\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16019\ : std_logic;
signal \N__16018\ : std_logic;
signal \N__16017\ : std_logic;
signal \N__16014\ : std_logic;
signal \N__16011\ : std_logic;
signal \N__16008\ : std_logic;
signal \N__16003\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15987\ : std_logic;
signal \N__15984\ : std_logic;
signal \N__15979\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15971\ : std_logic;
signal \N__15970\ : std_logic;
signal \N__15969\ : std_logic;
signal \N__15966\ : std_logic;
signal \N__15963\ : std_logic;
signal \N__15960\ : std_logic;
signal \N__15953\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15949\ : std_logic;
signal \N__15948\ : std_logic;
signal \N__15945\ : std_logic;
signal \N__15942\ : std_logic;
signal \N__15939\ : std_logic;
signal \N__15932\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15928\ : std_logic;
signal \N__15927\ : std_logic;
signal \N__15924\ : std_logic;
signal \N__15921\ : std_logic;
signal \N__15918\ : std_logic;
signal \N__15913\ : std_logic;
signal \N__15908\ : std_logic;
signal \N__15905\ : std_logic;
signal \N__15904\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15900\ : std_logic;
signal \N__15897\ : std_logic;
signal \N__15894\ : std_logic;
signal \N__15889\ : std_logic;
signal \N__15884\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15880\ : std_logic;
signal \N__15879\ : std_logic;
signal \N__15876\ : std_logic;
signal \N__15871\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15863\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15861\ : std_logic;
signal \N__15858\ : std_logic;
signal \N__15853\ : std_logic;
signal \N__15848\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15843\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15833\ : std_logic;
signal \N__15832\ : std_logic;
signal \N__15831\ : std_logic;
signal \N__15830\ : std_logic;
signal \N__15829\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15816\ : std_logic;
signal \N__15813\ : std_logic;
signal \N__15810\ : std_logic;
signal \N__15803\ : std_logic;
signal \N__15802\ : std_logic;
signal \N__15801\ : std_logic;
signal \N__15800\ : std_logic;
signal \N__15799\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15791\ : std_logic;
signal \N__15786\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15776\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15772\ : std_logic;
signal \N__15771\ : std_logic;
signal \N__15768\ : std_logic;
signal \N__15765\ : std_logic;
signal \N__15762\ : std_logic;
signal \N__15759\ : std_logic;
signal \N__15756\ : std_logic;
signal \N__15753\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15743\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15739\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15732\ : std_logic;
signal \N__15729\ : std_logic;
signal \N__15726\ : std_logic;
signal \N__15723\ : std_logic;
signal \N__15720\ : std_logic;
signal \N__15717\ : std_logic;
signal \N__15714\ : std_logic;
signal \N__15707\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15703\ : std_logic;
signal \N__15700\ : std_logic;
signal \N__15699\ : std_logic;
signal \N__15696\ : std_logic;
signal \N__15695\ : std_logic;
signal \N__15692\ : std_logic;
signal \N__15689\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15683\ : std_logic;
signal \N__15678\ : std_logic;
signal \N__15671\ : std_logic;
signal \N__15668\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15662\ : std_logic;
signal \N__15659\ : std_logic;
signal \N__15658\ : std_logic;
signal \N__15657\ : std_logic;
signal \N__15654\ : std_logic;
signal \N__15651\ : std_logic;
signal \N__15648\ : std_logic;
signal \N__15643\ : std_logic;
signal \N__15638\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15634\ : std_logic;
signal \N__15633\ : std_logic;
signal \N__15630\ : std_logic;
signal \N__15627\ : std_logic;
signal \N__15624\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15614\ : std_logic;
signal \N__15611\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15609\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15601\ : std_logic;
signal \N__15596\ : std_logic;
signal \N__15593\ : std_logic;
signal \N__15590\ : std_logic;
signal \N__15589\ : std_logic;
signal \N__15584\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15578\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15572\ : std_logic;
signal \N__15569\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15559\ : std_logic;
signal \N__15554\ : std_logic;
signal \N__15551\ : std_logic;
signal \N__15548\ : std_logic;
signal \N__15545\ : std_logic;
signal \N__15542\ : std_logic;
signal \N__15539\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15537\ : std_logic;
signal \N__15534\ : std_logic;
signal \N__15533\ : std_logic;
signal \N__15532\ : std_logic;
signal \N__15531\ : std_logic;
signal \N__15530\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15524\ : std_logic;
signal \N__15517\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15509\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15499\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15492\ : std_logic;
signal \N__15489\ : std_logic;
signal \N__15482\ : std_logic;
signal \N__15479\ : std_logic;
signal \N__15478\ : std_logic;
signal \N__15475\ : std_logic;
signal \N__15472\ : std_logic;
signal \N__15471\ : std_logic;
signal \N__15470\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15468\ : std_logic;
signal \N__15467\ : std_logic;
signal \N__15466\ : std_logic;
signal \N__15463\ : std_logic;
signal \N__15460\ : std_logic;
signal \N__15459\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15456\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15454\ : std_logic;
signal \N__15453\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15437\ : std_logic;
signal \N__15436\ : std_logic;
signal \N__15435\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15433\ : std_logic;
signal \N__15432\ : std_logic;
signal \N__15429\ : std_logic;
signal \N__15426\ : std_logic;
signal \N__15421\ : std_logic;
signal \N__15420\ : std_logic;
signal \N__15405\ : std_logic;
signal \N__15402\ : std_logic;
signal \N__15399\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15395\ : std_logic;
signal \N__15392\ : std_logic;
signal \N__15385\ : std_logic;
signal \N__15382\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15367\ : std_logic;
signal \N__15364\ : std_logic;
signal \N__15347\ : std_logic;
signal \N__15346\ : std_logic;
signal \N__15345\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15343\ : std_logic;
signal \N__15342\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15338\ : std_logic;
signal \N__15337\ : std_logic;
signal \N__15336\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15334\ : std_logic;
signal \N__15331\ : std_logic;
signal \N__15330\ : std_logic;
signal \N__15327\ : std_logic;
signal \N__15324\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15320\ : std_logic;
signal \N__15319\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15317\ : std_logic;
signal \N__15316\ : std_logic;
signal \N__15313\ : std_logic;
signal \N__15310\ : std_logic;
signal \N__15307\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15305\ : std_logic;
signal \N__15304\ : std_logic;
signal \N__15303\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15297\ : std_logic;
signal \N__15294\ : std_logic;
signal \N__15291\ : std_logic;
signal \N__15286\ : std_logic;
signal \N__15285\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15275\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15259\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15235\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15227\ : std_logic;
signal \N__15222\ : std_logic;
signal \N__15221\ : std_logic;
signal \N__15218\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15212\ : std_logic;
signal \N__15209\ : std_logic;
signal \N__15204\ : std_logic;
signal \N__15201\ : std_logic;
signal \N__15196\ : std_logic;
signal \N__15185\ : std_logic;
signal \N__15184\ : std_logic;
signal \N__15181\ : std_logic;
signal \N__15178\ : std_logic;
signal \N__15177\ : std_logic;
signal \N__15172\ : std_logic;
signal \N__15169\ : std_logic;
signal \N__15168\ : std_logic;
signal \N__15167\ : std_logic;
signal \N__15164\ : std_logic;
signal \N__15161\ : std_logic;
signal \N__15156\ : std_logic;
signal \N__15149\ : std_logic;
signal \N__15148\ : std_logic;
signal \N__15147\ : std_logic;
signal \N__15146\ : std_logic;
signal \N__15145\ : std_logic;
signal \N__15144\ : std_logic;
signal \N__15143\ : std_logic;
signal \N__15142\ : std_logic;
signal \N__15141\ : std_logic;
signal \N__15140\ : std_logic;
signal \N__15137\ : std_logic;
signal \N__15136\ : std_logic;
signal \N__15135\ : std_logic;
signal \N__15134\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15131\ : std_logic;
signal \N__15130\ : std_logic;
signal \N__15129\ : std_logic;
signal \N__15124\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15108\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15105\ : std_logic;
signal \N__15104\ : std_logic;
signal \N__15103\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15078\ : std_logic;
signal \N__15075\ : std_logic;
signal \N__15074\ : std_logic;
signal \N__15071\ : std_logic;
signal \N__15068\ : std_logic;
signal \N__15063\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15051\ : std_logic;
signal \N__15048\ : std_logic;
signal \N__15035\ : std_logic;
signal \N__15034\ : std_logic;
signal \N__15031\ : std_logic;
signal \N__15028\ : std_logic;
signal \N__15025\ : std_logic;
signal \N__15022\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15014\ : std_logic;
signal \N__15011\ : std_logic;
signal \N__15008\ : std_logic;
signal \N__15005\ : std_logic;
signal \N__15002\ : std_logic;
signal \N__15001\ : std_logic;
signal \N__15000\ : std_logic;
signal \N__14997\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14987\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14983\ : std_logic;
signal \N__14980\ : std_logic;
signal \N__14977\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14969\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14963\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14959\ : std_logic;
signal \N__14956\ : std_logic;
signal \N__14953\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14936\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14932\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14921\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14915\ : std_logic;
signal \N__14912\ : std_logic;
signal \N__14911\ : std_logic;
signal \N__14908\ : std_logic;
signal \N__14905\ : std_logic;
signal \N__14902\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14894\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14888\ : std_logic;
signal \N__14887\ : std_logic;
signal \N__14884\ : std_logic;
signal \N__14881\ : std_logic;
signal \N__14880\ : std_logic;
signal \N__14879\ : std_logic;
signal \N__14876\ : std_logic;
signal \N__14873\ : std_logic;
signal \N__14868\ : std_logic;
signal \N__14865\ : std_logic;
signal \N__14862\ : std_logic;
signal \N__14859\ : std_logic;
signal \N__14852\ : std_logic;
signal \N__14849\ : std_logic;
signal \N__14848\ : std_logic;
signal \N__14847\ : std_logic;
signal \N__14846\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14836\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14827\ : std_logic;
signal \N__14826\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14824\ : std_logic;
signal \N__14823\ : std_logic;
signal \N__14816\ : std_logic;
signal \N__14815\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14807\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14799\ : std_logic;
signal \N__14798\ : std_logic;
signal \N__14795\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14788\ : std_logic;
signal \N__14775\ : std_logic;
signal \N__14772\ : std_logic;
signal \N__14769\ : std_logic;
signal \N__14766\ : std_logic;
signal \N__14759\ : std_logic;
signal \N__14758\ : std_logic;
signal \N__14757\ : std_logic;
signal \N__14756\ : std_logic;
signal \N__14751\ : std_logic;
signal \N__14746\ : std_logic;
signal \N__14745\ : std_logic;
signal \N__14742\ : std_logic;
signal \N__14739\ : std_logic;
signal \N__14736\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14722\ : std_logic;
signal \N__14721\ : std_logic;
signal \N__14720\ : std_logic;
signal \N__14719\ : std_logic;
signal \N__14718\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14716\ : std_logic;
signal \N__14709\ : std_logic;
signal \N__14698\ : std_logic;
signal \N__14697\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14695\ : std_logic;
signal \N__14694\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14692\ : std_logic;
signal \N__14691\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14667\ : std_logic;
signal \N__14664\ : std_logic;
signal \N__14661\ : std_logic;
signal \N__14658\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14650\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14636\ : std_logic;
signal \N__14633\ : std_logic;
signal \N__14630\ : std_logic;
signal \N__14627\ : std_logic;
signal \N__14624\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14620\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14600\ : std_logic;
signal \N__14597\ : std_logic;
signal \N__14596\ : std_logic;
signal \N__14593\ : std_logic;
signal \N__14590\ : std_logic;
signal \N__14587\ : std_logic;
signal \N__14582\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14576\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14560\ : std_logic;
signal \N__14555\ : std_logic;
signal \N__14552\ : std_logic;
signal \N__14549\ : std_logic;
signal \N__14546\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14528\ : std_logic;
signal \N__14525\ : std_logic;
signal \N__14522\ : std_logic;
signal \N__14519\ : std_logic;
signal \N__14516\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14498\ : std_logic;
signal \N__14495\ : std_logic;
signal \N__14492\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14485\ : std_logic;
signal \N__14482\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14474\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14468\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14464\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14458\ : std_logic;
signal \N__14455\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14444\ : std_logic;
signal \N__14441\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14433\ : std_logic;
signal \N__14430\ : std_logic;
signal \N__14427\ : std_logic;
signal \N__14424\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14411\ : std_logic;
signal \N__14408\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14402\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14381\ : std_logic;
signal \N__14378\ : std_logic;
signal \N__14375\ : std_logic;
signal \N__14372\ : std_logic;
signal \N__14369\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14357\ : std_logic;
signal \N__14354\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14348\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14342\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14336\ : std_logic;
signal \N__14333\ : std_logic;
signal \N__14330\ : std_logic;
signal \N__14327\ : std_logic;
signal \N__14324\ : std_logic;
signal \N__14321\ : std_logic;
signal \N__14320\ : std_logic;
signal \N__14317\ : std_logic;
signal \N__14314\ : std_logic;
signal \N__14309\ : std_logic;
signal \N__14306\ : std_logic;
signal \N__14303\ : std_logic;
signal \N__14300\ : std_logic;
signal \N__14297\ : std_logic;
signal \N__14294\ : std_logic;
signal \N__14291\ : std_logic;
signal \N__14288\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14281\ : std_logic;
signal \N__14276\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14264\ : std_logic;
signal \N__14261\ : std_logic;
signal \N__14258\ : std_logic;
signal \N__14255\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14243\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14231\ : std_logic;
signal \N__14228\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14215\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14207\ : std_logic;
signal \N__14204\ : std_logic;
signal \N__14201\ : std_logic;
signal \N__14198\ : std_logic;
signal \N__14195\ : std_logic;
signal \N__14192\ : std_logic;
signal \N__14189\ : std_logic;
signal \N__14186\ : std_logic;
signal \N__14183\ : std_logic;
signal \N__14180\ : std_logic;
signal \N__14177\ : std_logic;
signal \N__14174\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14172\ : std_logic;
signal \N__14171\ : std_logic;
signal \N__14162\ : std_logic;
signal \N__14159\ : std_logic;
signal \N__14156\ : std_logic;
signal \N__14153\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14147\ : std_logic;
signal \N__14144\ : std_logic;
signal \N__14141\ : std_logic;
signal \N__14138\ : std_logic;
signal \N__14135\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14129\ : std_logic;
signal \N__14126\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14120\ : std_logic;
signal \N__14117\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14111\ : std_logic;
signal \N__14108\ : std_logic;
signal \N__14105\ : std_logic;
signal \N__14102\ : std_logic;
signal \N__14099\ : std_logic;
signal \N__14096\ : std_logic;
signal \N__14095\ : std_logic;
signal \N__14092\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14088\ : std_logic;
signal \N__14085\ : std_logic;
signal \N__14082\ : std_logic;
signal \N__14079\ : std_logic;
signal \N__14076\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14066\ : std_logic;
signal \N__14063\ : std_logic;
signal \N__14062\ : std_logic;
signal \N__14061\ : std_logic;
signal \N__14058\ : std_logic;
signal \N__14055\ : std_logic;
signal \N__14054\ : std_logic;
signal \N__14051\ : std_logic;
signal \N__14048\ : std_logic;
signal \N__14045\ : std_logic;
signal \N__14042\ : std_logic;
signal \N__14039\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14029\ : std_logic;
signal \N__14024\ : std_logic;
signal \N__14021\ : std_logic;
signal \N__14020\ : std_logic;
signal \N__14019\ : std_logic;
signal \N__14016\ : std_logic;
signal \N__14015\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14009\ : std_logic;
signal \N__14006\ : std_logic;
signal \N__14003\ : std_logic;
signal \N__14000\ : std_logic;
signal \N__13997\ : std_logic;
signal \N__13994\ : std_logic;
signal \N__13991\ : std_logic;
signal \N__13986\ : std_logic;
signal \N__13979\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13974\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13970\ : std_logic;
signal \N__13967\ : std_logic;
signal \N__13966\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13958\ : std_logic;
signal \N__13955\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13942\ : std_logic;
signal \N__13939\ : std_logic;
signal \N__13934\ : std_logic;
signal \N__13933\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13926\ : std_logic;
signal \N__13923\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13919\ : std_logic;
signal \N__13916\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13910\ : std_logic;
signal \N__13907\ : std_logic;
signal \N__13904\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13893\ : std_logic;
signal \N__13888\ : std_logic;
signal \N__13883\ : std_logic;
signal \N__13882\ : std_logic;
signal \N__13881\ : std_logic;
signal \N__13878\ : std_logic;
signal \N__13875\ : std_logic;
signal \N__13872\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13863\ : std_logic;
signal \N__13860\ : std_logic;
signal \N__13857\ : std_logic;
signal \N__13854\ : std_logic;
signal \N__13847\ : std_logic;
signal \N__13846\ : std_logic;
signal \N__13843\ : std_logic;
signal \N__13842\ : std_logic;
signal \N__13839\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13832\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13826\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13808\ : std_logic;
signal \N__13805\ : std_logic;
signal \N__13802\ : std_logic;
signal \N__13799\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13791\ : std_logic;
signal \N__13788\ : std_logic;
signal \N__13785\ : std_logic;
signal \N__13782\ : std_logic;
signal \N__13775\ : std_logic;
signal \N__13772\ : std_logic;
signal \N__13769\ : std_logic;
signal \N__13768\ : std_logic;
signal \N__13765\ : std_logic;
signal \N__13762\ : std_logic;
signal \N__13761\ : std_logic;
signal \N__13758\ : std_logic;
signal \N__13755\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13745\ : std_logic;
signal \N__13742\ : std_logic;
signal \N__13741\ : std_logic;
signal \N__13738\ : std_logic;
signal \N__13735\ : std_logic;
signal \N__13732\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13719\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13713\ : std_logic;
signal \N__13708\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13700\ : std_logic;
signal \N__13699\ : std_logic;
signal \N__13696\ : std_logic;
signal \N__13693\ : std_logic;
signal \N__13692\ : std_logic;
signal \N__13689\ : std_logic;
signal \N__13686\ : std_logic;
signal \N__13683\ : std_logic;
signal \N__13676\ : std_logic;
signal \N__13673\ : std_logic;
signal \N__13672\ : std_logic;
signal \N__13671\ : std_logic;
signal \N__13670\ : std_logic;
signal \N__13669\ : std_logic;
signal \N__13666\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13652\ : std_logic;
signal \N__13649\ : std_logic;
signal \N__13648\ : std_logic;
signal \N__13645\ : std_logic;
signal \N__13642\ : std_logic;
signal \N__13639\ : std_logic;
signal \N__13636\ : std_logic;
signal \N__13633\ : std_logic;
signal \N__13630\ : std_logic;
signal \N__13627\ : std_logic;
signal \N__13624\ : std_logic;
signal \N__13619\ : std_logic;
signal \N__13618\ : std_logic;
signal \N__13615\ : std_logic;
signal \N__13612\ : std_logic;
signal \N__13611\ : std_logic;
signal \N__13608\ : std_logic;
signal \N__13605\ : std_logic;
signal \N__13602\ : std_logic;
signal \N__13599\ : std_logic;
signal \N__13594\ : std_logic;
signal \N__13589\ : std_logic;
signal \N__13586\ : std_logic;
signal \N__13585\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13581\ : std_logic;
signal \N__13578\ : std_logic;
signal \N__13575\ : std_logic;
signal \N__13572\ : std_logic;
signal \N__13569\ : std_logic;
signal \N__13566\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13555\ : std_logic;
signal \N__13554\ : std_logic;
signal \N__13553\ : std_logic;
signal \N__13552\ : std_logic;
signal \N__13551\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13543\ : std_logic;
signal \N__13542\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13540\ : std_logic;
signal \N__13537\ : std_logic;
signal \N__13530\ : std_logic;
signal \N__13527\ : std_logic;
signal \N__13522\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13507\ : std_logic;
signal \N__13502\ : std_logic;
signal \N__13499\ : std_logic;
signal \N__13498\ : std_logic;
signal \N__13495\ : std_logic;
signal \N__13492\ : std_logic;
signal \N__13491\ : std_logic;
signal \N__13490\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13458\ : std_logic;
signal \N__13455\ : std_logic;
signal \N__13452\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13421\ : std_logic;
signal \N__13418\ : std_logic;
signal \N__13417\ : std_logic;
signal \N__13416\ : std_logic;
signal \N__13413\ : std_logic;
signal \N__13410\ : std_logic;
signal \N__13407\ : std_logic;
signal \N__13404\ : std_logic;
signal \N__13401\ : std_logic;
signal \N__13398\ : std_logic;
signal \N__13395\ : std_logic;
signal \N__13392\ : std_logic;
signal \N__13389\ : std_logic;
signal \N__13382\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13378\ : std_logic;
signal \N__13377\ : std_logic;
signal \N__13374\ : std_logic;
signal \N__13371\ : std_logic;
signal \N__13368\ : std_logic;
signal \N__13365\ : std_logic;
signal \N__13362\ : std_logic;
signal \N__13359\ : std_logic;
signal \N__13356\ : std_logic;
signal \N__13353\ : std_logic;
signal \N__13350\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13336\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13332\ : std_logic;
signal \N__13329\ : std_logic;
signal \N__13326\ : std_logic;
signal \N__13323\ : std_logic;
signal \N__13320\ : std_logic;
signal \N__13317\ : std_logic;
signal \N__13314\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13303\ : std_logic;
signal \N__13302\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13294\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13288\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13282\ : std_logic;
signal \N__13281\ : std_logic;
signal \N__13278\ : std_logic;
signal \N__13275\ : std_logic;
signal \N__13272\ : std_logic;
signal \N__13267\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13244\ : std_logic;
signal \N__13241\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13235\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13216\ : std_logic;
signal \N__13213\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13204\ : std_logic;
signal \N__13201\ : std_logic;
signal \N__13198\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13187\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13181\ : std_logic;
signal \N__13178\ : std_logic;
signal \N__13175\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13169\ : std_logic;
signal \N__13166\ : std_logic;
signal \N__13163\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13159\ : std_logic;
signal \N__13154\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13150\ : std_logic;
signal \N__13147\ : std_logic;
signal \N__13144\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13138\ : std_logic;
signal \N__13133\ : std_logic;
signal \N__13130\ : std_logic;
signal \N__13127\ : std_logic;
signal \N__13126\ : std_logic;
signal \N__13125\ : std_logic;
signal \N__13122\ : std_logic;
signal \N__13119\ : std_logic;
signal \N__13116\ : std_logic;
signal \N__13113\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13105\ : std_logic;
signal \N__13102\ : std_logic;
signal \N__13099\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13093\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13085\ : std_logic;
signal \N__13084\ : std_logic;
signal \N__13083\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13075\ : std_logic;
signal \N__13072\ : std_logic;
signal \N__13071\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13065\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13059\ : std_logic;
signal \N__13058\ : std_logic;
signal \N__13057\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13035\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13025\ : std_logic;
signal \N__13022\ : std_logic;
signal \N__13019\ : std_logic;
signal \N__13016\ : std_logic;
signal \N__13015\ : std_logic;
signal \N__13014\ : std_logic;
signal \N__13011\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13005\ : std_logic;
signal \N__13002\ : std_logic;
signal \N__12997\ : std_logic;
signal \N__12992\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12983\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12974\ : std_logic;
signal \N__12971\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12965\ : std_logic;
signal \N__12962\ : std_logic;
signal \N__12961\ : std_logic;
signal \N__12960\ : std_logic;
signal \N__12955\ : std_logic;
signal \N__12952\ : std_logic;
signal \N__12947\ : std_logic;
signal \N__12944\ : std_logic;
signal \N__12941\ : std_logic;
signal \N__12940\ : std_logic;
signal \N__12937\ : std_logic;
signal \N__12936\ : std_logic;
signal \N__12931\ : std_logic;
signal \N__12928\ : std_logic;
signal \N__12927\ : std_logic;
signal \N__12924\ : std_logic;
signal \N__12919\ : std_logic;
signal \N__12914\ : std_logic;
signal \N__12913\ : std_logic;
signal \N__12912\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12910\ : std_logic;
signal \N__12909\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12907\ : std_logic;
signal \N__12906\ : std_logic;
signal \N__12905\ : std_logic;
signal \N__12904\ : std_logic;
signal \N__12903\ : std_logic;
signal \N__12902\ : std_logic;
signal \N__12899\ : std_logic;
signal \N__12896\ : std_logic;
signal \N__12893\ : std_logic;
signal \N__12892\ : std_logic;
signal \N__12889\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12885\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12880\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12869\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12863\ : std_logic;
signal \N__12862\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12858\ : std_logic;
signal \N__12855\ : std_logic;
signal \N__12854\ : std_logic;
signal \N__12853\ : std_logic;
signal \N__12844\ : std_logic;
signal \N__12835\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12813\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12803\ : std_logic;
signal \N__12800\ : std_logic;
signal \N__12799\ : std_logic;
signal \N__12794\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12777\ : std_logic;
signal \N__12774\ : std_logic;
signal \N__12769\ : std_logic;
signal \N__12764\ : std_logic;
signal \N__12755\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12740\ : std_logic;
signal \N__12737\ : std_logic;
signal \N__12736\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12728\ : std_logic;
signal \N__12727\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12724\ : std_logic;
signal \N__12723\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12721\ : std_logic;
signal \N__12718\ : std_logic;
signal \N__12707\ : std_logic;
signal \N__12702\ : std_logic;
signal \N__12695\ : std_logic;
signal \N__12692\ : std_logic;
signal \N__12689\ : std_logic;
signal \N__12686\ : std_logic;
signal \N__12683\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12677\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12668\ : std_logic;
signal \N__12667\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12660\ : std_logic;
signal \N__12657\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12649\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12629\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12614\ : std_logic;
signal \N__12611\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12605\ : std_logic;
signal \N__12602\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12596\ : std_logic;
signal \N__12593\ : std_logic;
signal \N__12590\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12578\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12557\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12551\ : std_logic;
signal \N__12548\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12542\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12527\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12518\ : std_logic;
signal \N__12515\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12494\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12488\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12452\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12443\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12428\ : std_logic;
signal \N__12425\ : std_logic;
signal \N__12422\ : std_logic;
signal \N__12419\ : std_logic;
signal \N__12416\ : std_logic;
signal \N__12413\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12404\ : std_logic;
signal \N__12401\ : std_logic;
signal \N__12398\ : std_logic;
signal \N__12395\ : std_logic;
signal \N__12392\ : std_logic;
signal \N__12389\ : std_logic;
signal \N__12386\ : std_logic;
signal \N__12383\ : std_logic;
signal \N__12380\ : std_logic;
signal \N__12379\ : std_logic;
signal \N__12378\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12359\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12355\ : std_logic;
signal \N__12352\ : std_logic;
signal \N__12347\ : std_logic;
signal \N__12346\ : std_logic;
signal \N__12341\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12336\ : std_logic;
signal \N__12333\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12323\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12311\ : std_logic;
signal \N__12308\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12290\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12284\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12272\ : std_logic;
signal \N__12267\ : std_logic;
signal \N__12264\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12253\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12244\ : std_logic;
signal \N__12243\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12238\ : std_logic;
signal \N__12235\ : std_logic;
signal \N__12232\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12229\ : std_logic;
signal \N__12228\ : std_logic;
signal \N__12227\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12220\ : std_logic;
signal \N__12217\ : std_logic;
signal \N__12214\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12193\ : std_logic;
signal \N__12190\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12186\ : std_logic;
signal \N__12185\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12183\ : std_logic;
signal \N__12180\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12171\ : std_logic;
signal \N__12170\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12161\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12128\ : std_logic;
signal \N__12127\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12101\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12043\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12027\ : std_logic;
signal \N__12024\ : std_logic;
signal \N__12021\ : std_logic;
signal \N__12016\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12010\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__11999\ : std_logic;
signal \N__11996\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11992\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11985\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11969\ : std_logic;
signal \N__11966\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11959\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11949\ : std_logic;
signal \N__11942\ : std_logic;
signal \N__11941\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11939\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11937\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11934\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11932\ : std_logic;
signal \N__11929\ : std_logic;
signal \N__11928\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11916\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11903\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11889\ : std_logic;
signal \N__11888\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11817\ : std_logic;
signal \N__11814\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11800\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11786\ : std_logic;
signal \N__11783\ : std_logic;
signal \N__11780\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11733\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11720\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11714\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11696\ : std_logic;
signal \N__11687\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11644\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11635\ : std_logic;
signal \N__11634\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11556\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11534\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11486\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11404\ : std_logic;
signal \N__11403\ : std_logic;
signal \N__11402\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11377\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11330\ : std_logic;
signal \N__11327\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11312\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11294\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11270\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11237\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11159\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11145\ : std_logic;
signal \N__11142\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11133\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11107\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11098\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10979\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10907\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10891\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10882\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10876\ : std_logic;
signal \N__10875\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10873\ : std_logic;
signal \N__10872\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10818\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10806\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10800\ : std_logic;
signal \N__10797\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10780\ : std_logic;
signal \N__10779\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10777\ : std_logic;
signal \N__10776\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10774\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10768\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10765\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10729\ : std_logic;
signal \N__10722\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10711\ : std_logic;
signal \N__10710\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10699\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10690\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10615\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10588\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10522\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10480\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10474\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10466\ : std_logic;
signal \N__10463\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10438\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10366\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10348\ : std_logic;
signal \N__10345\ : std_logic;
signal \N__10342\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10192\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10122\ : std_logic;
signal \N__10119\ : std_logic;
signal \N__10116\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10033\ : std_logic;
signal \N__10030\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9994\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9913\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9907\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9889\ : std_logic;
signal \N__9886\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9871\ : std_logic;
signal \N__9868\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9850\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9788\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9742\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9708\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9699\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9609\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9547\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9474\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9466\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9390\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9384\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9348\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9242\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9176\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9061\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9040\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8860\ : std_logic;
signal \N__8857\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8839\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8372\ : std_logic;
signal \N__8369\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8360\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8312\ : std_logic;
signal \N__8309\ : std_logic;
signal \N__8306\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8273\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8246\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8210\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8198\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \bfn_1_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\ : std_logic;
signal \bfn_1_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\ : std_logic;
signal \bfn_1_16_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\ : std_logic;
signal \bfn_1_17_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\ : std_logic;
signal \bfn_1_18_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\ : std_logic;
signal \bfn_1_19_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \rgb_drv_RNOZ0\ : std_logic;
signal \N_39_i_i\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.time_passed11_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.time_passed11_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\ : std_logic;
signal \bfn_2_23_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7\ : std_logic;
signal \bfn_2_24_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15\ : std_logic;
signal \bfn_2_25_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.time_passed11_cascade_\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_3_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_3_16_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_17\ : std_logic;
signal \bfn_3_17_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_3_19_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_3_20_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_17\ : std_logic;
signal \bfn_3_21_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_3_25_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_3_26_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_17\ : std_logic;
signal \bfn_3_27_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\ : std_logic;
signal clk_12mhz : std_logic;
signal \GB_BUFFER_clk_12mhz_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_tr.time_passed11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_hc.time_passed11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_6_f0_0_a2_4Z0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_6_f0_0_a2_3Z0Z_3_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_144_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_0Z0Z_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2Z0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2Z0Z_9_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_6_i_o2Z0Z_15_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_1Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_1Z0Z_6_cascade_\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_122\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a3_0Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_144\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_o2Z0Z_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_0Z0Z_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_o2Z0Z_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_6_i_o2Z0Z_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa\ : std_logic;
signal \phase_controller_slave.stoper_hc.time_passed11\ : std_logic;
signal \phase_controller_slave.stoper_hc.time_passed_1_sqmuxa\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst1.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst1.N_110\ : std_logic;
signal \phase_controller_inst1.N_112\ : std_logic;
signal \phase_controller_inst1.tr_time_passed\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst1.hc_time_passed\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_4\ : std_logic;
signal \phase_controller_inst1.N_107\ : std_logic;
signal \phase_controller_inst1.start_timer_trZ0\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_5_17_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_5_18_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_17\ : std_logic;
signal \bfn_5_19_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO_cascade_\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_38\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa\ : std_logic;
signal \phase_controller_slave.start_timer_tr_0_sqmuxa\ : std_logic;
signal \phase_controller_slave.tr_time_passed\ : std_logic;
signal \phase_controller_slave.stateZ0Z_0\ : std_logic;
signal \phase_controller_slave.state_RNIVDE2Z0Z_0\ : std_logic;
signal start_stop_c : std_logic;
signal shift_flag_start : std_logic;
signal il_max_comp2_c : std_logic;
signal \il_max_comp2_D1\ : std_logic;
signal \phase_controller_slave.state_RNO_0Z0Z_3\ : std_logic;
signal \il_max_comp2_D2\ : std_logic;
signal \phase_controller_slave.start_timer_hc_0_sqmuxa\ : std_logic;
signal \phase_controller_slave.stateZ0Z_4\ : std_logic;
signal \phase_controller_slave.start_timer_hcZ0\ : std_logic;
signal \phase_controller_slave.stateZ0Z_2\ : std_logic;
signal \phase_controller_slave.hc_time_passed\ : std_logic;
signal \phase_controller_slave.start_timer_hc_RNOZ0Z_0\ : std_logic;
signal il_max_comp1_c : std_logic;
signal il_min_comp2_c : std_logic;
signal \il_max_comp1_D1\ : std_logic;
signal \il_max_comp1_D2\ : std_logic;
signal \phase_controller_inst1.start_timer_hc_0_sqmuxa\ : std_logic;
signal il_min_comp1_c : std_logic;
signal \il_min_comp1_D1\ : std_logic;
signal \il_min_comp1_D2\ : std_logic;
signal \phase_controller_inst1.T01_0_sqmuxa\ : std_logic;
signal \phase_controller_slave.stoper_tr.time_passed_1_sqmuxa\ : std_logic;
signal \il_min_comp2_D1\ : std_logic;
signal \il_min_comp2_D2\ : std_logic;
signal measured_delay_hc_5 : std_logic;
signal measured_delay_hc_2 : std_logic;
signal measured_delay_hc_11 : std_logic;
signal measured_delay_hc_12 : std_logic;
signal measured_delay_hc_3 : std_logic;
signal measured_delay_hc_4 : std_logic;
signal \delay_measurement_inst.delay_hc_reg_3_0_a2_0_6\ : std_logic;
signal measured_delay_hc_1 : std_logic;
signal measured_delay_hc_10 : std_logic;
signal measured_delay_hc_9 : std_logic;
signal measured_delay_hc_15 : std_logic;
signal measured_delay_hc_19 : std_logic;
signal measured_delay_hc_6 : std_logic;
signal measured_delay_hc_17 : std_logic;
signal measured_delay_hc_16 : std_logic;
signal measured_delay_hc_14 : std_logic;
signal measured_delay_hc_18 : std_logic;
signal measured_delay_hc_7 : std_logic;
signal measured_delay_hc_8 : std_logic;
signal \bfn_8_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_7\ : std_logic;
signal \bfn_8_14_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_15\ : std_logic;
signal \bfn_8_15_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_23\ : std_logic;
signal \bfn_8_16_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_256_i_g\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\ : std_logic;
signal \bfn_8_17_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9\ : std_logic;
signal \bfn_8_18_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17\ : std_logic;
signal \bfn_8_19_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_55\ : std_logic;
signal \phase_controller_slave.stoper_tr.time_passed11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_50\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_32\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_32_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_33\ : std_logic;
signal \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_slave.start_timer_trZ0\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_0_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_0_3\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_232_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_6_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_0_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_7\ : std_logic;
signal \delay_measurement_inst.un3_elapsed_time_hc_0_i\ : std_logic;
signal \delay_measurement_inst.un3_elapsed_time_hc_0_i_cascade_\ : std_logic;
signal \delay_measurement_inst.N_219\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_237_cascade_\ : std_logic;
signal \delay_measurement_inst.N_209\ : std_logic;
signal \delay_measurement_inst.N_207\ : std_logic;
signal \delay_measurement_inst.N_207_cascade_\ : std_logic;
signal \delay_measurement_inst.N_243\ : std_logic;
signal \delay_measurement_inst.N_247\ : std_logic;
signal \delay_measurement_inst.N_216_1\ : std_logic;
signal measured_delay_hc_13 : std_logic;
signal \delay_measurement_inst.un3_elapsed_time_hc_0_i_0\ : std_logic;
signal \phase_controller_slave.stateZ0Z_1\ : std_logic;
signal s4_phy_c : std_logic;
signal \bfn_9_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\ : std_logic;
signal \bfn_9_14_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\ : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\ : std_logic;
signal \bfn_9_16_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal measured_delay_tr_1 : std_logic;
signal measured_delay_tr_2 : std_logic;
signal measured_delay_tr_3 : std_logic;
signal measured_delay_tr_6 : std_logic;
signal measured_delay_tr_18 : std_logic;
signal measured_delay_tr_17 : std_logic;
signal measured_delay_tr_16 : std_logic;
signal measured_delay_tr_12 : std_logic;
signal measured_delay_tr_11 : std_logic;
signal measured_delay_tr_13 : std_logic;
signal measured_delay_tr_10 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_0_6\ : std_logic;
signal measured_delay_tr_9 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_0_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_9_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_0_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_97\ : std_logic;
signal measured_delay_tr_4 : std_logic;
signal measured_delay_tr_14 : std_logic;
signal measured_delay_tr_15 : std_logic;
signal measured_delay_tr_5 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_3\ : std_logic;
signal s1_phy_c : std_logic;
signal \bfn_9_21_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_7\ : std_logic;
signal \bfn_9_22_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_15\ : std_logic;
signal \bfn_9_23_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_23\ : std_logic;
signal \bfn_9_24_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_28\ : std_logic;
signal \phase_controller_slave.stateZ0Z_3\ : std_logic;
signal s3_phy_c : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_255_i_g\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.running_i\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_5\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_4\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_3\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_1\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_5_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_177_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3_cascade_\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_16\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_17\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_12\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_11\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_13\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6\ : std_logic;
signal \delay_measurement_inst.N_35_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_7\ : std_logic;
signal \delay_measurement_inst.N_164\ : std_logic;
signal \delay_measurement_inst.N_187\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_7\ : std_logic;
signal \delay_measurement_inst.N_187_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_177\ : std_logic;
signal \delay_measurement_inst.un3_elapsed_time_tr_0_i_cascade_\ : std_logic;
signal \delay_measurement_inst.N_162_1\ : std_logic;
signal \delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_reg3lto9\ : std_logic;
signal \delay_measurement_inst.delay_tr_reg3lto14\ : std_logic;
signal \delay_measurement_inst.N_39\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_180_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_reg3lto6\ : std_logic;
signal \delay_measurement_inst.delay_tr_reg3lto15\ : std_logic;
signal \delay_measurement_inst.delay_tr_reg_5_0_a2_0_6\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_7\ : std_logic;
signal measured_delay_tr_7 : std_logic;
signal \delay_measurement_inst.un3_elapsed_time_tr_0_i\ : std_logic;
signal \delay_measurement_inst.N_41\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_8\ : std_logic;
signal measured_delay_tr_8 : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_31\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_19\ : std_logic;
signal \delay_measurement_inst.N_35\ : std_logic;
signal measured_delay_tr_19 : std_logic;
signal \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_3\ : std_logic;
signal \bfn_10_21_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_11\ : std_logic;
signal \bfn_10_22_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_19\ : std_logic;
signal \bfn_10_23_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\ : std_logic;
signal \bfn_10_24_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_253_i_g\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_255_i\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_1\ : std_logic;
signal s2_phy_c : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_o2_7_19_cascade_\ : std_logic;
signal \delay_measurement_inst.N_276\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_o2_6_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_o2_0_19\ : std_logic;
signal \delay_measurement_inst.start_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_256_i\ : std_logic;
signal delay_tr_input_c : std_logic;
signal delay_tr_d1 : std_logic;
signal delay_tr_d2 : std_logic;
signal \delay_measurement_inst.prev_tr_sigZ0\ : std_logic;
signal \delay_measurement_inst.tr_stateZ0Z_0\ : std_logic;
signal delay_hc_input_c : std_logic;
signal delay_hc_d1 : std_logic;
signal \delay_measurement_inst.prev_hc_sigZ0\ : std_logic;
signal \delay_measurement_inst.hc_stateZ0Z_0\ : std_logic;
signal delay_hc_d2 : std_logic;
signal clk_100mhz : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_253_i\ : std_logic;
signal \delay_measurement_inst.start_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_254_i_g\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.running_i\ : std_logic;
signal red_c_g : std_logic;
signal red_c_i : std_logic;
signal \_gnd_net_\ : std_logic;

signal reset_wire : std_logic;
signal il_min_comp2_wire : std_logic;
signal s1_phy_wire : std_logic;
signal s4_phy_wire : std_logic;
signal start_stop_wire : std_logic;
signal il_max_comp2_wire : std_logic;
signal pwm_output_wire : std_logic;
signal il_max_comp1_wire : std_logic;
signal il_min_comp1_wire : std_logic;
signal s2_phy_wire : std_logic;
signal s3_phy_wire : std_logic;
signal delay_hc_input_wire : std_logic;
signal delay_tr_input_wire : std_logic;
signal rgb_r_wire : std_logic;
signal rgb_b_wire : std_logic;
signal rgb_g_wire : std_logic;
signal \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    reset_wire <= reset;
    il_min_comp2_wire <= il_min_comp2;
    s1_phy <= s1_phy_wire;
    s4_phy <= s4_phy_wire;
    start_stop_wire <= start_stop;
    il_max_comp2_wire <= il_max_comp2;
    pwm_output <= pwm_output_wire;
    il_max_comp1_wire <= il_max_comp1;
    il_min_comp1_wire <= il_min_comp1;
    s2_phy <= s2_phy_wire;
    s3_phy <= s3_phy_wire;
    delay_hc_input_wire <= delay_hc_input;
    delay_tr_input_wire <= delay_tr_input;
    rgb_r <= rgb_r_wire;
    rgb_b <= rgb_b_wire;
    rgb_g <= rgb_g_wire;
    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__10667\,
            RESETB => \N__20181\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => clk_100mhz
        );

    \reset_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__21135\,
            GLOBALBUFFEROUTPUT => red_c_g
        );

    \reset_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21137\,
            DIN => \N__21136\,
            DOUT => \N__21135\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__21137\,
            PADOUT => \N__21136\,
            PADIN => \N__21135\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21126\,
            DIN => \N__21125\,
            DOUT => \N__21124\,
            PACKAGEPIN => il_min_comp2_wire
        );

    \il_min_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__21126\,
            PADOUT => \N__21125\,
            PADIN => \N__21124\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s1_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21117\,
            DIN => \N__21116\,
            DOUT => \N__21115\,
            PACKAGEPIN => s1_phy_wire
        );

    \s1_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__21117\,
            PADOUT => \N__21116\,
            PADIN => \N__21115\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__16859\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s4_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21108\,
            DIN => \N__21107\,
            DOUT => \N__21106\,
            PACKAGEPIN => s4_phy_wire
        );

    \s4_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__21108\,
            PADOUT => \N__21107\,
            PADIN => \N__21106\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__15671\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \start_stop_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21099\,
            DIN => \N__21098\,
            DOUT => \N__21097\,
            PACKAGEPIN => start_stop_wire
        );

    \start_stop_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__21099\,
            PADOUT => \N__21098\,
            PADIN => \N__21097\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => start_stop_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21090\,
            DIN => \N__21089\,
            DOUT => \N__21088\,
            PACKAGEPIN => il_max_comp2_wire
        );

    \il_max_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__21090\,
            PADOUT => \N__21089\,
            PADIN => \N__21088\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21081\,
            DIN => \N__21080\,
            DOUT => \N__21079\,
            PACKAGEPIN => pwm_output_wire
        );

    \pwm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__21081\,
            PADOUT => \N__21080\,
            PADIN => \N__21079\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21072\,
            DIN => \N__21071\,
            DOUT => \N__21070\,
            PACKAGEPIN => il_max_comp1_wire
        );

    \il_max_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__21072\,
            PADOUT => \N__21071\,
            PADIN => \N__21070\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21063\,
            DIN => \N__21062\,
            DOUT => \N__21061\,
            PACKAGEPIN => il_min_comp1_wire
        );

    \il_min_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__21063\,
            PADOUT => \N__21062\,
            PADIN => \N__21061\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s2_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21054\,
            DIN => \N__21053\,
            DOUT => \N__21052\,
            PACKAGEPIN => s2_phy_wire
        );

    \s2_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__21054\,
            PADOUT => \N__21053\,
            PADIN => \N__21052\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__19883\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s3_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21045\,
            DIN => \N__21044\,
            DOUT => \N__21043\,
            PACKAGEPIN => s3_phy_wire
        );

    \s3_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__21045\,
            PADOUT => \N__21044\,
            PADIN => \N__21043\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17243\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_hc_input_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21036\,
            DIN => \N__21035\,
            DOUT => \N__21034\,
            PACKAGEPIN => delay_hc_input_wire
        );

    \delay_hc_input_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__21036\,
            PADOUT => \N__21035\,
            PADIN => \N__21034\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_hc_input_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_tr_input_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21027\,
            DIN => \N__21026\,
            DOUT => \N__21025\,
            PACKAGEPIN => delay_tr_input_wire
        );

    \delay_tr_input_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__21027\,
            PADOUT => \N__21026\,
            PADIN => \N__21025\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_tr_input_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__4965\ : InMux
    port map (
            O => \N__21008\,
            I => \N__21005\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__21005\,
            I => \N__21000\
        );

    \I__4963\ : InMux
    port map (
            O => \N__21004\,
            I => \N__20997\
        );

    \I__4962\ : InMux
    port map (
            O => \N__21003\,
            I => \N__20994\
        );

    \I__4961\ : Odrv4
    port map (
            O => \N__21000\,
            I => \delay_measurement_inst.prev_hc_sigZ0\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__20997\,
            I => \delay_measurement_inst.prev_hc_sigZ0\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__20994\,
            I => \delay_measurement_inst.prev_hc_sigZ0\
        );

    \I__4958\ : InMux
    port map (
            O => \N__20987\,
            I => \N__20984\
        );

    \I__4957\ : LocalMux
    port map (
            O => \N__20984\,
            I => \N__20979\
        );

    \I__4956\ : InMux
    port map (
            O => \N__20983\,
            I => \N__20976\
        );

    \I__4955\ : InMux
    port map (
            O => \N__20982\,
            I => \N__20973\
        );

    \I__4954\ : Odrv4
    port map (
            O => \N__20979\,
            I => \delay_measurement_inst.hc_stateZ0Z_0\
        );

    \I__4953\ : LocalMux
    port map (
            O => \N__20976\,
            I => \delay_measurement_inst.hc_stateZ0Z_0\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__20973\,
            I => \delay_measurement_inst.hc_stateZ0Z_0\
        );

    \I__4951\ : InMux
    port map (
            O => \N__20966\,
            I => \N__20959\
        );

    \I__4950\ : InMux
    port map (
            O => \N__20965\,
            I => \N__20959\
        );

    \I__4949\ : InMux
    port map (
            O => \N__20964\,
            I => \N__20956\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__20959\,
            I => \N__20950\
        );

    \I__4947\ : LocalMux
    port map (
            O => \N__20956\,
            I => \N__20950\
        );

    \I__4946\ : InMux
    port map (
            O => \N__20955\,
            I => \N__20947\
        );

    \I__4945\ : Odrv4
    port map (
            O => \N__20950\,
            I => delay_hc_d2
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__20947\,
            I => delay_hc_d2
        );

    \I__4943\ : ClkMux
    port map (
            O => \N__20942\,
            I => \N__20705\
        );

    \I__4942\ : ClkMux
    port map (
            O => \N__20941\,
            I => \N__20705\
        );

    \I__4941\ : ClkMux
    port map (
            O => \N__20940\,
            I => \N__20705\
        );

    \I__4940\ : ClkMux
    port map (
            O => \N__20939\,
            I => \N__20705\
        );

    \I__4939\ : ClkMux
    port map (
            O => \N__20938\,
            I => \N__20705\
        );

    \I__4938\ : ClkMux
    port map (
            O => \N__20937\,
            I => \N__20705\
        );

    \I__4937\ : ClkMux
    port map (
            O => \N__20936\,
            I => \N__20705\
        );

    \I__4936\ : ClkMux
    port map (
            O => \N__20935\,
            I => \N__20705\
        );

    \I__4935\ : ClkMux
    port map (
            O => \N__20934\,
            I => \N__20705\
        );

    \I__4934\ : ClkMux
    port map (
            O => \N__20933\,
            I => \N__20705\
        );

    \I__4933\ : ClkMux
    port map (
            O => \N__20932\,
            I => \N__20705\
        );

    \I__4932\ : ClkMux
    port map (
            O => \N__20931\,
            I => \N__20705\
        );

    \I__4931\ : ClkMux
    port map (
            O => \N__20930\,
            I => \N__20705\
        );

    \I__4930\ : ClkMux
    port map (
            O => \N__20929\,
            I => \N__20705\
        );

    \I__4929\ : ClkMux
    port map (
            O => \N__20928\,
            I => \N__20705\
        );

    \I__4928\ : ClkMux
    port map (
            O => \N__20927\,
            I => \N__20705\
        );

    \I__4927\ : ClkMux
    port map (
            O => \N__20926\,
            I => \N__20705\
        );

    \I__4926\ : ClkMux
    port map (
            O => \N__20925\,
            I => \N__20705\
        );

    \I__4925\ : ClkMux
    port map (
            O => \N__20924\,
            I => \N__20705\
        );

    \I__4924\ : ClkMux
    port map (
            O => \N__20923\,
            I => \N__20705\
        );

    \I__4923\ : ClkMux
    port map (
            O => \N__20922\,
            I => \N__20705\
        );

    \I__4922\ : ClkMux
    port map (
            O => \N__20921\,
            I => \N__20705\
        );

    \I__4921\ : ClkMux
    port map (
            O => \N__20920\,
            I => \N__20705\
        );

    \I__4920\ : ClkMux
    port map (
            O => \N__20919\,
            I => \N__20705\
        );

    \I__4919\ : ClkMux
    port map (
            O => \N__20918\,
            I => \N__20705\
        );

    \I__4918\ : ClkMux
    port map (
            O => \N__20917\,
            I => \N__20705\
        );

    \I__4917\ : ClkMux
    port map (
            O => \N__20916\,
            I => \N__20705\
        );

    \I__4916\ : ClkMux
    port map (
            O => \N__20915\,
            I => \N__20705\
        );

    \I__4915\ : ClkMux
    port map (
            O => \N__20914\,
            I => \N__20705\
        );

    \I__4914\ : ClkMux
    port map (
            O => \N__20913\,
            I => \N__20705\
        );

    \I__4913\ : ClkMux
    port map (
            O => \N__20912\,
            I => \N__20705\
        );

    \I__4912\ : ClkMux
    port map (
            O => \N__20911\,
            I => \N__20705\
        );

    \I__4911\ : ClkMux
    port map (
            O => \N__20910\,
            I => \N__20705\
        );

    \I__4910\ : ClkMux
    port map (
            O => \N__20909\,
            I => \N__20705\
        );

    \I__4909\ : ClkMux
    port map (
            O => \N__20908\,
            I => \N__20705\
        );

    \I__4908\ : ClkMux
    port map (
            O => \N__20907\,
            I => \N__20705\
        );

    \I__4907\ : ClkMux
    port map (
            O => \N__20906\,
            I => \N__20705\
        );

    \I__4906\ : ClkMux
    port map (
            O => \N__20905\,
            I => \N__20705\
        );

    \I__4905\ : ClkMux
    port map (
            O => \N__20904\,
            I => \N__20705\
        );

    \I__4904\ : ClkMux
    port map (
            O => \N__20903\,
            I => \N__20705\
        );

    \I__4903\ : ClkMux
    port map (
            O => \N__20902\,
            I => \N__20705\
        );

    \I__4902\ : ClkMux
    port map (
            O => \N__20901\,
            I => \N__20705\
        );

    \I__4901\ : ClkMux
    port map (
            O => \N__20900\,
            I => \N__20705\
        );

    \I__4900\ : ClkMux
    port map (
            O => \N__20899\,
            I => \N__20705\
        );

    \I__4899\ : ClkMux
    port map (
            O => \N__20898\,
            I => \N__20705\
        );

    \I__4898\ : ClkMux
    port map (
            O => \N__20897\,
            I => \N__20705\
        );

    \I__4897\ : ClkMux
    port map (
            O => \N__20896\,
            I => \N__20705\
        );

    \I__4896\ : ClkMux
    port map (
            O => \N__20895\,
            I => \N__20705\
        );

    \I__4895\ : ClkMux
    port map (
            O => \N__20894\,
            I => \N__20705\
        );

    \I__4894\ : ClkMux
    port map (
            O => \N__20893\,
            I => \N__20705\
        );

    \I__4893\ : ClkMux
    port map (
            O => \N__20892\,
            I => \N__20705\
        );

    \I__4892\ : ClkMux
    port map (
            O => \N__20891\,
            I => \N__20705\
        );

    \I__4891\ : ClkMux
    port map (
            O => \N__20890\,
            I => \N__20705\
        );

    \I__4890\ : ClkMux
    port map (
            O => \N__20889\,
            I => \N__20705\
        );

    \I__4889\ : ClkMux
    port map (
            O => \N__20888\,
            I => \N__20705\
        );

    \I__4888\ : ClkMux
    port map (
            O => \N__20887\,
            I => \N__20705\
        );

    \I__4887\ : ClkMux
    port map (
            O => \N__20886\,
            I => \N__20705\
        );

    \I__4886\ : ClkMux
    port map (
            O => \N__20885\,
            I => \N__20705\
        );

    \I__4885\ : ClkMux
    port map (
            O => \N__20884\,
            I => \N__20705\
        );

    \I__4884\ : ClkMux
    port map (
            O => \N__20883\,
            I => \N__20705\
        );

    \I__4883\ : ClkMux
    port map (
            O => \N__20882\,
            I => \N__20705\
        );

    \I__4882\ : ClkMux
    port map (
            O => \N__20881\,
            I => \N__20705\
        );

    \I__4881\ : ClkMux
    port map (
            O => \N__20880\,
            I => \N__20705\
        );

    \I__4880\ : ClkMux
    port map (
            O => \N__20879\,
            I => \N__20705\
        );

    \I__4879\ : ClkMux
    port map (
            O => \N__20878\,
            I => \N__20705\
        );

    \I__4878\ : ClkMux
    port map (
            O => \N__20877\,
            I => \N__20705\
        );

    \I__4877\ : ClkMux
    port map (
            O => \N__20876\,
            I => \N__20705\
        );

    \I__4876\ : ClkMux
    port map (
            O => \N__20875\,
            I => \N__20705\
        );

    \I__4875\ : ClkMux
    port map (
            O => \N__20874\,
            I => \N__20705\
        );

    \I__4874\ : ClkMux
    port map (
            O => \N__20873\,
            I => \N__20705\
        );

    \I__4873\ : ClkMux
    port map (
            O => \N__20872\,
            I => \N__20705\
        );

    \I__4872\ : ClkMux
    port map (
            O => \N__20871\,
            I => \N__20705\
        );

    \I__4871\ : ClkMux
    port map (
            O => \N__20870\,
            I => \N__20705\
        );

    \I__4870\ : ClkMux
    port map (
            O => \N__20869\,
            I => \N__20705\
        );

    \I__4869\ : ClkMux
    port map (
            O => \N__20868\,
            I => \N__20705\
        );

    \I__4868\ : ClkMux
    port map (
            O => \N__20867\,
            I => \N__20705\
        );

    \I__4867\ : ClkMux
    port map (
            O => \N__20866\,
            I => \N__20705\
        );

    \I__4866\ : ClkMux
    port map (
            O => \N__20865\,
            I => \N__20705\
        );

    \I__4865\ : ClkMux
    port map (
            O => \N__20864\,
            I => \N__20705\
        );

    \I__4864\ : GlobalMux
    port map (
            O => \N__20705\,
            I => clk_100mhz
        );

    \I__4863\ : IoInMux
    port map (
            O => \N__20702\,
            I => \N__20699\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__20699\,
            I => \N__20696\
        );

    \I__4861\ : Odrv12
    port map (
            O => \N__20696\,
            I => \delay_measurement_inst.delay_hc_timer.N_253_i\
        );

    \I__4860\ : InMux
    port map (
            O => \N__20693\,
            I => \N__20689\
        );

    \I__4859\ : InMux
    port map (
            O => \N__20692\,
            I => \N__20686\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__20689\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__20686\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__4856\ : InMux
    port map (
            O => \N__20681\,
            I => \N__20674\
        );

    \I__4855\ : InMux
    port map (
            O => \N__20680\,
            I => \N__20674\
        );

    \I__4854\ : InMux
    port map (
            O => \N__20679\,
            I => \N__20671\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__20674\,
            I => \N__20668\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__20671\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__4851\ : Odrv4
    port map (
            O => \N__20668\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__4850\ : CEMux
    port map (
            O => \N__20663\,
            I => \N__20660\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__20660\,
            I => \N__20655\
        );

    \I__4848\ : CEMux
    port map (
            O => \N__20659\,
            I => \N__20652\
        );

    \I__4847\ : CEMux
    port map (
            O => \N__20658\,
            I => \N__20648\
        );

    \I__4846\ : Span4Mux_v
    port map (
            O => \N__20655\,
            I => \N__20643\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__20652\,
            I => \N__20643\
        );

    \I__4844\ : CEMux
    port map (
            O => \N__20651\,
            I => \N__20640\
        );

    \I__4843\ : LocalMux
    port map (
            O => \N__20648\,
            I => \N__20637\
        );

    \I__4842\ : Span4Mux_h
    port map (
            O => \N__20643\,
            I => \N__20634\
        );

    \I__4841\ : LocalMux
    port map (
            O => \N__20640\,
            I => \N__20631\
        );

    \I__4840\ : Span4Mux_v
    port map (
            O => \N__20637\,
            I => \N__20628\
        );

    \I__4839\ : Span4Mux_h
    port map (
            O => \N__20634\,
            I => \N__20625\
        );

    \I__4838\ : Sp12to4
    port map (
            O => \N__20631\,
            I => \N__20622\
        );

    \I__4837\ : Odrv4
    port map (
            O => \N__20628\,
            I => \delay_measurement_inst.delay_hc_timer.N_254_i_g\
        );

    \I__4836\ : Odrv4
    port map (
            O => \N__20625\,
            I => \delay_measurement_inst.delay_hc_timer.N_254_i_g\
        );

    \I__4835\ : Odrv12
    port map (
            O => \N__20622\,
            I => \delay_measurement_inst.delay_hc_timer.N_254_i_g\
        );

    \I__4834\ : InMux
    port map (
            O => \N__20615\,
            I => \N__20609\
        );

    \I__4833\ : InMux
    port map (
            O => \N__20614\,
            I => \N__20602\
        );

    \I__4832\ : InMux
    port map (
            O => \N__20613\,
            I => \N__20602\
        );

    \I__4831\ : InMux
    port map (
            O => \N__20612\,
            I => \N__20602\
        );

    \I__4830\ : LocalMux
    port map (
            O => \N__20609\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__4829\ : LocalMux
    port map (
            O => \N__20602\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__4828\ : InMux
    port map (
            O => \N__20597\,
            I => \N__20569\
        );

    \I__4827\ : InMux
    port map (
            O => \N__20596\,
            I => \N__20569\
        );

    \I__4826\ : InMux
    port map (
            O => \N__20595\,
            I => \N__20569\
        );

    \I__4825\ : InMux
    port map (
            O => \N__20594\,
            I => \N__20569\
        );

    \I__4824\ : InMux
    port map (
            O => \N__20593\,
            I => \N__20560\
        );

    \I__4823\ : InMux
    port map (
            O => \N__20592\,
            I => \N__20560\
        );

    \I__4822\ : InMux
    port map (
            O => \N__20591\,
            I => \N__20560\
        );

    \I__4821\ : InMux
    port map (
            O => \N__20590\,
            I => \N__20560\
        );

    \I__4820\ : InMux
    port map (
            O => \N__20589\,
            I => \N__20551\
        );

    \I__4819\ : InMux
    port map (
            O => \N__20588\,
            I => \N__20551\
        );

    \I__4818\ : InMux
    port map (
            O => \N__20587\,
            I => \N__20551\
        );

    \I__4817\ : InMux
    port map (
            O => \N__20586\,
            I => \N__20551\
        );

    \I__4816\ : InMux
    port map (
            O => \N__20585\,
            I => \N__20542\
        );

    \I__4815\ : InMux
    port map (
            O => \N__20584\,
            I => \N__20542\
        );

    \I__4814\ : InMux
    port map (
            O => \N__20583\,
            I => \N__20542\
        );

    \I__4813\ : InMux
    port map (
            O => \N__20582\,
            I => \N__20542\
        );

    \I__4812\ : InMux
    port map (
            O => \N__20581\,
            I => \N__20533\
        );

    \I__4811\ : InMux
    port map (
            O => \N__20580\,
            I => \N__20533\
        );

    \I__4810\ : InMux
    port map (
            O => \N__20579\,
            I => \N__20533\
        );

    \I__4809\ : InMux
    port map (
            O => \N__20578\,
            I => \N__20533\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__20569\,
            I => \N__20518\
        );

    \I__4807\ : LocalMux
    port map (
            O => \N__20560\,
            I => \N__20518\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__20551\,
            I => \N__20511\
        );

    \I__4805\ : LocalMux
    port map (
            O => \N__20542\,
            I => \N__20511\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__20533\,
            I => \N__20511\
        );

    \I__4803\ : InMux
    port map (
            O => \N__20532\,
            I => \N__20506\
        );

    \I__4802\ : InMux
    port map (
            O => \N__20531\,
            I => \N__20506\
        );

    \I__4801\ : InMux
    port map (
            O => \N__20530\,
            I => \N__20497\
        );

    \I__4800\ : InMux
    port map (
            O => \N__20529\,
            I => \N__20497\
        );

    \I__4799\ : InMux
    port map (
            O => \N__20528\,
            I => \N__20497\
        );

    \I__4798\ : InMux
    port map (
            O => \N__20527\,
            I => \N__20497\
        );

    \I__4797\ : InMux
    port map (
            O => \N__20526\,
            I => \N__20488\
        );

    \I__4796\ : InMux
    port map (
            O => \N__20525\,
            I => \N__20488\
        );

    \I__4795\ : InMux
    port map (
            O => \N__20524\,
            I => \N__20488\
        );

    \I__4794\ : InMux
    port map (
            O => \N__20523\,
            I => \N__20488\
        );

    \I__4793\ : Span4Mux_v
    port map (
            O => \N__20518\,
            I => \N__20479\
        );

    \I__4792\ : Span4Mux_v
    port map (
            O => \N__20511\,
            I => \N__20479\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__20506\,
            I => \N__20479\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__20497\,
            I => \N__20479\
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__20488\,
            I => \N__20476\
        );

    \I__4788\ : Span4Mux_h
    port map (
            O => \N__20479\,
            I => \N__20473\
        );

    \I__4787\ : Odrv12
    port map (
            O => \N__20476\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__4786\ : Odrv4
    port map (
            O => \N__20473\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__4785\ : CascadeMux
    port map (
            O => \N__20468\,
            I => \N__20458\
        );

    \I__4784\ : CascadeMux
    port map (
            O => \N__20467\,
            I => \N__20455\
        );

    \I__4783\ : InMux
    port map (
            O => \N__20466\,
            I => \N__20452\
        );

    \I__4782\ : InMux
    port map (
            O => \N__20465\,
            I => \N__20447\
        );

    \I__4781\ : InMux
    port map (
            O => \N__20464\,
            I => \N__20447\
        );

    \I__4780\ : InMux
    port map (
            O => \N__20463\,
            I => \N__20444\
        );

    \I__4779\ : InMux
    port map (
            O => \N__20462\,
            I => \N__20441\
        );

    \I__4778\ : InMux
    port map (
            O => \N__20461\,
            I => \N__20438\
        );

    \I__4777\ : InMux
    port map (
            O => \N__20458\,
            I => \N__20435\
        );

    \I__4776\ : InMux
    port map (
            O => \N__20455\,
            I => \N__20432\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__20452\,
            I => \N__20429\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__20447\,
            I => \N__20426\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__20444\,
            I => \N__20402\
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__20441\,
            I => \N__20386\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__20438\,
            I => \N__20363\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__20435\,
            I => \N__20357\
        );

    \I__4769\ : LocalMux
    port map (
            O => \N__20432\,
            I => \N__20347\
        );

    \I__4768\ : Glb2LocalMux
    port map (
            O => \N__20429\,
            I => \N__20201\
        );

    \I__4767\ : Glb2LocalMux
    port map (
            O => \N__20426\,
            I => \N__20201\
        );

    \I__4766\ : SRMux
    port map (
            O => \N__20425\,
            I => \N__20201\
        );

    \I__4765\ : SRMux
    port map (
            O => \N__20424\,
            I => \N__20201\
        );

    \I__4764\ : SRMux
    port map (
            O => \N__20423\,
            I => \N__20201\
        );

    \I__4763\ : SRMux
    port map (
            O => \N__20422\,
            I => \N__20201\
        );

    \I__4762\ : SRMux
    port map (
            O => \N__20421\,
            I => \N__20201\
        );

    \I__4761\ : SRMux
    port map (
            O => \N__20420\,
            I => \N__20201\
        );

    \I__4760\ : SRMux
    port map (
            O => \N__20419\,
            I => \N__20201\
        );

    \I__4759\ : SRMux
    port map (
            O => \N__20418\,
            I => \N__20201\
        );

    \I__4758\ : SRMux
    port map (
            O => \N__20417\,
            I => \N__20201\
        );

    \I__4757\ : SRMux
    port map (
            O => \N__20416\,
            I => \N__20201\
        );

    \I__4756\ : SRMux
    port map (
            O => \N__20415\,
            I => \N__20201\
        );

    \I__4755\ : SRMux
    port map (
            O => \N__20414\,
            I => \N__20201\
        );

    \I__4754\ : SRMux
    port map (
            O => \N__20413\,
            I => \N__20201\
        );

    \I__4753\ : SRMux
    port map (
            O => \N__20412\,
            I => \N__20201\
        );

    \I__4752\ : SRMux
    port map (
            O => \N__20411\,
            I => \N__20201\
        );

    \I__4751\ : SRMux
    port map (
            O => \N__20410\,
            I => \N__20201\
        );

    \I__4750\ : SRMux
    port map (
            O => \N__20409\,
            I => \N__20201\
        );

    \I__4749\ : SRMux
    port map (
            O => \N__20408\,
            I => \N__20201\
        );

    \I__4748\ : SRMux
    port map (
            O => \N__20407\,
            I => \N__20201\
        );

    \I__4747\ : SRMux
    port map (
            O => \N__20406\,
            I => \N__20201\
        );

    \I__4746\ : SRMux
    port map (
            O => \N__20405\,
            I => \N__20201\
        );

    \I__4745\ : Glb2LocalMux
    port map (
            O => \N__20402\,
            I => \N__20201\
        );

    \I__4744\ : SRMux
    port map (
            O => \N__20401\,
            I => \N__20201\
        );

    \I__4743\ : SRMux
    port map (
            O => \N__20400\,
            I => \N__20201\
        );

    \I__4742\ : SRMux
    port map (
            O => \N__20399\,
            I => \N__20201\
        );

    \I__4741\ : SRMux
    port map (
            O => \N__20398\,
            I => \N__20201\
        );

    \I__4740\ : SRMux
    port map (
            O => \N__20397\,
            I => \N__20201\
        );

    \I__4739\ : SRMux
    port map (
            O => \N__20396\,
            I => \N__20201\
        );

    \I__4738\ : SRMux
    port map (
            O => \N__20395\,
            I => \N__20201\
        );

    \I__4737\ : SRMux
    port map (
            O => \N__20394\,
            I => \N__20201\
        );

    \I__4736\ : SRMux
    port map (
            O => \N__20393\,
            I => \N__20201\
        );

    \I__4735\ : SRMux
    port map (
            O => \N__20392\,
            I => \N__20201\
        );

    \I__4734\ : SRMux
    port map (
            O => \N__20391\,
            I => \N__20201\
        );

    \I__4733\ : SRMux
    port map (
            O => \N__20390\,
            I => \N__20201\
        );

    \I__4732\ : SRMux
    port map (
            O => \N__20389\,
            I => \N__20201\
        );

    \I__4731\ : Glb2LocalMux
    port map (
            O => \N__20386\,
            I => \N__20201\
        );

    \I__4730\ : SRMux
    port map (
            O => \N__20385\,
            I => \N__20201\
        );

    \I__4729\ : SRMux
    port map (
            O => \N__20384\,
            I => \N__20201\
        );

    \I__4728\ : SRMux
    port map (
            O => \N__20383\,
            I => \N__20201\
        );

    \I__4727\ : SRMux
    port map (
            O => \N__20382\,
            I => \N__20201\
        );

    \I__4726\ : SRMux
    port map (
            O => \N__20381\,
            I => \N__20201\
        );

    \I__4725\ : SRMux
    port map (
            O => \N__20380\,
            I => \N__20201\
        );

    \I__4724\ : SRMux
    port map (
            O => \N__20379\,
            I => \N__20201\
        );

    \I__4723\ : SRMux
    port map (
            O => \N__20378\,
            I => \N__20201\
        );

    \I__4722\ : SRMux
    port map (
            O => \N__20377\,
            I => \N__20201\
        );

    \I__4721\ : SRMux
    port map (
            O => \N__20376\,
            I => \N__20201\
        );

    \I__4720\ : SRMux
    port map (
            O => \N__20375\,
            I => \N__20201\
        );

    \I__4719\ : SRMux
    port map (
            O => \N__20374\,
            I => \N__20201\
        );

    \I__4718\ : SRMux
    port map (
            O => \N__20373\,
            I => \N__20201\
        );

    \I__4717\ : SRMux
    port map (
            O => \N__20372\,
            I => \N__20201\
        );

    \I__4716\ : SRMux
    port map (
            O => \N__20371\,
            I => \N__20201\
        );

    \I__4715\ : SRMux
    port map (
            O => \N__20370\,
            I => \N__20201\
        );

    \I__4714\ : SRMux
    port map (
            O => \N__20369\,
            I => \N__20201\
        );

    \I__4713\ : SRMux
    port map (
            O => \N__20368\,
            I => \N__20201\
        );

    \I__4712\ : SRMux
    port map (
            O => \N__20367\,
            I => \N__20201\
        );

    \I__4711\ : SRMux
    port map (
            O => \N__20366\,
            I => \N__20201\
        );

    \I__4710\ : Glb2LocalMux
    port map (
            O => \N__20363\,
            I => \N__20201\
        );

    \I__4709\ : SRMux
    port map (
            O => \N__20362\,
            I => \N__20201\
        );

    \I__4708\ : SRMux
    port map (
            O => \N__20361\,
            I => \N__20201\
        );

    \I__4707\ : SRMux
    port map (
            O => \N__20360\,
            I => \N__20201\
        );

    \I__4706\ : Glb2LocalMux
    port map (
            O => \N__20357\,
            I => \N__20201\
        );

    \I__4705\ : SRMux
    port map (
            O => \N__20356\,
            I => \N__20201\
        );

    \I__4704\ : SRMux
    port map (
            O => \N__20355\,
            I => \N__20201\
        );

    \I__4703\ : SRMux
    port map (
            O => \N__20354\,
            I => \N__20201\
        );

    \I__4702\ : SRMux
    port map (
            O => \N__20353\,
            I => \N__20201\
        );

    \I__4701\ : SRMux
    port map (
            O => \N__20352\,
            I => \N__20201\
        );

    \I__4700\ : SRMux
    port map (
            O => \N__20351\,
            I => \N__20201\
        );

    \I__4699\ : SRMux
    port map (
            O => \N__20350\,
            I => \N__20201\
        );

    \I__4698\ : Glb2LocalMux
    port map (
            O => \N__20347\,
            I => \N__20201\
        );

    \I__4697\ : SRMux
    port map (
            O => \N__20346\,
            I => \N__20201\
        );

    \I__4696\ : GlobalMux
    port map (
            O => \N__20201\,
            I => \N__20198\
        );

    \I__4695\ : gio2CtrlBuf
    port map (
            O => \N__20198\,
            I => red_c_g
        );

    \I__4694\ : CEMux
    port map (
            O => \N__20195\,
            I => \N__20192\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__20192\,
            I => \N__20185\
        );

    \I__4692\ : CEMux
    port map (
            O => \N__20191\,
            I => \N__20182\
        );

    \I__4691\ : CEMux
    port map (
            O => \N__20190\,
            I => \N__20178\
        );

    \I__4690\ : CEMux
    port map (
            O => \N__20189\,
            I => \N__20175\
        );

    \I__4689\ : CEMux
    port map (
            O => \N__20188\,
            I => \N__20172\
        );

    \I__4688\ : Span4Mux_v
    port map (
            O => \N__20185\,
            I => \N__20168\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__20182\,
            I => \N__20165\
        );

    \I__4686\ : IoInMux
    port map (
            O => \N__20181\,
            I => \N__20162\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__20178\,
            I => \N__20159\
        );

    \I__4684\ : LocalMux
    port map (
            O => \N__20175\,
            I => \N__20156\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__20172\,
            I => \N__20153\
        );

    \I__4682\ : CEMux
    port map (
            O => \N__20171\,
            I => \N__20150\
        );

    \I__4681\ : Span4Mux_v
    port map (
            O => \N__20168\,
            I => \N__20147\
        );

    \I__4680\ : Span4Mux_h
    port map (
            O => \N__20165\,
            I => \N__20144\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__20162\,
            I => \N__20141\
        );

    \I__4678\ : Span4Mux_h
    port map (
            O => \N__20159\,
            I => \N__20136\
        );

    \I__4677\ : Span4Mux_h
    port map (
            O => \N__20156\,
            I => \N__20136\
        );

    \I__4676\ : Span4Mux_v
    port map (
            O => \N__20153\,
            I => \N__20131\
        );

    \I__4675\ : LocalMux
    port map (
            O => \N__20150\,
            I => \N__20131\
        );

    \I__4674\ : Span4Mux_h
    port map (
            O => \N__20147\,
            I => \N__20128\
        );

    \I__4673\ : Span4Mux_h
    port map (
            O => \N__20144\,
            I => \N__20125\
        );

    \I__4672\ : IoSpan4Mux
    port map (
            O => \N__20141\,
            I => \N__20122\
        );

    \I__4671\ : Span4Mux_h
    port map (
            O => \N__20136\,
            I => \N__20117\
        );

    \I__4670\ : Span4Mux_v
    port map (
            O => \N__20131\,
            I => \N__20117\
        );

    \I__4669\ : Span4Mux_h
    port map (
            O => \N__20128\,
            I => \N__20114\
        );

    \I__4668\ : Span4Mux_h
    port map (
            O => \N__20125\,
            I => \N__20107\
        );

    \I__4667\ : Span4Mux_s2_v
    port map (
            O => \N__20122\,
            I => \N__20107\
        );

    \I__4666\ : Span4Mux_v
    port map (
            O => \N__20117\,
            I => \N__20107\
        );

    \I__4665\ : Odrv4
    port map (
            O => \N__20114\,
            I => red_c_i
        );

    \I__4664\ : Odrv4
    port map (
            O => \N__20107\,
            I => red_c_i
        );

    \I__4663\ : InMux
    port map (
            O => \N__20102\,
            I => \N__20098\
        );

    \I__4662\ : InMux
    port map (
            O => \N__20101\,
            I => \N__20095\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__20098\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__20095\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__4659\ : InMux
    port map (
            O => \N__20090\,
            I => \N__20085\
        );

    \I__4658\ : InMux
    port map (
            O => \N__20089\,
            I => \N__20082\
        );

    \I__4657\ : InMux
    port map (
            O => \N__20088\,
            I => \N__20079\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__20085\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__4655\ : LocalMux
    port map (
            O => \N__20082\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__20079\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__4653\ : InMux
    port map (
            O => \N__20072\,
            I => \N__20066\
        );

    \I__4652\ : InMux
    port map (
            O => \N__20071\,
            I => \N__20063\
        );

    \I__4651\ : InMux
    port map (
            O => \N__20070\,
            I => \N__20060\
        );

    \I__4650\ : InMux
    port map (
            O => \N__20069\,
            I => \N__20057\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__20066\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__20063\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__20060\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__20057\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__4645\ : IoInMux
    port map (
            O => \N__20048\,
            I => \N__20045\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__20045\,
            I => \N__20042\
        );

    \I__4643\ : Span12Mux_s5_v
    port map (
            O => \N__20042\,
            I => \N__20039\
        );

    \I__4642\ : Odrv12
    port map (
            O => \N__20039\,
            I => \delay_measurement_inst.delay_tr_timer.N_256_i\
        );

    \I__4641\ : InMux
    port map (
            O => \N__20036\,
            I => \N__20033\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__20033\,
            I => \N__20030\
        );

    \I__4639\ : Span4Mux_v
    port map (
            O => \N__20030\,
            I => \N__20027\
        );

    \I__4638\ : Sp12to4
    port map (
            O => \N__20027\,
            I => \N__20024\
        );

    \I__4637\ : Span12Mux_s10_h
    port map (
            O => \N__20024\,
            I => \N__20021\
        );

    \I__4636\ : Odrv12
    port map (
            O => \N__20021\,
            I => delay_tr_input_c
        );

    \I__4635\ : InMux
    port map (
            O => \N__20018\,
            I => \N__20015\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__20015\,
            I => delay_tr_d1
        );

    \I__4633\ : InMux
    port map (
            O => \N__20012\,
            I => \N__20006\
        );

    \I__4632\ : InMux
    port map (
            O => \N__20011\,
            I => \N__20003\
        );

    \I__4631\ : InMux
    port map (
            O => \N__20010\,
            I => \N__19998\
        );

    \I__4630\ : InMux
    port map (
            O => \N__20009\,
            I => \N__19998\
        );

    \I__4629\ : LocalMux
    port map (
            O => \N__20006\,
            I => delay_tr_d2
        );

    \I__4628\ : LocalMux
    port map (
            O => \N__20003\,
            I => delay_tr_d2
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__19998\,
            I => delay_tr_d2
        );

    \I__4626\ : InMux
    port map (
            O => \N__19991\,
            I => \N__19986\
        );

    \I__4625\ : InMux
    port map (
            O => \N__19990\,
            I => \N__19983\
        );

    \I__4624\ : InMux
    port map (
            O => \N__19989\,
            I => \N__19980\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__19986\,
            I => \delay_measurement_inst.prev_tr_sigZ0\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__19983\,
            I => \delay_measurement_inst.prev_tr_sigZ0\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__19980\,
            I => \delay_measurement_inst.prev_tr_sigZ0\
        );

    \I__4620\ : InMux
    port map (
            O => \N__19973\,
            I => \N__19968\
        );

    \I__4619\ : InMux
    port map (
            O => \N__19972\,
            I => \N__19965\
        );

    \I__4618\ : InMux
    port map (
            O => \N__19971\,
            I => \N__19962\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__19968\,
            I => \delay_measurement_inst.tr_stateZ0Z_0\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__19965\,
            I => \delay_measurement_inst.tr_stateZ0Z_0\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__19962\,
            I => \delay_measurement_inst.tr_stateZ0Z_0\
        );

    \I__4614\ : InMux
    port map (
            O => \N__19955\,
            I => \N__19952\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__19952\,
            I => \N__19949\
        );

    \I__4612\ : Span12Mux_h
    port map (
            O => \N__19949\,
            I => \N__19946\
        );

    \I__4611\ : Span12Mux_v
    port map (
            O => \N__19946\,
            I => \N__19943\
        );

    \I__4610\ : Odrv12
    port map (
            O => \N__19943\,
            I => delay_hc_input_c
        );

    \I__4609\ : InMux
    port map (
            O => \N__19940\,
            I => \N__19937\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__19937\,
            I => delay_hc_d1
        );

    \I__4607\ : IoInMux
    port map (
            O => \N__19934\,
            I => \N__19931\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__19931\,
            I => \N__19928\
        );

    \I__4605\ : Span12Mux_s4_v
    port map (
            O => \N__19928\,
            I => \N__19925\
        );

    \I__4604\ : Span12Mux_v
    port map (
            O => \N__19925\,
            I => \N__19922\
        );

    \I__4603\ : Odrv12
    port map (
            O => \N__19922\,
            I => \delay_measurement_inst.delay_tr_timer.N_255_i\
        );

    \I__4602\ : InMux
    port map (
            O => \N__19919\,
            I => \N__19916\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__19916\,
            I => \N__19911\
        );

    \I__4600\ : CascadeMux
    port map (
            O => \N__19915\,
            I => \N__19907\
        );

    \I__4599\ : CascadeMux
    port map (
            O => \N__19914\,
            I => \N__19904\
        );

    \I__4598\ : Span4Mux_h
    port map (
            O => \N__19911\,
            I => \N__19901\
        );

    \I__4597\ : InMux
    port map (
            O => \N__19910\,
            I => \N__19898\
        );

    \I__4596\ : InMux
    port map (
            O => \N__19907\,
            I => \N__19893\
        );

    \I__4595\ : InMux
    port map (
            O => \N__19904\,
            I => \N__19893\
        );

    \I__4594\ : Span4Mux_v
    port map (
            O => \N__19901\,
            I => \N__19888\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__19898\,
            I => \N__19888\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__19893\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__4591\ : Odrv4
    port map (
            O => \N__19888\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__4590\ : IoInMux
    port map (
            O => \N__19883\,
            I => \N__19880\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__19880\,
            I => \N__19877\
        );

    \I__4588\ : Span4Mux_s3_v
    port map (
            O => \N__19877\,
            I => \N__19874\
        );

    \I__4587\ : Span4Mux_v
    port map (
            O => \N__19874\,
            I => \N__19871\
        );

    \I__4586\ : Span4Mux_v
    port map (
            O => \N__19871\,
            I => \N__19868\
        );

    \I__4585\ : Odrv4
    port map (
            O => \N__19868\,
            I => s2_phy_c
        );

    \I__4584\ : InMux
    port map (
            O => \N__19865\,
            I => \N__19862\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__19862\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__4582\ : InMux
    port map (
            O => \N__19859\,
            I => \N__19856\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__19856\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__4580\ : CascadeMux
    port map (
            O => \N__19853\,
            I => \N__19850\
        );

    \I__4579\ : InMux
    port map (
            O => \N__19850\,
            I => \N__19847\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__19847\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__4577\ : InMux
    port map (
            O => \N__19844\,
            I => \N__19841\
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__19841\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__4575\ : InMux
    port map (
            O => \N__19838\,
            I => \N__19835\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__19835\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__4573\ : CascadeMux
    port map (
            O => \N__19832\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_o2_7_19_cascade_\
        );

    \I__4572\ : InMux
    port map (
            O => \N__19829\,
            I => \N__19810\
        );

    \I__4571\ : InMux
    port map (
            O => \N__19828\,
            I => \N__19810\
        );

    \I__4570\ : InMux
    port map (
            O => \N__19827\,
            I => \N__19810\
        );

    \I__4569\ : InMux
    port map (
            O => \N__19826\,
            I => \N__19810\
        );

    \I__4568\ : InMux
    port map (
            O => \N__19825\,
            I => \N__19810\
        );

    \I__4567\ : InMux
    port map (
            O => \N__19824\,
            I => \N__19801\
        );

    \I__4566\ : InMux
    port map (
            O => \N__19823\,
            I => \N__19801\
        );

    \I__4565\ : InMux
    port map (
            O => \N__19822\,
            I => \N__19801\
        );

    \I__4564\ : InMux
    port map (
            O => \N__19821\,
            I => \N__19801\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__19810\,
            I => \N__19798\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__19801\,
            I => \N__19795\
        );

    \I__4561\ : Odrv12
    port map (
            O => \N__19798\,
            I => \delay_measurement_inst.N_276\
        );

    \I__4560\ : Odrv4
    port map (
            O => \N__19795\,
            I => \delay_measurement_inst.N_276\
        );

    \I__4559\ : InMux
    port map (
            O => \N__19790\,
            I => \N__19787\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__19787\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__4557\ : InMux
    port map (
            O => \N__19784\,
            I => \N__19781\
        );

    \I__4556\ : LocalMux
    port map (
            O => \N__19781\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__4555\ : CascadeMux
    port map (
            O => \N__19778\,
            I => \N__19775\
        );

    \I__4554\ : InMux
    port map (
            O => \N__19775\,
            I => \N__19772\
        );

    \I__4553\ : LocalMux
    port map (
            O => \N__19772\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__4552\ : InMux
    port map (
            O => \N__19769\,
            I => \N__19766\
        );

    \I__4551\ : LocalMux
    port map (
            O => \N__19766\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__4550\ : InMux
    port map (
            O => \N__19763\,
            I => \N__19760\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__19760\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_o2_6_19\
        );

    \I__4548\ : InMux
    port map (
            O => \N__19757\,
            I => \N__19754\
        );

    \I__4547\ : LocalMux
    port map (
            O => \N__19754\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_30\
        );

    \I__4546\ : InMux
    port map (
            O => \N__19751\,
            I => \N__19748\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__19748\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__4544\ : InMux
    port map (
            O => \N__19745\,
            I => \N__19742\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__19742\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_o2_0_19\
        );

    \I__4542\ : InMux
    port map (
            O => \N__19739\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__4541\ : CascadeMux
    port map (
            O => \N__19736\,
            I => \N__19731\
        );

    \I__4540\ : CascadeMux
    port map (
            O => \N__19735\,
            I => \N__19728\
        );

    \I__4539\ : InMux
    port map (
            O => \N__19734\,
            I => \N__19725\
        );

    \I__4538\ : InMux
    port map (
            O => \N__19731\,
            I => \N__19720\
        );

    \I__4537\ : InMux
    port map (
            O => \N__19728\,
            I => \N__19720\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__19725\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__4535\ : LocalMux
    port map (
            O => \N__19720\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__4534\ : InMux
    port map (
            O => \N__19715\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__4533\ : CascadeMux
    port map (
            O => \N__19712\,
            I => \N__19707\
        );

    \I__4532\ : CascadeMux
    port map (
            O => \N__19711\,
            I => \N__19704\
        );

    \I__4531\ : InMux
    port map (
            O => \N__19710\,
            I => \N__19701\
        );

    \I__4530\ : InMux
    port map (
            O => \N__19707\,
            I => \N__19696\
        );

    \I__4529\ : InMux
    port map (
            O => \N__19704\,
            I => \N__19696\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__19701\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__19696\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__4526\ : InMux
    port map (
            O => \N__19691\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__4525\ : InMux
    port map (
            O => \N__19688\,
            I => \N__19683\
        );

    \I__4524\ : InMux
    port map (
            O => \N__19687\,
            I => \N__19680\
        );

    \I__4523\ : InMux
    port map (
            O => \N__19686\,
            I => \N__19677\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__19683\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__19680\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__19677\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__4519\ : InMux
    port map (
            O => \N__19670\,
            I => \bfn_10_24_0_\
        );

    \I__4518\ : InMux
    port map (
            O => \N__19667\,
            I => \N__19662\
        );

    \I__4517\ : InMux
    port map (
            O => \N__19666\,
            I => \N__19659\
        );

    \I__4516\ : InMux
    port map (
            O => \N__19665\,
            I => \N__19656\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__19662\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__19659\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__19656\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__4512\ : InMux
    port map (
            O => \N__19649\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__4511\ : InMux
    port map (
            O => \N__19646\,
            I => \N__19642\
        );

    \I__4510\ : InMux
    port map (
            O => \N__19645\,
            I => \N__19639\
        );

    \I__4509\ : LocalMux
    port map (
            O => \N__19642\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__19639\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__4507\ : CascadeMux
    port map (
            O => \N__19634\,
            I => \N__19629\
        );

    \I__4506\ : CascadeMux
    port map (
            O => \N__19633\,
            I => \N__19626\
        );

    \I__4505\ : InMux
    port map (
            O => \N__19632\,
            I => \N__19623\
        );

    \I__4504\ : InMux
    port map (
            O => \N__19629\,
            I => \N__19618\
        );

    \I__4503\ : InMux
    port map (
            O => \N__19626\,
            I => \N__19618\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__19623\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__19618\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__4500\ : InMux
    port map (
            O => \N__19613\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__4499\ : InMux
    port map (
            O => \N__19610\,
            I => \N__19606\
        );

    \I__4498\ : InMux
    port map (
            O => \N__19609\,
            I => \N__19603\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__19606\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__4496\ : LocalMux
    port map (
            O => \N__19603\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__4495\ : CascadeMux
    port map (
            O => \N__19598\,
            I => \N__19593\
        );

    \I__4494\ : CascadeMux
    port map (
            O => \N__19597\,
            I => \N__19590\
        );

    \I__4493\ : InMux
    port map (
            O => \N__19596\,
            I => \N__19587\
        );

    \I__4492\ : InMux
    port map (
            O => \N__19593\,
            I => \N__19582\
        );

    \I__4491\ : InMux
    port map (
            O => \N__19590\,
            I => \N__19582\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__19587\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__4489\ : LocalMux
    port map (
            O => \N__19582\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__4488\ : InMux
    port map (
            O => \N__19577\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__4487\ : InMux
    port map (
            O => \N__19574\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__4486\ : CascadeMux
    port map (
            O => \N__19571\,
            I => \N__19563\
        );

    \I__4485\ : CascadeMux
    port map (
            O => \N__19570\,
            I => \N__19554\
        );

    \I__4484\ : InMux
    port map (
            O => \N__19569\,
            I => \N__19546\
        );

    \I__4483\ : InMux
    port map (
            O => \N__19568\,
            I => \N__19546\
        );

    \I__4482\ : InMux
    port map (
            O => \N__19567\,
            I => \N__19546\
        );

    \I__4481\ : InMux
    port map (
            O => \N__19566\,
            I => \N__19543\
        );

    \I__4480\ : InMux
    port map (
            O => \N__19563\,
            I => \N__19532\
        );

    \I__4479\ : InMux
    port map (
            O => \N__19562\,
            I => \N__19532\
        );

    \I__4478\ : InMux
    port map (
            O => \N__19561\,
            I => \N__19532\
        );

    \I__4477\ : InMux
    port map (
            O => \N__19560\,
            I => \N__19532\
        );

    \I__4476\ : InMux
    port map (
            O => \N__19559\,
            I => \N__19532\
        );

    \I__4475\ : InMux
    port map (
            O => \N__19558\,
            I => \N__19527\
        );

    \I__4474\ : InMux
    port map (
            O => \N__19557\,
            I => \N__19527\
        );

    \I__4473\ : InMux
    port map (
            O => \N__19554\,
            I => \N__19524\
        );

    \I__4472\ : InMux
    port map (
            O => \N__19553\,
            I => \N__19521\
        );

    \I__4471\ : LocalMux
    port map (
            O => \N__19546\,
            I => \N__19516\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__19543\,
            I => \N__19516\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__19532\,
            I => \N__19509\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__19527\,
            I => \N__19509\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__19524\,
            I => \N__19509\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__19521\,
            I => \N__19504\
        );

    \I__4465\ : Span4Mux_v
    port map (
            O => \N__19516\,
            I => \N__19504\
        );

    \I__4464\ : Span4Mux_h
    port map (
            O => \N__19509\,
            I => \N__19501\
        );

    \I__4463\ : Odrv4
    port map (
            O => \N__19504\,
            I => \delay_measurement_inst.elapsed_time_hc_31\
        );

    \I__4462\ : Odrv4
    port map (
            O => \N__19501\,
            I => \delay_measurement_inst.elapsed_time_hc_31\
        );

    \I__4461\ : CEMux
    port map (
            O => \N__19496\,
            I => \N__19481\
        );

    \I__4460\ : CEMux
    port map (
            O => \N__19495\,
            I => \N__19481\
        );

    \I__4459\ : CEMux
    port map (
            O => \N__19494\,
            I => \N__19481\
        );

    \I__4458\ : CEMux
    port map (
            O => \N__19493\,
            I => \N__19481\
        );

    \I__4457\ : CEMux
    port map (
            O => \N__19492\,
            I => \N__19481\
        );

    \I__4456\ : GlobalMux
    port map (
            O => \N__19481\,
            I => \N__19478\
        );

    \I__4455\ : gio2CtrlBuf
    port map (
            O => \N__19478\,
            I => \delay_measurement_inst.delay_hc_timer.N_253_i_g\
        );

    \I__4454\ : InMux
    port map (
            O => \N__19475\,
            I => \N__19470\
        );

    \I__4453\ : InMux
    port map (
            O => \N__19474\,
            I => \N__19465\
        );

    \I__4452\ : InMux
    port map (
            O => \N__19473\,
            I => \N__19465\
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__19470\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__4450\ : LocalMux
    port map (
            O => \N__19465\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__4449\ : InMux
    port map (
            O => \N__19460\,
            I => \N__19455\
        );

    \I__4448\ : InMux
    port map (
            O => \N__19459\,
            I => \N__19452\
        );

    \I__4447\ : InMux
    port map (
            O => \N__19458\,
            I => \N__19449\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__19455\,
            I => \N__19446\
        );

    \I__4445\ : LocalMux
    port map (
            O => \N__19452\,
            I => \N__19441\
        );

    \I__4444\ : LocalMux
    port map (
            O => \N__19449\,
            I => \N__19441\
        );

    \I__4443\ : Span4Mux_v
    port map (
            O => \N__19446\,
            I => \N__19436\
        );

    \I__4442\ : Span4Mux_v
    port map (
            O => \N__19441\,
            I => \N__19436\
        );

    \I__4441\ : Odrv4
    port map (
            O => \N__19436\,
            I => \delay_measurement_inst.elapsed_time_hc_16\
        );

    \I__4440\ : InMux
    port map (
            O => \N__19433\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__4439\ : CascadeMux
    port map (
            O => \N__19430\,
            I => \N__19425\
        );

    \I__4438\ : CascadeMux
    port map (
            O => \N__19429\,
            I => \N__19422\
        );

    \I__4437\ : InMux
    port map (
            O => \N__19428\,
            I => \N__19419\
        );

    \I__4436\ : InMux
    port map (
            O => \N__19425\,
            I => \N__19414\
        );

    \I__4435\ : InMux
    port map (
            O => \N__19422\,
            I => \N__19414\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__19419\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__4433\ : LocalMux
    port map (
            O => \N__19414\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__4432\ : CascadeMux
    port map (
            O => \N__19409\,
            I => \N__19405\
        );

    \I__4431\ : InMux
    port map (
            O => \N__19408\,
            I => \N__19401\
        );

    \I__4430\ : InMux
    port map (
            O => \N__19405\,
            I => \N__19398\
        );

    \I__4429\ : InMux
    port map (
            O => \N__19404\,
            I => \N__19395\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__19401\,
            I => \N__19390\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__19398\,
            I => \N__19390\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__19395\,
            I => \N__19387\
        );

    \I__4425\ : Span4Mux_h
    port map (
            O => \N__19390\,
            I => \N__19384\
        );

    \I__4424\ : Odrv4
    port map (
            O => \N__19387\,
            I => \delay_measurement_inst.elapsed_time_hc_17\
        );

    \I__4423\ : Odrv4
    port map (
            O => \N__19384\,
            I => \delay_measurement_inst.elapsed_time_hc_17\
        );

    \I__4422\ : InMux
    port map (
            O => \N__19379\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__4421\ : CascadeMux
    port map (
            O => \N__19376\,
            I => \N__19371\
        );

    \I__4420\ : CascadeMux
    port map (
            O => \N__19375\,
            I => \N__19368\
        );

    \I__4419\ : InMux
    port map (
            O => \N__19374\,
            I => \N__19365\
        );

    \I__4418\ : InMux
    port map (
            O => \N__19371\,
            I => \N__19360\
        );

    \I__4417\ : InMux
    port map (
            O => \N__19368\,
            I => \N__19360\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__19365\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__19360\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__4414\ : InMux
    port map (
            O => \N__19355\,
            I => \N__19351\
        );

    \I__4413\ : InMux
    port map (
            O => \N__19354\,
            I => \N__19348\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__19351\,
            I => \N__19342\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__19348\,
            I => \N__19342\
        );

    \I__4410\ : InMux
    port map (
            O => \N__19347\,
            I => \N__19339\
        );

    \I__4409\ : Span4Mux_v
    port map (
            O => \N__19342\,
            I => \N__19334\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__19339\,
            I => \N__19334\
        );

    \I__4407\ : Odrv4
    port map (
            O => \N__19334\,
            I => \delay_measurement_inst.elapsed_time_hc_18\
        );

    \I__4406\ : InMux
    port map (
            O => \N__19331\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__4405\ : InMux
    port map (
            O => \N__19328\,
            I => \N__19323\
        );

    \I__4404\ : InMux
    port map (
            O => \N__19327\,
            I => \N__19320\
        );

    \I__4403\ : InMux
    port map (
            O => \N__19326\,
            I => \N__19317\
        );

    \I__4402\ : LocalMux
    port map (
            O => \N__19323\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__19320\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__19317\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__4399\ : CascadeMux
    port map (
            O => \N__19310\,
            I => \N__19305\
        );

    \I__4398\ : InMux
    port map (
            O => \N__19309\,
            I => \N__19302\
        );

    \I__4397\ : InMux
    port map (
            O => \N__19308\,
            I => \N__19299\
        );

    \I__4396\ : InMux
    port map (
            O => \N__19305\,
            I => \N__19296\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__19302\,
            I => \N__19293\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__19299\,
            I => \N__19288\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__19296\,
            I => \N__19288\
        );

    \I__4392\ : Span4Mux_h
    port map (
            O => \N__19293\,
            I => \N__19283\
        );

    \I__4391\ : Span4Mux_v
    port map (
            O => \N__19288\,
            I => \N__19283\
        );

    \I__4390\ : Odrv4
    port map (
            O => \N__19283\,
            I => \delay_measurement_inst.elapsed_time_hc_19\
        );

    \I__4389\ : InMux
    port map (
            O => \N__19280\,
            I => \bfn_10_23_0_\
        );

    \I__4388\ : InMux
    port map (
            O => \N__19277\,
            I => \N__19272\
        );

    \I__4387\ : InMux
    port map (
            O => \N__19276\,
            I => \N__19269\
        );

    \I__4386\ : InMux
    port map (
            O => \N__19275\,
            I => \N__19266\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__19272\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__19269\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__19266\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__4382\ : InMux
    port map (
            O => \N__19259\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__4381\ : CascadeMux
    port map (
            O => \N__19256\,
            I => \N__19251\
        );

    \I__4380\ : CascadeMux
    port map (
            O => \N__19255\,
            I => \N__19248\
        );

    \I__4379\ : InMux
    port map (
            O => \N__19254\,
            I => \N__19245\
        );

    \I__4378\ : InMux
    port map (
            O => \N__19251\,
            I => \N__19240\
        );

    \I__4377\ : InMux
    port map (
            O => \N__19248\,
            I => \N__19240\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__19245\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__19240\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__4374\ : InMux
    port map (
            O => \N__19235\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__4373\ : CascadeMux
    port map (
            O => \N__19232\,
            I => \N__19227\
        );

    \I__4372\ : CascadeMux
    port map (
            O => \N__19231\,
            I => \N__19224\
        );

    \I__4371\ : InMux
    port map (
            O => \N__19230\,
            I => \N__19221\
        );

    \I__4370\ : InMux
    port map (
            O => \N__19227\,
            I => \N__19216\
        );

    \I__4369\ : InMux
    port map (
            O => \N__19224\,
            I => \N__19216\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__19221\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__19216\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__4366\ : InMux
    port map (
            O => \N__19211\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__4365\ : InMux
    port map (
            O => \N__19208\,
            I => \N__19203\
        );

    \I__4364\ : InMux
    port map (
            O => \N__19207\,
            I => \N__19198\
        );

    \I__4363\ : InMux
    port map (
            O => \N__19206\,
            I => \N__19198\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__19203\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__4361\ : LocalMux
    port map (
            O => \N__19198\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__4360\ : InMux
    port map (
            O => \N__19193\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__4359\ : InMux
    port map (
            O => \N__19190\,
            I => \N__19185\
        );

    \I__4358\ : InMux
    port map (
            O => \N__19189\,
            I => \N__19180\
        );

    \I__4357\ : InMux
    port map (
            O => \N__19188\,
            I => \N__19180\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__19185\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__19180\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__4354\ : CascadeMux
    port map (
            O => \N__19175\,
            I => \N__19170\
        );

    \I__4353\ : CascadeMux
    port map (
            O => \N__19174\,
            I => \N__19167\
        );

    \I__4352\ : InMux
    port map (
            O => \N__19173\,
            I => \N__19164\
        );

    \I__4351\ : InMux
    port map (
            O => \N__19170\,
            I => \N__19159\
        );

    \I__4350\ : InMux
    port map (
            O => \N__19167\,
            I => \N__19159\
        );

    \I__4349\ : LocalMux
    port map (
            O => \N__19164\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__19159\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__4347\ : CascadeMux
    port map (
            O => \N__19154\,
            I => \N__19150\
        );

    \I__4346\ : CascadeMux
    port map (
            O => \N__19153\,
            I => \N__19147\
        );

    \I__4345\ : InMux
    port map (
            O => \N__19150\,
            I => \N__19141\
        );

    \I__4344\ : InMux
    port map (
            O => \N__19147\,
            I => \N__19136\
        );

    \I__4343\ : InMux
    port map (
            O => \N__19146\,
            I => \N__19136\
        );

    \I__4342\ : InMux
    port map (
            O => \N__19145\,
            I => \N__19131\
        );

    \I__4341\ : InMux
    port map (
            O => \N__19144\,
            I => \N__19131\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__19141\,
            I => \N__19128\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__19136\,
            I => \N__19125\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__19131\,
            I => \N__19122\
        );

    \I__4337\ : Span4Mux_h
    port map (
            O => \N__19128\,
            I => \N__19117\
        );

    \I__4336\ : Span4Mux_h
    port map (
            O => \N__19125\,
            I => \N__19117\
        );

    \I__4335\ : Span4Mux_h
    port map (
            O => \N__19122\,
            I => \N__19114\
        );

    \I__4334\ : Odrv4
    port map (
            O => \N__19117\,
            I => \delay_measurement_inst.delay_hc_reg3lto9\
        );

    \I__4333\ : Odrv4
    port map (
            O => \N__19114\,
            I => \delay_measurement_inst.delay_hc_reg3lto9\
        );

    \I__4332\ : InMux
    port map (
            O => \N__19109\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__4331\ : CascadeMux
    port map (
            O => \N__19106\,
            I => \N__19101\
        );

    \I__4330\ : CascadeMux
    port map (
            O => \N__19105\,
            I => \N__19098\
        );

    \I__4329\ : InMux
    port map (
            O => \N__19104\,
            I => \N__19095\
        );

    \I__4328\ : InMux
    port map (
            O => \N__19101\,
            I => \N__19090\
        );

    \I__4327\ : InMux
    port map (
            O => \N__19098\,
            I => \N__19090\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__19095\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__19090\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__4324\ : InMux
    port map (
            O => \N__19085\,
            I => \N__19081\
        );

    \I__4323\ : InMux
    port map (
            O => \N__19084\,
            I => \N__19078\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__19081\,
            I => \N__19073\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__19078\,
            I => \N__19073\
        );

    \I__4320\ : Span4Mux_h
    port map (
            O => \N__19073\,
            I => \N__19070\
        );

    \I__4319\ : Odrv4
    port map (
            O => \N__19070\,
            I => \delay_measurement_inst.elapsed_time_hc_10\
        );

    \I__4318\ : InMux
    port map (
            O => \N__19067\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__4317\ : InMux
    port map (
            O => \N__19064\,
            I => \N__19059\
        );

    \I__4316\ : InMux
    port map (
            O => \N__19063\,
            I => \N__19056\
        );

    \I__4315\ : InMux
    port map (
            O => \N__19062\,
            I => \N__19053\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__19059\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__19056\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__19053\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__4311\ : InMux
    port map (
            O => \N__19046\,
            I => \N__19042\
        );

    \I__4310\ : InMux
    port map (
            O => \N__19045\,
            I => \N__19039\
        );

    \I__4309\ : LocalMux
    port map (
            O => \N__19042\,
            I => \N__19036\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__19039\,
            I => \N__19033\
        );

    \I__4307\ : Odrv12
    port map (
            O => \N__19036\,
            I => \delay_measurement_inst.elapsed_time_hc_11\
        );

    \I__4306\ : Odrv4
    port map (
            O => \N__19033\,
            I => \delay_measurement_inst.elapsed_time_hc_11\
        );

    \I__4305\ : InMux
    port map (
            O => \N__19028\,
            I => \bfn_10_22_0_\
        );

    \I__4304\ : InMux
    port map (
            O => \N__19025\,
            I => \N__19020\
        );

    \I__4303\ : InMux
    port map (
            O => \N__19024\,
            I => \N__19017\
        );

    \I__4302\ : InMux
    port map (
            O => \N__19023\,
            I => \N__19014\
        );

    \I__4301\ : LocalMux
    port map (
            O => \N__19020\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__19017\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__19014\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__4298\ : InMux
    port map (
            O => \N__19007\,
            I => \N__19004\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__19004\,
            I => \N__19000\
        );

    \I__4296\ : InMux
    port map (
            O => \N__19003\,
            I => \N__18997\
        );

    \I__4295\ : Span4Mux_h
    port map (
            O => \N__19000\,
            I => \N__18992\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__18997\,
            I => \N__18992\
        );

    \I__4293\ : Odrv4
    port map (
            O => \N__18992\,
            I => \delay_measurement_inst.elapsed_time_hc_12\
        );

    \I__4292\ : InMux
    port map (
            O => \N__18989\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__4291\ : CascadeMux
    port map (
            O => \N__18986\,
            I => \N__18981\
        );

    \I__4290\ : CascadeMux
    port map (
            O => \N__18985\,
            I => \N__18978\
        );

    \I__4289\ : InMux
    port map (
            O => \N__18984\,
            I => \N__18975\
        );

    \I__4288\ : InMux
    port map (
            O => \N__18981\,
            I => \N__18970\
        );

    \I__4287\ : InMux
    port map (
            O => \N__18978\,
            I => \N__18970\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__18975\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__4285\ : LocalMux
    port map (
            O => \N__18970\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__4284\ : InMux
    port map (
            O => \N__18965\,
            I => \N__18961\
        );

    \I__4283\ : CascadeMux
    port map (
            O => \N__18964\,
            I => \N__18958\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__18961\,
            I => \N__18955\
        );

    \I__4281\ : InMux
    port map (
            O => \N__18958\,
            I => \N__18952\
        );

    \I__4280\ : Span4Mux_v
    port map (
            O => \N__18955\,
            I => \N__18949\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__18952\,
            I => \N__18946\
        );

    \I__4278\ : Odrv4
    port map (
            O => \N__18949\,
            I => \delay_measurement_inst.elapsed_time_hc_13\
        );

    \I__4277\ : Odrv4
    port map (
            O => \N__18946\,
            I => \delay_measurement_inst.elapsed_time_hc_13\
        );

    \I__4276\ : InMux
    port map (
            O => \N__18941\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__4275\ : CascadeMux
    port map (
            O => \N__18938\,
            I => \N__18933\
        );

    \I__4274\ : CascadeMux
    port map (
            O => \N__18937\,
            I => \N__18930\
        );

    \I__4273\ : InMux
    port map (
            O => \N__18936\,
            I => \N__18927\
        );

    \I__4272\ : InMux
    port map (
            O => \N__18933\,
            I => \N__18922\
        );

    \I__4271\ : InMux
    port map (
            O => \N__18930\,
            I => \N__18922\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__18927\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__18922\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__4268\ : CascadeMux
    port map (
            O => \N__18917\,
            I => \N__18912\
        );

    \I__4267\ : InMux
    port map (
            O => \N__18916\,
            I => \N__18907\
        );

    \I__4266\ : InMux
    port map (
            O => \N__18915\,
            I => \N__18902\
        );

    \I__4265\ : InMux
    port map (
            O => \N__18912\,
            I => \N__18902\
        );

    \I__4264\ : InMux
    port map (
            O => \N__18911\,
            I => \N__18899\
        );

    \I__4263\ : InMux
    port map (
            O => \N__18910\,
            I => \N__18896\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__18907\,
            I => \N__18893\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__18902\,
            I => \N__18890\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__18899\,
            I => \N__18885\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__18896\,
            I => \N__18885\
        );

    \I__4258\ : Span4Mux_h
    port map (
            O => \N__18893\,
            I => \N__18882\
        );

    \I__4257\ : Span4Mux_v
    port map (
            O => \N__18890\,
            I => \N__18877\
        );

    \I__4256\ : Span4Mux_h
    port map (
            O => \N__18885\,
            I => \N__18877\
        );

    \I__4255\ : Odrv4
    port map (
            O => \N__18882\,
            I => \delay_measurement_inst.delay_hc_reg3lto14\
        );

    \I__4254\ : Odrv4
    port map (
            O => \N__18877\,
            I => \delay_measurement_inst.delay_hc_reg3lto14\
        );

    \I__4253\ : InMux
    port map (
            O => \N__18872\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__4252\ : InMux
    port map (
            O => \N__18869\,
            I => \N__18864\
        );

    \I__4251\ : InMux
    port map (
            O => \N__18868\,
            I => \N__18859\
        );

    \I__4250\ : InMux
    port map (
            O => \N__18867\,
            I => \N__18859\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__18864\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__18859\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__4247\ : InMux
    port map (
            O => \N__18854\,
            I => \N__18846\
        );

    \I__4246\ : InMux
    port map (
            O => \N__18853\,
            I => \N__18846\
        );

    \I__4245\ : InMux
    port map (
            O => \N__18852\,
            I => \N__18840\
        );

    \I__4244\ : InMux
    port map (
            O => \N__18851\,
            I => \N__18840\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__18846\,
            I => \N__18834\
        );

    \I__4242\ : InMux
    port map (
            O => \N__18845\,
            I => \N__18831\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__18840\,
            I => \N__18828\
        );

    \I__4240\ : InMux
    port map (
            O => \N__18839\,
            I => \N__18825\
        );

    \I__4239\ : InMux
    port map (
            O => \N__18838\,
            I => \N__18820\
        );

    \I__4238\ : InMux
    port map (
            O => \N__18837\,
            I => \N__18820\
        );

    \I__4237\ : Span4Mux_v
    port map (
            O => \N__18834\,
            I => \N__18815\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__18831\,
            I => \N__18815\
        );

    \I__4235\ : Span4Mux_v
    port map (
            O => \N__18828\,
            I => \N__18812\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__18825\,
            I => \N__18809\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__18820\,
            I => \N__18806\
        );

    \I__4232\ : Span4Mux_v
    port map (
            O => \N__18815\,
            I => \N__18799\
        );

    \I__4231\ : Span4Mux_h
    port map (
            O => \N__18812\,
            I => \N__18799\
        );

    \I__4230\ : Span4Mux_v
    port map (
            O => \N__18809\,
            I => \N__18799\
        );

    \I__4229\ : Span4Mux_h
    port map (
            O => \N__18806\,
            I => \N__18796\
        );

    \I__4228\ : Odrv4
    port map (
            O => \N__18799\,
            I => \delay_measurement_inst.delay_hc_reg3lto15\
        );

    \I__4227\ : Odrv4
    port map (
            O => \N__18796\,
            I => \delay_measurement_inst.delay_hc_reg3lto15\
        );

    \I__4226\ : InMux
    port map (
            O => \N__18791\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__4225\ : InMux
    port map (
            O => \N__18788\,
            I => \N__18782\
        );

    \I__4224\ : InMux
    port map (
            O => \N__18787\,
            I => \N__18782\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__18782\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i\
        );

    \I__4222\ : InMux
    port map (
            O => \N__18779\,
            I => \N__18759\
        );

    \I__4221\ : InMux
    port map (
            O => \N__18778\,
            I => \N__18759\
        );

    \I__4220\ : InMux
    port map (
            O => \N__18777\,
            I => \N__18759\
        );

    \I__4219\ : InMux
    port map (
            O => \N__18776\,
            I => \N__18759\
        );

    \I__4218\ : InMux
    port map (
            O => \N__18775\,
            I => \N__18759\
        );

    \I__4217\ : InMux
    port map (
            O => \N__18774\,
            I => \N__18759\
        );

    \I__4216\ : InMux
    port map (
            O => \N__18773\,
            I => \N__18754\
        );

    \I__4215\ : InMux
    port map (
            O => \N__18772\,
            I => \N__18754\
        );

    \I__4214\ : LocalMux
    port map (
            O => \N__18759\,
            I => \delay_measurement_inst.N_41\
        );

    \I__4213\ : LocalMux
    port map (
            O => \N__18754\,
            I => \delay_measurement_inst.N_41\
        );

    \I__4212\ : InMux
    port map (
            O => \N__18749\,
            I => \N__18745\
        );

    \I__4211\ : InMux
    port map (
            O => \N__18748\,
            I => \N__18742\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__18745\,
            I => \N__18736\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__18742\,
            I => \N__18736\
        );

    \I__4208\ : InMux
    port map (
            O => \N__18741\,
            I => \N__18733\
        );

    \I__4207\ : Span4Mux_v
    port map (
            O => \N__18736\,
            I => \N__18728\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__18733\,
            I => \N__18728\
        );

    \I__4205\ : Odrv4
    port map (
            O => \N__18728\,
            I => \delay_measurement_inst.elapsed_time_tr_8\
        );

    \I__4204\ : InMux
    port map (
            O => \N__18725\,
            I => \N__18722\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__18722\,
            I => \N__18718\
        );

    \I__4202\ : CascadeMux
    port map (
            O => \N__18721\,
            I => \N__18714\
        );

    \I__4201\ : Span4Mux_v
    port map (
            O => \N__18718\,
            I => \N__18711\
        );

    \I__4200\ : InMux
    port map (
            O => \N__18717\,
            I => \N__18708\
        );

    \I__4199\ : InMux
    port map (
            O => \N__18714\,
            I => \N__18704\
        );

    \I__4198\ : Sp12to4
    port map (
            O => \N__18711\,
            I => \N__18699\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__18708\,
            I => \N__18699\
        );

    \I__4196\ : InMux
    port map (
            O => \N__18707\,
            I => \N__18696\
        );

    \I__4195\ : LocalMux
    port map (
            O => \N__18704\,
            I => measured_delay_tr_8
        );

    \I__4194\ : Odrv12
    port map (
            O => \N__18699\,
            I => measured_delay_tr_8
        );

    \I__4193\ : LocalMux
    port map (
            O => \N__18696\,
            I => measured_delay_tr_8
        );

    \I__4192\ : CascadeMux
    port map (
            O => \N__18689\,
            I => \N__18684\
        );

    \I__4191\ : CascadeMux
    port map (
            O => \N__18688\,
            I => \N__18673\
        );

    \I__4190\ : InMux
    port map (
            O => \N__18687\,
            I => \N__18670\
        );

    \I__4189\ : InMux
    port map (
            O => \N__18684\,
            I => \N__18667\
        );

    \I__4188\ : InMux
    port map (
            O => \N__18683\,
            I => \N__18664\
        );

    \I__4187\ : InMux
    port map (
            O => \N__18682\,
            I => \N__18649\
        );

    \I__4186\ : InMux
    port map (
            O => \N__18681\,
            I => \N__18649\
        );

    \I__4185\ : InMux
    port map (
            O => \N__18680\,
            I => \N__18649\
        );

    \I__4184\ : InMux
    port map (
            O => \N__18679\,
            I => \N__18649\
        );

    \I__4183\ : InMux
    port map (
            O => \N__18678\,
            I => \N__18649\
        );

    \I__4182\ : InMux
    port map (
            O => \N__18677\,
            I => \N__18649\
        );

    \I__4181\ : InMux
    port map (
            O => \N__18676\,
            I => \N__18649\
        );

    \I__4180\ : InMux
    port map (
            O => \N__18673\,
            I => \N__18644\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__18670\,
            I => \N__18641\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__18667\,
            I => \N__18634\
        );

    \I__4177\ : LocalMux
    port map (
            O => \N__18664\,
            I => \N__18634\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__18649\,
            I => \N__18634\
        );

    \I__4175\ : InMux
    port map (
            O => \N__18648\,
            I => \N__18629\
        );

    \I__4174\ : InMux
    port map (
            O => \N__18647\,
            I => \N__18629\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__18644\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__4172\ : Odrv4
    port map (
            O => \N__18641\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__4171\ : Odrv4
    port map (
            O => \N__18634\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__18629\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__4169\ : InMux
    port map (
            O => \N__18620\,
            I => \N__18617\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__18617\,
            I => \N__18613\
        );

    \I__4167\ : CascadeMux
    port map (
            O => \N__18616\,
            I => \N__18609\
        );

    \I__4166\ : Span4Mux_v
    port map (
            O => \N__18613\,
            I => \N__18606\
        );

    \I__4165\ : InMux
    port map (
            O => \N__18612\,
            I => \N__18603\
        );

    \I__4164\ : InMux
    port map (
            O => \N__18609\,
            I => \N__18600\
        );

    \I__4163\ : Odrv4
    port map (
            O => \N__18606\,
            I => \delay_measurement_inst.elapsed_time_tr_19\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__18603\,
            I => \delay_measurement_inst.elapsed_time_tr_19\
        );

    \I__4161\ : LocalMux
    port map (
            O => \N__18600\,
            I => \delay_measurement_inst.elapsed_time_tr_19\
        );

    \I__4160\ : InMux
    port map (
            O => \N__18593\,
            I => \N__18583\
        );

    \I__4159\ : InMux
    port map (
            O => \N__18592\,
            I => \N__18583\
        );

    \I__4158\ : InMux
    port map (
            O => \N__18591\,
            I => \N__18583\
        );

    \I__4157\ : InMux
    port map (
            O => \N__18590\,
            I => \N__18580\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__18583\,
            I => \N__18570\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__18580\,
            I => \N__18570\
        );

    \I__4154\ : InMux
    port map (
            O => \N__18579\,
            I => \N__18567\
        );

    \I__4153\ : InMux
    port map (
            O => \N__18578\,
            I => \N__18558\
        );

    \I__4152\ : InMux
    port map (
            O => \N__18577\,
            I => \N__18558\
        );

    \I__4151\ : InMux
    port map (
            O => \N__18576\,
            I => \N__18558\
        );

    \I__4150\ : InMux
    port map (
            O => \N__18575\,
            I => \N__18558\
        );

    \I__4149\ : Odrv4
    port map (
            O => \N__18570\,
            I => \delay_measurement_inst.N_35\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__18567\,
            I => \delay_measurement_inst.N_35\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__18558\,
            I => \delay_measurement_inst.N_35\
        );

    \I__4146\ : InMux
    port map (
            O => \N__18551\,
            I => \N__18548\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__18548\,
            I => \N__18543\
        );

    \I__4144\ : InMux
    port map (
            O => \N__18547\,
            I => \N__18540\
        );

    \I__4143\ : CascadeMux
    port map (
            O => \N__18546\,
            I => \N__18537\
        );

    \I__4142\ : Span4Mux_v
    port map (
            O => \N__18543\,
            I => \N__18534\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__18540\,
            I => \N__18531\
        );

    \I__4140\ : InMux
    port map (
            O => \N__18537\,
            I => \N__18528\
        );

    \I__4139\ : Span4Mux_h
    port map (
            O => \N__18534\,
            I => \N__18520\
        );

    \I__4138\ : Span4Mux_v
    port map (
            O => \N__18531\,
            I => \N__18520\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__18528\,
            I => \N__18520\
        );

    \I__4136\ : CascadeMux
    port map (
            O => \N__18527\,
            I => \N__18517\
        );

    \I__4135\ : Span4Mux_h
    port map (
            O => \N__18520\,
            I => \N__18514\
        );

    \I__4134\ : InMux
    port map (
            O => \N__18517\,
            I => \N__18511\
        );

    \I__4133\ : Odrv4
    port map (
            O => \N__18514\,
            I => measured_delay_tr_19
        );

    \I__4132\ : LocalMux
    port map (
            O => \N__18511\,
            I => measured_delay_tr_19
        );

    \I__4131\ : CEMux
    port map (
            O => \N__18506\,
            I => \N__18502\
        );

    \I__4130\ : CEMux
    port map (
            O => \N__18505\,
            I => \N__18498\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__18502\,
            I => \N__18495\
        );

    \I__4128\ : CEMux
    port map (
            O => \N__18501\,
            I => \N__18492\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__18498\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\
        );

    \I__4126\ : Odrv12
    port map (
            O => \N__18495\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__18492\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\
        );

    \I__4124\ : InMux
    port map (
            O => \N__18485\,
            I => \N__18480\
        );

    \I__4123\ : InMux
    port map (
            O => \N__18484\,
            I => \N__18477\
        );

    \I__4122\ : InMux
    port map (
            O => \N__18483\,
            I => \N__18474\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__18480\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__18477\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__18474\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__4118\ : CascadeMux
    port map (
            O => \N__18467\,
            I => \N__18464\
        );

    \I__4117\ : InMux
    port map (
            O => \N__18464\,
            I => \N__18459\
        );

    \I__4116\ : InMux
    port map (
            O => \N__18463\,
            I => \N__18454\
        );

    \I__4115\ : InMux
    port map (
            O => \N__18462\,
            I => \N__18454\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__18459\,
            I => \N__18449\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__18454\,
            I => \N__18449\
        );

    \I__4112\ : Span4Mux_h
    port map (
            O => \N__18449\,
            I => \N__18446\
        );

    \I__4111\ : Odrv4
    port map (
            O => \N__18446\,
            I => \delay_measurement_inst.elapsed_time_hc_3\
        );

    \I__4110\ : InMux
    port map (
            O => \N__18443\,
            I => \N__18438\
        );

    \I__4109\ : InMux
    port map (
            O => \N__18442\,
            I => \N__18435\
        );

    \I__4108\ : InMux
    port map (
            O => \N__18441\,
            I => \N__18432\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__18438\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__18435\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__18432\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__4104\ : CascadeMux
    port map (
            O => \N__18425\,
            I => \N__18422\
        );

    \I__4103\ : InMux
    port map (
            O => \N__18422\,
            I => \N__18419\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__18419\,
            I => \N__18416\
        );

    \I__4101\ : Span4Mux_v
    port map (
            O => \N__18416\,
            I => \N__18412\
        );

    \I__4100\ : InMux
    port map (
            O => \N__18415\,
            I => \N__18409\
        );

    \I__4099\ : Sp12to4
    port map (
            O => \N__18412\,
            I => \N__18404\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__18409\,
            I => \N__18404\
        );

    \I__4097\ : Odrv12
    port map (
            O => \N__18404\,
            I => \delay_measurement_inst.elapsed_time_hc_4\
        );

    \I__4096\ : InMux
    port map (
            O => \N__18401\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__4095\ : CascadeMux
    port map (
            O => \N__18398\,
            I => \N__18393\
        );

    \I__4094\ : CascadeMux
    port map (
            O => \N__18397\,
            I => \N__18390\
        );

    \I__4093\ : InMux
    port map (
            O => \N__18396\,
            I => \N__18387\
        );

    \I__4092\ : InMux
    port map (
            O => \N__18393\,
            I => \N__18382\
        );

    \I__4091\ : InMux
    port map (
            O => \N__18390\,
            I => \N__18382\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__18387\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__18382\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__4088\ : InMux
    port map (
            O => \N__18377\,
            I => \N__18374\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__18374\,
            I => \N__18370\
        );

    \I__4086\ : InMux
    port map (
            O => \N__18373\,
            I => \N__18367\
        );

    \I__4085\ : Span4Mux_v
    port map (
            O => \N__18370\,
            I => \N__18362\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__18367\,
            I => \N__18362\
        );

    \I__4083\ : Odrv4
    port map (
            O => \N__18362\,
            I => \delay_measurement_inst.elapsed_time_hc_5\
        );

    \I__4082\ : InMux
    port map (
            O => \N__18359\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__4081\ : CascadeMux
    port map (
            O => \N__18356\,
            I => \N__18351\
        );

    \I__4080\ : CascadeMux
    port map (
            O => \N__18355\,
            I => \N__18348\
        );

    \I__4079\ : InMux
    port map (
            O => \N__18354\,
            I => \N__18345\
        );

    \I__4078\ : InMux
    port map (
            O => \N__18351\,
            I => \N__18340\
        );

    \I__4077\ : InMux
    port map (
            O => \N__18348\,
            I => \N__18340\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__18345\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__18340\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__4074\ : CascadeMux
    port map (
            O => \N__18335\,
            I => \N__18332\
        );

    \I__4073\ : InMux
    port map (
            O => \N__18332\,
            I => \N__18327\
        );

    \I__4072\ : InMux
    port map (
            O => \N__18331\,
            I => \N__18321\
        );

    \I__4071\ : InMux
    port map (
            O => \N__18330\,
            I => \N__18321\
        );

    \I__4070\ : LocalMux
    port map (
            O => \N__18327\,
            I => \N__18318\
        );

    \I__4069\ : InMux
    port map (
            O => \N__18326\,
            I => \N__18315\
        );

    \I__4068\ : LocalMux
    port map (
            O => \N__18321\,
            I => \N__18312\
        );

    \I__4067\ : Span4Mux_v
    port map (
            O => \N__18318\,
            I => \N__18307\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__18315\,
            I => \N__18307\
        );

    \I__4065\ : Span4Mux_h
    port map (
            O => \N__18312\,
            I => \N__18304\
        );

    \I__4064\ : Odrv4
    port map (
            O => \N__18307\,
            I => \delay_measurement_inst.delay_hc_reg3lto6\
        );

    \I__4063\ : Odrv4
    port map (
            O => \N__18304\,
            I => \delay_measurement_inst.delay_hc_reg3lto6\
        );

    \I__4062\ : InMux
    port map (
            O => \N__18299\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__4061\ : InMux
    port map (
            O => \N__18296\,
            I => \N__18291\
        );

    \I__4060\ : InMux
    port map (
            O => \N__18295\,
            I => \N__18286\
        );

    \I__4059\ : InMux
    port map (
            O => \N__18294\,
            I => \N__18286\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__18291\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__18286\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__4056\ : CascadeMux
    port map (
            O => \N__18281\,
            I => \N__18278\
        );

    \I__4055\ : InMux
    port map (
            O => \N__18278\,
            I => \N__18274\
        );

    \I__4054\ : InMux
    port map (
            O => \N__18277\,
            I => \N__18271\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__18274\,
            I => \N__18268\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__18271\,
            I => \N__18265\
        );

    \I__4051\ : Span4Mux_h
    port map (
            O => \N__18268\,
            I => \N__18262\
        );

    \I__4050\ : Span4Mux_h
    port map (
            O => \N__18265\,
            I => \N__18259\
        );

    \I__4049\ : Odrv4
    port map (
            O => \N__18262\,
            I => \delay_measurement_inst.elapsed_time_hc_7\
        );

    \I__4048\ : Odrv4
    port map (
            O => \N__18259\,
            I => \delay_measurement_inst.elapsed_time_hc_7\
        );

    \I__4047\ : InMux
    port map (
            O => \N__18254\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__4046\ : InMux
    port map (
            O => \N__18251\,
            I => \N__18246\
        );

    \I__4045\ : InMux
    port map (
            O => \N__18250\,
            I => \N__18241\
        );

    \I__4044\ : InMux
    port map (
            O => \N__18249\,
            I => \N__18241\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__18246\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__4042\ : LocalMux
    port map (
            O => \N__18241\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__4041\ : CascadeMux
    port map (
            O => \N__18236\,
            I => \N__18232\
        );

    \I__4040\ : CascadeMux
    port map (
            O => \N__18235\,
            I => \N__18229\
        );

    \I__4039\ : InMux
    port map (
            O => \N__18232\,
            I => \N__18226\
        );

    \I__4038\ : InMux
    port map (
            O => \N__18229\,
            I => \N__18223\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__18226\,
            I => \N__18220\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__18223\,
            I => \N__18217\
        );

    \I__4035\ : Span4Mux_h
    port map (
            O => \N__18220\,
            I => \N__18214\
        );

    \I__4034\ : Span4Mux_h
    port map (
            O => \N__18217\,
            I => \N__18211\
        );

    \I__4033\ : Odrv4
    port map (
            O => \N__18214\,
            I => \delay_measurement_inst.elapsed_time_hc_8\
        );

    \I__4032\ : Odrv4
    port map (
            O => \N__18211\,
            I => \delay_measurement_inst.elapsed_time_hc_8\
        );

    \I__4031\ : InMux
    port map (
            O => \N__18206\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__4030\ : InMux
    port map (
            O => \N__18203\,
            I => \N__18200\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__18200\,
            I => \delay_measurement_inst.N_164\
        );

    \I__4028\ : InMux
    port map (
            O => \N__18197\,
            I => \N__18179\
        );

    \I__4027\ : InMux
    port map (
            O => \N__18196\,
            I => \N__18179\
        );

    \I__4026\ : InMux
    port map (
            O => \N__18195\,
            I => \N__18179\
        );

    \I__4025\ : InMux
    port map (
            O => \N__18194\,
            I => \N__18179\
        );

    \I__4024\ : InMux
    port map (
            O => \N__18193\,
            I => \N__18179\
        );

    \I__4023\ : InMux
    port map (
            O => \N__18192\,
            I => \N__18179\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__18179\,
            I => \delay_measurement_inst.N_187\
        );

    \I__4021\ : InMux
    port map (
            O => \N__18176\,
            I => \N__18173\
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__18173\,
            I => \N__18170\
        );

    \I__4019\ : Odrv4
    port map (
            O => \N__18170\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_7\
        );

    \I__4018\ : CascadeMux
    port map (
            O => \N__18167\,
            I => \delay_measurement_inst.N_187_cascade_\
        );

    \I__4017\ : InMux
    port map (
            O => \N__18164\,
            I => \N__18161\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__18161\,
            I => \delay_measurement_inst.delay_tr_timer.N_177\
        );

    \I__4015\ : CascadeMux
    port map (
            O => \N__18158\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i_cascade_\
        );

    \I__4014\ : CascadeMux
    port map (
            O => \N__18155\,
            I => \N__18152\
        );

    \I__4013\ : InMux
    port map (
            O => \N__18152\,
            I => \N__18136\
        );

    \I__4012\ : InMux
    port map (
            O => \N__18151\,
            I => \N__18136\
        );

    \I__4011\ : InMux
    port map (
            O => \N__18150\,
            I => \N__18136\
        );

    \I__4010\ : InMux
    port map (
            O => \N__18149\,
            I => \N__18136\
        );

    \I__4009\ : InMux
    port map (
            O => \N__18148\,
            I => \N__18136\
        );

    \I__4008\ : InMux
    port map (
            O => \N__18147\,
            I => \N__18133\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__18136\,
            I => \delay_measurement_inst.N_162_1\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__18133\,
            I => \delay_measurement_inst.N_162_1\
        );

    \I__4005\ : CascadeMux
    port map (
            O => \N__18128\,
            I => \N__18123\
        );

    \I__4004\ : InMux
    port map (
            O => \N__18127\,
            I => \N__18115\
        );

    \I__4003\ : InMux
    port map (
            O => \N__18126\,
            I => \N__18115\
        );

    \I__4002\ : InMux
    port map (
            O => \N__18123\,
            I => \N__18115\
        );

    \I__4001\ : InMux
    port map (
            O => \N__18122\,
            I => \N__18112\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__18115\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__18112\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10\
        );

    \I__3998\ : CascadeMux
    port map (
            O => \N__18107\,
            I => \N__18102\
        );

    \I__3997\ : CascadeMux
    port map (
            O => \N__18106\,
            I => \N__18099\
        );

    \I__3996\ : InMux
    port map (
            O => \N__18105\,
            I => \N__18096\
        );

    \I__3995\ : InMux
    port map (
            O => \N__18102\,
            I => \N__18093\
        );

    \I__3994\ : InMux
    port map (
            O => \N__18099\,
            I => \N__18090\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__18096\,
            I => \N__18086\
        );

    \I__3992\ : LocalMux
    port map (
            O => \N__18093\,
            I => \N__18081\
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__18090\,
            I => \N__18081\
        );

    \I__3990\ : InMux
    port map (
            O => \N__18089\,
            I => \N__18078\
        );

    \I__3989\ : Span4Mux_v
    port map (
            O => \N__18086\,
            I => \N__18074\
        );

    \I__3988\ : Span4Mux_v
    port map (
            O => \N__18081\,
            I => \N__18069\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__18078\,
            I => \N__18069\
        );

    \I__3986\ : InMux
    port map (
            O => \N__18077\,
            I => \N__18066\
        );

    \I__3985\ : Odrv4
    port map (
            O => \N__18074\,
            I => \delay_measurement_inst.delay_tr_reg3lto9\
        );

    \I__3984\ : Odrv4
    port map (
            O => \N__18069\,
            I => \delay_measurement_inst.delay_tr_reg3lto9\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__18066\,
            I => \delay_measurement_inst.delay_tr_reg3lto9\
        );

    \I__3982\ : InMux
    port map (
            O => \N__18059\,
            I => \N__18053\
        );

    \I__3981\ : InMux
    port map (
            O => \N__18058\,
            I => \N__18050\
        );

    \I__3980\ : InMux
    port map (
            O => \N__18057\,
            I => \N__18047\
        );

    \I__3979\ : CascadeMux
    port map (
            O => \N__18056\,
            I => \N__18044\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__18053\,
            I => \N__18040\
        );

    \I__3977\ : LocalMux
    port map (
            O => \N__18050\,
            I => \N__18035\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__18047\,
            I => \N__18035\
        );

    \I__3975\ : InMux
    port map (
            O => \N__18044\,
            I => \N__18030\
        );

    \I__3974\ : InMux
    port map (
            O => \N__18043\,
            I => \N__18030\
        );

    \I__3973\ : Odrv12
    port map (
            O => \N__18040\,
            I => \delay_measurement_inst.delay_tr_reg3lto14\
        );

    \I__3972\ : Odrv4
    port map (
            O => \N__18035\,
            I => \delay_measurement_inst.delay_tr_reg3lto14\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__18030\,
            I => \delay_measurement_inst.delay_tr_reg3lto14\
        );

    \I__3970\ : InMux
    port map (
            O => \N__18023\,
            I => \N__18019\
        );

    \I__3969\ : CascadeMux
    port map (
            O => \N__18022\,
            I => \N__18015\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__18019\,
            I => \N__18012\
        );

    \I__3967\ : InMux
    port map (
            O => \N__18018\,
            I => \N__18009\
        );

    \I__3966\ : InMux
    port map (
            O => \N__18015\,
            I => \N__18006\
        );

    \I__3965\ : Span4Mux_h
    port map (
            O => \N__18012\,
            I => \N__18002\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__18009\,
            I => \N__17999\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__18006\,
            I => \N__17996\
        );

    \I__3962\ : InMux
    port map (
            O => \N__18005\,
            I => \N__17993\
        );

    \I__3961\ : Odrv4
    port map (
            O => \N__18002\,
            I => \delay_measurement_inst.N_39\
        );

    \I__3960\ : Odrv4
    port map (
            O => \N__17999\,
            I => \delay_measurement_inst.N_39\
        );

    \I__3959\ : Odrv4
    port map (
            O => \N__17996\,
            I => \delay_measurement_inst.N_39\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__17993\,
            I => \delay_measurement_inst.N_39\
        );

    \I__3957\ : CascadeMux
    port map (
            O => \N__17984\,
            I => \delay_measurement_inst.delay_tr_timer.N_180_cascade_\
        );

    \I__3956\ : CascadeMux
    port map (
            O => \N__17981\,
            I => \N__17978\
        );

    \I__3955\ : InMux
    port map (
            O => \N__17978\,
            I => \N__17974\
        );

    \I__3954\ : InMux
    port map (
            O => \N__17977\,
            I => \N__17971\
        );

    \I__3953\ : LocalMux
    port map (
            O => \N__17974\,
            I => \N__17967\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__17971\,
            I => \N__17964\
        );

    \I__3951\ : InMux
    port map (
            O => \N__17970\,
            I => \N__17961\
        );

    \I__3950\ : Span4Mux_v
    port map (
            O => \N__17967\,
            I => \N__17957\
        );

    \I__3949\ : Span4Mux_v
    port map (
            O => \N__17964\,
            I => \N__17952\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__17961\,
            I => \N__17952\
        );

    \I__3947\ : InMux
    port map (
            O => \N__17960\,
            I => \N__17949\
        );

    \I__3946\ : Odrv4
    port map (
            O => \N__17957\,
            I => \delay_measurement_inst.delay_tr_reg3lto6\
        );

    \I__3945\ : Odrv4
    port map (
            O => \N__17952\,
            I => \delay_measurement_inst.delay_tr_reg3lto6\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__17949\,
            I => \delay_measurement_inst.delay_tr_reg3lto6\
        );

    \I__3943\ : InMux
    port map (
            O => \N__17942\,
            I => \N__17932\
        );

    \I__3942\ : InMux
    port map (
            O => \N__17941\,
            I => \N__17932\
        );

    \I__3941\ : InMux
    port map (
            O => \N__17940\,
            I => \N__17927\
        );

    \I__3940\ : InMux
    port map (
            O => \N__17939\,
            I => \N__17927\
        );

    \I__3939\ : InMux
    port map (
            O => \N__17938\,
            I => \N__17922\
        );

    \I__3938\ : InMux
    port map (
            O => \N__17937\,
            I => \N__17922\
        );

    \I__3937\ : LocalMux
    port map (
            O => \N__17932\,
            I => \N__17913\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__17927\,
            I => \N__17913\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__17922\,
            I => \N__17913\
        );

    \I__3934\ : InMux
    port map (
            O => \N__17921\,
            I => \N__17908\
        );

    \I__3933\ : InMux
    port map (
            O => \N__17920\,
            I => \N__17908\
        );

    \I__3932\ : Odrv4
    port map (
            O => \N__17913\,
            I => \delay_measurement_inst.delay_tr_reg3lto15\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__17908\,
            I => \delay_measurement_inst.delay_tr_reg3lto15\
        );

    \I__3930\ : CascadeMux
    port map (
            O => \N__17903\,
            I => \N__17896\
        );

    \I__3929\ : CascadeMux
    port map (
            O => \N__17902\,
            I => \N__17893\
        );

    \I__3928\ : InMux
    port map (
            O => \N__17901\,
            I => \N__17882\
        );

    \I__3927\ : InMux
    port map (
            O => \N__17900\,
            I => \N__17882\
        );

    \I__3926\ : InMux
    port map (
            O => \N__17899\,
            I => \N__17882\
        );

    \I__3925\ : InMux
    port map (
            O => \N__17896\,
            I => \N__17882\
        );

    \I__3924\ : InMux
    port map (
            O => \N__17893\,
            I => \N__17882\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__17882\,
            I => \delay_measurement_inst.delay_tr_reg_5_0_a2_0_6\
        );

    \I__3922\ : InMux
    port map (
            O => \N__17879\,
            I => \N__17875\
        );

    \I__3921\ : InMux
    port map (
            O => \N__17878\,
            I => \N__17872\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__17875\,
            I => \N__17866\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__17872\,
            I => \N__17866\
        );

    \I__3918\ : InMux
    port map (
            O => \N__17871\,
            I => \N__17863\
        );

    \I__3917\ : Span4Mux_v
    port map (
            O => \N__17866\,
            I => \N__17858\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__17863\,
            I => \N__17858\
        );

    \I__3915\ : Odrv4
    port map (
            O => \N__17858\,
            I => \delay_measurement_inst.elapsed_time_tr_7\
        );

    \I__3914\ : InMux
    port map (
            O => \N__17855\,
            I => \N__17852\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__17852\,
            I => \N__17846\
        );

    \I__3912\ : InMux
    port map (
            O => \N__17851\,
            I => \N__17843\
        );

    \I__3911\ : CascadeMux
    port map (
            O => \N__17850\,
            I => \N__17840\
        );

    \I__3910\ : CascadeMux
    port map (
            O => \N__17849\,
            I => \N__17837\
        );

    \I__3909\ : Span4Mux_v
    port map (
            O => \N__17846\,
            I => \N__17834\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__17843\,
            I => \N__17831\
        );

    \I__3907\ : InMux
    port map (
            O => \N__17840\,
            I => \N__17828\
        );

    \I__3906\ : InMux
    port map (
            O => \N__17837\,
            I => \N__17825\
        );

    \I__3905\ : Span4Mux_h
    port map (
            O => \N__17834\,
            I => \N__17820\
        );

    \I__3904\ : Span4Mux_h
    port map (
            O => \N__17831\,
            I => \N__17820\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__17828\,
            I => \N__17817\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__17825\,
            I => measured_delay_tr_7
        );

    \I__3901\ : Odrv4
    port map (
            O => \N__17820\,
            I => measured_delay_tr_7
        );

    \I__3900\ : Odrv4
    port map (
            O => \N__17817\,
            I => measured_delay_tr_7
        );

    \I__3899\ : InMux
    port map (
            O => \N__17810\,
            I => \N__17804\
        );

    \I__3898\ : InMux
    port map (
            O => \N__17809\,
            I => \N__17804\
        );

    \I__3897\ : LocalMux
    port map (
            O => \N__17804\,
            I => \delay_measurement_inst.delay_tr_timer.N_177_4\
        );

    \I__3896\ : InMux
    port map (
            O => \N__17801\,
            I => \N__17798\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__17798\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_4\
        );

    \I__3894\ : CascadeMux
    port map (
            O => \N__17795\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3_cascade_\
        );

    \I__3893\ : InMux
    port map (
            O => \N__17792\,
            I => \N__17789\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__17789\,
            I => \N__17784\
        );

    \I__3891\ : InMux
    port map (
            O => \N__17788\,
            I => \N__17779\
        );

    \I__3890\ : InMux
    port map (
            O => \N__17787\,
            I => \N__17779\
        );

    \I__3889\ : Odrv12
    port map (
            O => \N__17784\,
            I => \delay_measurement_inst.elapsed_time_tr_16\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__17779\,
            I => \delay_measurement_inst.elapsed_time_tr_16\
        );

    \I__3887\ : InMux
    port map (
            O => \N__17774\,
            I => \N__17770\
        );

    \I__3886\ : CascadeMux
    port map (
            O => \N__17773\,
            I => \N__17766\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__17770\,
            I => \N__17763\
        );

    \I__3884\ : InMux
    port map (
            O => \N__17769\,
            I => \N__17760\
        );

    \I__3883\ : InMux
    port map (
            O => \N__17766\,
            I => \N__17757\
        );

    \I__3882\ : Odrv12
    port map (
            O => \N__17763\,
            I => \delay_measurement_inst.elapsed_time_tr_17\
        );

    \I__3881\ : LocalMux
    port map (
            O => \N__17760\,
            I => \delay_measurement_inst.elapsed_time_tr_17\
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__17757\,
            I => \delay_measurement_inst.elapsed_time_tr_17\
        );

    \I__3879\ : InMux
    port map (
            O => \N__17750\,
            I => \N__17747\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__17747\,
            I => \N__17742\
        );

    \I__3877\ : InMux
    port map (
            O => \N__17746\,
            I => \N__17739\
        );

    \I__3876\ : InMux
    port map (
            O => \N__17745\,
            I => \N__17736\
        );

    \I__3875\ : Odrv12
    port map (
            O => \N__17742\,
            I => \delay_measurement_inst.elapsed_time_tr_18\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__17739\,
            I => \delay_measurement_inst.elapsed_time_tr_18\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__17736\,
            I => \delay_measurement_inst.elapsed_time_tr_18\
        );

    \I__3872\ : InMux
    port map (
            O => \N__17729\,
            I => \N__17726\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__17726\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\
        );

    \I__3870\ : InMux
    port map (
            O => \N__17723\,
            I => \N__17720\
        );

    \I__3869\ : LocalMux
    port map (
            O => \N__17720\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__3868\ : InMux
    port map (
            O => \N__17717\,
            I => \N__17713\
        );

    \I__3867\ : InMux
    port map (
            O => \N__17716\,
            I => \N__17710\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__17713\,
            I => \N__17707\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__17710\,
            I => \N__17704\
        );

    \I__3864\ : Span4Mux_h
    port map (
            O => \N__17707\,
            I => \N__17701\
        );

    \I__3863\ : Odrv12
    port map (
            O => \N__17704\,
            I => \delay_measurement_inst.elapsed_time_tr_12\
        );

    \I__3862\ : Odrv4
    port map (
            O => \N__17701\,
            I => \delay_measurement_inst.elapsed_time_tr_12\
        );

    \I__3861\ : InMux
    port map (
            O => \N__17696\,
            I => \N__17692\
        );

    \I__3860\ : InMux
    port map (
            O => \N__17695\,
            I => \N__17689\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__17692\,
            I => \N__17686\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__17689\,
            I => \N__17683\
        );

    \I__3857\ : Span4Mux_h
    port map (
            O => \N__17686\,
            I => \N__17680\
        );

    \I__3856\ : Odrv12
    port map (
            O => \N__17683\,
            I => \delay_measurement_inst.elapsed_time_tr_11\
        );

    \I__3855\ : Odrv4
    port map (
            O => \N__17680\,
            I => \delay_measurement_inst.elapsed_time_tr_11\
        );

    \I__3854\ : InMux
    port map (
            O => \N__17675\,
            I => \N__17671\
        );

    \I__3853\ : CascadeMux
    port map (
            O => \N__17674\,
            I => \N__17668\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__17671\,
            I => \N__17665\
        );

    \I__3851\ : InMux
    port map (
            O => \N__17668\,
            I => \N__17662\
        );

    \I__3850\ : Span4Mux_v
    port map (
            O => \N__17665\,
            I => \N__17657\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__17662\,
            I => \N__17657\
        );

    \I__3848\ : Odrv4
    port map (
            O => \N__17657\,
            I => \delay_measurement_inst.elapsed_time_tr_13\
        );

    \I__3847\ : InMux
    port map (
            O => \N__17654\,
            I => \N__17650\
        );

    \I__3846\ : InMux
    port map (
            O => \N__17653\,
            I => \N__17647\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__17650\,
            I => \N__17644\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__17647\,
            I => \N__17641\
        );

    \I__3843\ : Odrv12
    port map (
            O => \N__17644\,
            I => \delay_measurement_inst.elapsed_time_tr_10\
        );

    \I__3842\ : Odrv4
    port map (
            O => \N__17641\,
            I => \delay_measurement_inst.elapsed_time_tr_10\
        );

    \I__3841\ : InMux
    port map (
            O => \N__17636\,
            I => \N__17633\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__17633\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__3839\ : InMux
    port map (
            O => \N__17630\,
            I => \N__17627\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__17627\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__3837\ : CascadeMux
    port map (
            O => \N__17624\,
            I => \N__17621\
        );

    \I__3836\ : InMux
    port map (
            O => \N__17621\,
            I => \N__17618\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__17618\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__3834\ : InMux
    port map (
            O => \N__17615\,
            I => \N__17612\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__17612\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__3832\ : InMux
    port map (
            O => \N__17609\,
            I => \N__17606\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__17606\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__3830\ : InMux
    port map (
            O => \N__17603\,
            I => \N__17600\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__17600\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19\
        );

    \I__3828\ : CascadeMux
    port map (
            O => \N__17597\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19_cascade_\
        );

    \I__3827\ : InMux
    port map (
            O => \N__17594\,
            I => \N__17591\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__17591\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19\
        );

    \I__3825\ : InMux
    port map (
            O => \N__17588\,
            I => \N__17585\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__17585\,
            I => \N__17582\
        );

    \I__3823\ : Odrv4
    port map (
            O => \N__17582\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6\
        );

    \I__3822\ : CascadeMux
    port map (
            O => \N__17579\,
            I => \delay_measurement_inst.N_35_cascade_\
        );

    \I__3821\ : InMux
    port map (
            O => \N__17576\,
            I => \N__17573\
        );

    \I__3820\ : LocalMux
    port map (
            O => \N__17573\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_7\
        );

    \I__3819\ : CascadeMux
    port map (
            O => \N__17570\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_\
        );

    \I__3818\ : InMux
    port map (
            O => \N__17567\,
            I => \N__17533\
        );

    \I__3817\ : InMux
    port map (
            O => \N__17566\,
            I => \N__17533\
        );

    \I__3816\ : InMux
    port map (
            O => \N__17565\,
            I => \N__17533\
        );

    \I__3815\ : InMux
    port map (
            O => \N__17564\,
            I => \N__17533\
        );

    \I__3814\ : InMux
    port map (
            O => \N__17563\,
            I => \N__17524\
        );

    \I__3813\ : InMux
    port map (
            O => \N__17562\,
            I => \N__17524\
        );

    \I__3812\ : InMux
    port map (
            O => \N__17561\,
            I => \N__17515\
        );

    \I__3811\ : InMux
    port map (
            O => \N__17560\,
            I => \N__17515\
        );

    \I__3810\ : InMux
    port map (
            O => \N__17559\,
            I => \N__17515\
        );

    \I__3809\ : InMux
    port map (
            O => \N__17558\,
            I => \N__17515\
        );

    \I__3808\ : InMux
    port map (
            O => \N__17557\,
            I => \N__17506\
        );

    \I__3807\ : InMux
    port map (
            O => \N__17556\,
            I => \N__17506\
        );

    \I__3806\ : InMux
    port map (
            O => \N__17555\,
            I => \N__17506\
        );

    \I__3805\ : InMux
    port map (
            O => \N__17554\,
            I => \N__17506\
        );

    \I__3804\ : InMux
    port map (
            O => \N__17553\,
            I => \N__17497\
        );

    \I__3803\ : InMux
    port map (
            O => \N__17552\,
            I => \N__17497\
        );

    \I__3802\ : InMux
    port map (
            O => \N__17551\,
            I => \N__17497\
        );

    \I__3801\ : InMux
    port map (
            O => \N__17550\,
            I => \N__17497\
        );

    \I__3800\ : InMux
    port map (
            O => \N__17549\,
            I => \N__17488\
        );

    \I__3799\ : InMux
    port map (
            O => \N__17548\,
            I => \N__17488\
        );

    \I__3798\ : InMux
    port map (
            O => \N__17547\,
            I => \N__17488\
        );

    \I__3797\ : InMux
    port map (
            O => \N__17546\,
            I => \N__17488\
        );

    \I__3796\ : InMux
    port map (
            O => \N__17545\,
            I => \N__17479\
        );

    \I__3795\ : InMux
    port map (
            O => \N__17544\,
            I => \N__17479\
        );

    \I__3794\ : InMux
    port map (
            O => \N__17543\,
            I => \N__17479\
        );

    \I__3793\ : InMux
    port map (
            O => \N__17542\,
            I => \N__17479\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__17533\,
            I => \N__17476\
        );

    \I__3791\ : InMux
    port map (
            O => \N__17532\,
            I => \N__17467\
        );

    \I__3790\ : InMux
    port map (
            O => \N__17531\,
            I => \N__17467\
        );

    \I__3789\ : InMux
    port map (
            O => \N__17530\,
            I => \N__17467\
        );

    \I__3788\ : InMux
    port map (
            O => \N__17529\,
            I => \N__17467\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__17524\,
            I => \N__17464\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__17515\,
            I => \N__17459\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__17506\,
            I => \N__17459\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__17497\,
            I => \N__17452\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__17488\,
            I => \N__17452\
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__17479\,
            I => \N__17452\
        );

    \I__3781\ : Span4Mux_v
    port map (
            O => \N__17476\,
            I => \N__17441\
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__17467\,
            I => \N__17441\
        );

    \I__3779\ : Span4Mux_v
    port map (
            O => \N__17464\,
            I => \N__17441\
        );

    \I__3778\ : Span4Mux_v
    port map (
            O => \N__17459\,
            I => \N__17441\
        );

    \I__3777\ : Span4Mux_v
    port map (
            O => \N__17452\,
            I => \N__17441\
        );

    \I__3776\ : Odrv4
    port map (
            O => \N__17441\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__3775\ : CascadeMux
    port map (
            O => \N__17438\,
            I => \N__17435\
        );

    \I__3774\ : InMux
    port map (
            O => \N__17435\,
            I => \N__17432\
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__17432\,
            I => \N__17429\
        );

    \I__3772\ : Span4Mux_v
    port map (
            O => \N__17429\,
            I => \N__17425\
        );

    \I__3771\ : InMux
    port map (
            O => \N__17428\,
            I => \N__17422\
        );

    \I__3770\ : Odrv4
    port map (
            O => \N__17425\,
            I => \delay_measurement_inst.elapsed_time_tr_5\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__17422\,
            I => \delay_measurement_inst.elapsed_time_tr_5\
        );

    \I__3768\ : InMux
    port map (
            O => \N__17417\,
            I => \N__17414\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__17414\,
            I => \N__17410\
        );

    \I__3766\ : InMux
    port map (
            O => \N__17413\,
            I => \N__17407\
        );

    \I__3765\ : Odrv12
    port map (
            O => \N__17410\,
            I => \delay_measurement_inst.elapsed_time_tr_4\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__17407\,
            I => \delay_measurement_inst.elapsed_time_tr_4\
        );

    \I__3763\ : CascadeMux
    port map (
            O => \N__17402\,
            I => \N__17399\
        );

    \I__3762\ : InMux
    port map (
            O => \N__17399\,
            I => \N__17396\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__17396\,
            I => \N__17392\
        );

    \I__3760\ : InMux
    port map (
            O => \N__17395\,
            I => \N__17389\
        );

    \I__3759\ : Span4Mux_v
    port map (
            O => \N__17392\,
            I => \N__17383\
        );

    \I__3758\ : LocalMux
    port map (
            O => \N__17389\,
            I => \N__17383\
        );

    \I__3757\ : InMux
    port map (
            O => \N__17388\,
            I => \N__17380\
        );

    \I__3756\ : Odrv4
    port map (
            O => \N__17383\,
            I => \delay_measurement_inst.elapsed_time_tr_3\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__17380\,
            I => \delay_measurement_inst.elapsed_time_tr_3\
        );

    \I__3754\ : CascadeMux
    port map (
            O => \N__17375\,
            I => \N__17372\
        );

    \I__3753\ : InMux
    port map (
            O => \N__17372\,
            I => \N__17368\
        );

    \I__3752\ : CascadeMux
    port map (
            O => \N__17371\,
            I => \N__17365\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__17368\,
            I => \N__17362\
        );

    \I__3750\ : InMux
    port map (
            O => \N__17365\,
            I => \N__17359\
        );

    \I__3749\ : Span4Mux_v
    port map (
            O => \N__17362\,
            I => \N__17356\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__17359\,
            I => \N__17353\
        );

    \I__3747\ : Odrv4
    port map (
            O => \N__17356\,
            I => \delay_measurement_inst.elapsed_time_tr_1\
        );

    \I__3746\ : Odrv12
    port map (
            O => \N__17353\,
            I => \delay_measurement_inst.elapsed_time_tr_1\
        );

    \I__3745\ : InMux
    port map (
            O => \N__17348\,
            I => \N__17345\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__17345\,
            I => \N__17341\
        );

    \I__3743\ : InMux
    port map (
            O => \N__17344\,
            I => \N__17338\
        );

    \I__3742\ : Span4Mux_v
    port map (
            O => \N__17341\,
            I => \N__17332\
        );

    \I__3741\ : LocalMux
    port map (
            O => \N__17338\,
            I => \N__17332\
        );

    \I__3740\ : InMux
    port map (
            O => \N__17337\,
            I => \N__17329\
        );

    \I__3739\ : Odrv4
    port map (
            O => \N__17332\,
            I => \delay_measurement_inst.elapsed_time_tr_2\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__17329\,
            I => \delay_measurement_inst.elapsed_time_tr_2\
        );

    \I__3737\ : InMux
    port map (
            O => \N__17324\,
            I => \N__17321\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__17321\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__3735\ : InMux
    port map (
            O => \N__17318\,
            I => \N__17315\
        );

    \I__3734\ : LocalMux
    port map (
            O => \N__17315\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__3733\ : CascadeMux
    port map (
            O => \N__17312\,
            I => \N__17309\
        );

    \I__3732\ : InMux
    port map (
            O => \N__17309\,
            I => \N__17306\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__17306\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__3730\ : InMux
    port map (
            O => \N__17303\,
            I => \N__17300\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__17300\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__3728\ : CascadeMux
    port map (
            O => \N__17297\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_5_cascade_\
        );

    \I__3727\ : InMux
    port map (
            O => \N__17294\,
            I => \bfn_9_24_0_\
        );

    \I__3726\ : InMux
    port map (
            O => \N__17291\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_24\
        );

    \I__3725\ : InMux
    port map (
            O => \N__17288\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_25\
        );

    \I__3724\ : InMux
    port map (
            O => \N__17285\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_26\
        );

    \I__3723\ : InMux
    port map (
            O => \N__17282\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_27\
        );

    \I__3722\ : InMux
    port map (
            O => \N__17279\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_28\
        );

    \I__3721\ : InMux
    port map (
            O => \N__17276\,
            I => \N__17273\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__17273\,
            I => \N__17270\
        );

    \I__3719\ : Span4Mux_s1_v
    port map (
            O => \N__17270\,
            I => \N__17267\
        );

    \I__3718\ : Span4Mux_v
    port map (
            O => \N__17267\,
            I => \N__17261\
        );

    \I__3717\ : InMux
    port map (
            O => \N__17266\,
            I => \N__17258\
        );

    \I__3716\ : InMux
    port map (
            O => \N__17265\,
            I => \N__17255\
        );

    \I__3715\ : InMux
    port map (
            O => \N__17264\,
            I => \N__17252\
        );

    \I__3714\ : Odrv4
    port map (
            O => \N__17261\,
            I => \phase_controller_slave.stateZ0Z_3\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__17258\,
            I => \phase_controller_slave.stateZ0Z_3\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__17255\,
            I => \phase_controller_slave.stateZ0Z_3\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__17252\,
            I => \phase_controller_slave.stateZ0Z_3\
        );

    \I__3710\ : IoInMux
    port map (
            O => \N__17243\,
            I => \N__17240\
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__17240\,
            I => s3_phy_c
        );

    \I__3708\ : InMux
    port map (
            O => \N__17237\,
            I => \N__17234\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__17234\,
            I => \N__17229\
        );

    \I__3706\ : InMux
    port map (
            O => \N__17233\,
            I => \N__17226\
        );

    \I__3705\ : InMux
    port map (
            O => \N__17232\,
            I => \N__17223\
        );

    \I__3704\ : Odrv4
    port map (
            O => \N__17229\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__17226\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__17223\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__3701\ : InMux
    port map (
            O => \N__17216\,
            I => \N__17213\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__17213\,
            I => \N__17208\
        );

    \I__3699\ : InMux
    port map (
            O => \N__17212\,
            I => \N__17205\
        );

    \I__3698\ : InMux
    port map (
            O => \N__17211\,
            I => \N__17202\
        );

    \I__3697\ : Odrv4
    port map (
            O => \N__17208\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__17205\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__17202\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__3694\ : CEMux
    port map (
            O => \N__17195\,
            I => \N__17180\
        );

    \I__3693\ : CEMux
    port map (
            O => \N__17194\,
            I => \N__17180\
        );

    \I__3692\ : CEMux
    port map (
            O => \N__17193\,
            I => \N__17180\
        );

    \I__3691\ : CEMux
    port map (
            O => \N__17192\,
            I => \N__17180\
        );

    \I__3690\ : CEMux
    port map (
            O => \N__17191\,
            I => \N__17180\
        );

    \I__3689\ : GlobalMux
    port map (
            O => \N__17180\,
            I => \N__17177\
        );

    \I__3688\ : gio2CtrlBuf
    port map (
            O => \N__17177\,
            I => \delay_measurement_inst.delay_tr_timer.N_255_i_g\
        );

    \I__3687\ : InMux
    port map (
            O => \N__17174\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_14\
        );

    \I__3686\ : InMux
    port map (
            O => \N__17171\,
            I => \bfn_9_23_0_\
        );

    \I__3685\ : InMux
    port map (
            O => \N__17168\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_16\
        );

    \I__3684\ : InMux
    port map (
            O => \N__17165\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_17\
        );

    \I__3683\ : InMux
    port map (
            O => \N__17162\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_18\
        );

    \I__3682\ : InMux
    port map (
            O => \N__17159\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_19\
        );

    \I__3681\ : InMux
    port map (
            O => \N__17156\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_20\
        );

    \I__3680\ : InMux
    port map (
            O => \N__17153\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_21\
        );

    \I__3679\ : InMux
    port map (
            O => \N__17150\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_22\
        );

    \I__3678\ : InMux
    port map (
            O => \N__17147\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_5\
        );

    \I__3677\ : InMux
    port map (
            O => \N__17144\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_6\
        );

    \I__3676\ : InMux
    port map (
            O => \N__17141\,
            I => \bfn_9_22_0_\
        );

    \I__3675\ : InMux
    port map (
            O => \N__17138\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_8\
        );

    \I__3674\ : InMux
    port map (
            O => \N__17135\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_9\
        );

    \I__3673\ : InMux
    port map (
            O => \N__17132\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_10\
        );

    \I__3672\ : InMux
    port map (
            O => \N__17129\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_11\
        );

    \I__3671\ : InMux
    port map (
            O => \N__17126\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_12\
        );

    \I__3670\ : InMux
    port map (
            O => \N__17123\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_13\
        );

    \I__3669\ : InMux
    port map (
            O => \N__17120\,
            I => \N__17117\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__17117\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3\
        );

    \I__3667\ : CascadeMux
    port map (
            O => \N__17114\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_9_cascade_\
        );

    \I__3666\ : InMux
    port map (
            O => \N__17111\,
            I => \N__17107\
        );

    \I__3665\ : InMux
    port map (
            O => \N__17110\,
            I => \N__17104\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__17107\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_0_6\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__17104\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_0_6\
        );

    \I__3662\ : InMux
    port map (
            O => \N__17099\,
            I => \N__17096\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__17096\,
            I => \N__17093\
        );

    \I__3660\ : Span4Mux_h
    port map (
            O => \N__17093\,
            I => \N__17089\
        );

    \I__3659\ : InMux
    port map (
            O => \N__17092\,
            I => \N__17086\
        );

    \I__3658\ : Span4Mux_h
    port map (
            O => \N__17089\,
            I => \N__17082\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__17086\,
            I => \N__17079\
        );

    \I__3656\ : InMux
    port map (
            O => \N__17085\,
            I => \N__17076\
        );

    \I__3655\ : Odrv4
    port map (
            O => \N__17082\,
            I => \phase_controller_inst1.stoper_tr.N_97\
        );

    \I__3654\ : Odrv12
    port map (
            O => \N__17079\,
            I => \phase_controller_inst1.stoper_tr.N_97\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__17076\,
            I => \phase_controller_inst1.stoper_tr.N_97\
        );

    \I__3652\ : InMux
    port map (
            O => \N__17069\,
            I => \N__17065\
        );

    \I__3651\ : InMux
    port map (
            O => \N__17068\,
            I => \N__17062\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__17065\,
            I => \N__17058\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__17062\,
            I => \N__17055\
        );

    \I__3648\ : InMux
    port map (
            O => \N__17061\,
            I => \N__17052\
        );

    \I__3647\ : Span12Mux_s9_h
    port map (
            O => \N__17058\,
            I => \N__17049\
        );

    \I__3646\ : Span4Mux_h
    port map (
            O => \N__17055\,
            I => \N__17044\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__17052\,
            I => \N__17044\
        );

    \I__3644\ : Odrv12
    port map (
            O => \N__17049\,
            I => measured_delay_tr_4
        );

    \I__3643\ : Odrv4
    port map (
            O => \N__17044\,
            I => measured_delay_tr_4
        );

    \I__3642\ : InMux
    port map (
            O => \N__17039\,
            I => \N__17035\
        );

    \I__3641\ : InMux
    port map (
            O => \N__17038\,
            I => \N__17032\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__17035\,
            I => \N__17026\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__17032\,
            I => \N__17026\
        );

    \I__3638\ : InMux
    port map (
            O => \N__17031\,
            I => \N__17023\
        );

    \I__3637\ : Span4Mux_v
    port map (
            O => \N__17026\,
            I => \N__17017\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__17023\,
            I => \N__17017\
        );

    \I__3635\ : InMux
    port map (
            O => \N__17022\,
            I => \N__17013\
        );

    \I__3634\ : Span4Mux_h
    port map (
            O => \N__17017\,
            I => \N__17010\
        );

    \I__3633\ : InMux
    port map (
            O => \N__17016\,
            I => \N__17007\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__17013\,
            I => measured_delay_tr_14
        );

    \I__3631\ : Odrv4
    port map (
            O => \N__17010\,
            I => measured_delay_tr_14
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__17007\,
            I => measured_delay_tr_14
        );

    \I__3629\ : InMux
    port map (
            O => \N__17000\,
            I => \N__16987\
        );

    \I__3628\ : InMux
    port map (
            O => \N__16999\,
            I => \N__16987\
        );

    \I__3627\ : InMux
    port map (
            O => \N__16998\,
            I => \N__16987\
        );

    \I__3626\ : InMux
    port map (
            O => \N__16997\,
            I => \N__16984\
        );

    \I__3625\ : InMux
    port map (
            O => \N__16996\,
            I => \N__16979\
        );

    \I__3624\ : InMux
    port map (
            O => \N__16995\,
            I => \N__16979\
        );

    \I__3623\ : InMux
    port map (
            O => \N__16994\,
            I => \N__16976\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__16987\,
            I => \N__16973\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__16984\,
            I => \N__16966\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__16979\,
            I => \N__16966\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__16976\,
            I => \N__16966\
        );

    \I__3618\ : Span4Mux_v
    port map (
            O => \N__16973\,
            I => \N__16960\
        );

    \I__3617\ : Span4Mux_v
    port map (
            O => \N__16966\,
            I => \N__16957\
        );

    \I__3616\ : InMux
    port map (
            O => \N__16965\,
            I => \N__16952\
        );

    \I__3615\ : InMux
    port map (
            O => \N__16964\,
            I => \N__16952\
        );

    \I__3614\ : CascadeMux
    port map (
            O => \N__16963\,
            I => \N__16949\
        );

    \I__3613\ : Span4Mux_h
    port map (
            O => \N__16960\,
            I => \N__16942\
        );

    \I__3612\ : Span4Mux_h
    port map (
            O => \N__16957\,
            I => \N__16942\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__16952\,
            I => \N__16942\
        );

    \I__3610\ : InMux
    port map (
            O => \N__16949\,
            I => \N__16939\
        );

    \I__3609\ : Sp12to4
    port map (
            O => \N__16942\,
            I => \N__16934\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__16939\,
            I => \N__16934\
        );

    \I__3607\ : Odrv12
    port map (
            O => \N__16934\,
            I => measured_delay_tr_15
        );

    \I__3606\ : InMux
    port map (
            O => \N__16931\,
            I => \N__16928\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__16928\,
            I => \N__16924\
        );

    \I__3604\ : InMux
    port map (
            O => \N__16927\,
            I => \N__16921\
        );

    \I__3603\ : Span4Mux_v
    port map (
            O => \N__16924\,
            I => \N__16915\
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__16921\,
            I => \N__16915\
        );

    \I__3601\ : InMux
    port map (
            O => \N__16920\,
            I => \N__16912\
        );

    \I__3600\ : Span4Mux_h
    port map (
            O => \N__16915\,
            I => \N__16907\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__16912\,
            I => \N__16907\
        );

    \I__3598\ : Odrv4
    port map (
            O => \N__16907\,
            I => measured_delay_tr_5
        );

    \I__3597\ : InMux
    port map (
            O => \N__16904\,
            I => \N__16901\
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__16901\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3\
        );

    \I__3595\ : InMux
    port map (
            O => \N__16898\,
            I => \N__16895\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__16895\,
            I => \N__16892\
        );

    \I__3593\ : Span4Mux_h
    port map (
            O => \N__16892\,
            I => \N__16886\
        );

    \I__3592\ : CascadeMux
    port map (
            O => \N__16891\,
            I => \N__16883\
        );

    \I__3591\ : CascadeMux
    port map (
            O => \N__16890\,
            I => \N__16880\
        );

    \I__3590\ : InMux
    port map (
            O => \N__16889\,
            I => \N__16877\
        );

    \I__3589\ : Span4Mux_v
    port map (
            O => \N__16886\,
            I => \N__16874\
        );

    \I__3588\ : InMux
    port map (
            O => \N__16883\,
            I => \N__16869\
        );

    \I__3587\ : InMux
    port map (
            O => \N__16880\,
            I => \N__16869\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__16877\,
            I => \N__16866\
        );

    \I__3585\ : Odrv4
    port map (
            O => \N__16874\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__16869\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__3583\ : Odrv4
    port map (
            O => \N__16866\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__3582\ : IoInMux
    port map (
            O => \N__16859\,
            I => \N__16856\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__16856\,
            I => \N__16853\
        );

    \I__3580\ : Span4Mux_s2_v
    port map (
            O => \N__16853\,
            I => \N__16850\
        );

    \I__3579\ : Span4Mux_h
    port map (
            O => \N__16850\,
            I => \N__16847\
        );

    \I__3578\ : Span4Mux_v
    port map (
            O => \N__16847\,
            I => \N__16844\
        );

    \I__3577\ : Span4Mux_v
    port map (
            O => \N__16844\,
            I => \N__16841\
        );

    \I__3576\ : Odrv4
    port map (
            O => \N__16841\,
            I => s1_phy_c
        );

    \I__3575\ : InMux
    port map (
            O => \N__16838\,
            I => \bfn_9_21_0_\
        );

    \I__3574\ : InMux
    port map (
            O => \N__16835\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_0\
        );

    \I__3573\ : InMux
    port map (
            O => \N__16832\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_1\
        );

    \I__3572\ : InMux
    port map (
            O => \N__16829\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_2\
        );

    \I__3571\ : InMux
    port map (
            O => \N__16826\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_3\
        );

    \I__3570\ : InMux
    port map (
            O => \N__16823\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_4\
        );

    \I__3569\ : InMux
    port map (
            O => \N__16820\,
            I => \N__16816\
        );

    \I__3568\ : InMux
    port map (
            O => \N__16819\,
            I => \N__16813\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__16816\,
            I => \N__16808\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__16813\,
            I => \N__16808\
        );

    \I__3565\ : Span4Mux_v
    port map (
            O => \N__16808\,
            I => \N__16804\
        );

    \I__3564\ : InMux
    port map (
            O => \N__16807\,
            I => \N__16801\
        );

    \I__3563\ : Span4Mux_h
    port map (
            O => \N__16804\,
            I => \N__16796\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__16801\,
            I => \N__16796\
        );

    \I__3561\ : Odrv4
    port map (
            O => \N__16796\,
            I => measured_delay_tr_6
        );

    \I__3560\ : InMux
    port map (
            O => \N__16793\,
            I => \N__16789\
        );

    \I__3559\ : InMux
    port map (
            O => \N__16792\,
            I => \N__16786\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__16789\,
            I => \N__16783\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__16786\,
            I => \N__16779\
        );

    \I__3556\ : Span4Mux_h
    port map (
            O => \N__16783\,
            I => \N__16775\
        );

    \I__3555\ : InMux
    port map (
            O => \N__16782\,
            I => \N__16772\
        );

    \I__3554\ : Span4Mux_h
    port map (
            O => \N__16779\,
            I => \N__16769\
        );

    \I__3553\ : InMux
    port map (
            O => \N__16778\,
            I => \N__16766\
        );

    \I__3552\ : Span4Mux_h
    port map (
            O => \N__16775\,
            I => \N__16761\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__16772\,
            I => \N__16761\
        );

    \I__3550\ : Odrv4
    port map (
            O => \N__16769\,
            I => measured_delay_tr_18
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__16766\,
            I => measured_delay_tr_18
        );

    \I__3548\ : Odrv4
    port map (
            O => \N__16761\,
            I => measured_delay_tr_18
        );

    \I__3547\ : InMux
    port map (
            O => \N__16754\,
            I => \N__16751\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__16751\,
            I => \N__16747\
        );

    \I__3545\ : InMux
    port map (
            O => \N__16750\,
            I => \N__16744\
        );

    \I__3544\ : Span4Mux_h
    port map (
            O => \N__16747\,
            I => \N__16741\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__16744\,
            I => \N__16738\
        );

    \I__3542\ : Span4Mux_h
    port map (
            O => \N__16741\,
            I => \N__16733\
        );

    \I__3541\ : Span4Mux_h
    port map (
            O => \N__16738\,
            I => \N__16730\
        );

    \I__3540\ : InMux
    port map (
            O => \N__16737\,
            I => \N__16727\
        );

    \I__3539\ : InMux
    port map (
            O => \N__16736\,
            I => \N__16724\
        );

    \I__3538\ : Odrv4
    port map (
            O => \N__16733\,
            I => measured_delay_tr_17
        );

    \I__3537\ : Odrv4
    port map (
            O => \N__16730\,
            I => measured_delay_tr_17
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__16727\,
            I => measured_delay_tr_17
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__16724\,
            I => measured_delay_tr_17
        );

    \I__3534\ : InMux
    port map (
            O => \N__16715\,
            I => \N__16712\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__16712\,
            I => \N__16708\
        );

    \I__3532\ : InMux
    port map (
            O => \N__16711\,
            I => \N__16705\
        );

    \I__3531\ : Span4Mux_v
    port map (
            O => \N__16708\,
            I => \N__16702\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__16705\,
            I => \N__16699\
        );

    \I__3529\ : Span4Mux_h
    port map (
            O => \N__16702\,
            I => \N__16694\
        );

    \I__3528\ : Span4Mux_v
    port map (
            O => \N__16699\,
            I => \N__16691\
        );

    \I__3527\ : InMux
    port map (
            O => \N__16698\,
            I => \N__16688\
        );

    \I__3526\ : InMux
    port map (
            O => \N__16697\,
            I => \N__16685\
        );

    \I__3525\ : Odrv4
    port map (
            O => \N__16694\,
            I => measured_delay_tr_16
        );

    \I__3524\ : Odrv4
    port map (
            O => \N__16691\,
            I => measured_delay_tr_16
        );

    \I__3523\ : LocalMux
    port map (
            O => \N__16688\,
            I => measured_delay_tr_16
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__16685\,
            I => measured_delay_tr_16
        );

    \I__3521\ : InMux
    port map (
            O => \N__16676\,
            I => \N__16673\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__16673\,
            I => \N__16669\
        );

    \I__3519\ : InMux
    port map (
            O => \N__16672\,
            I => \N__16666\
        );

    \I__3518\ : Span12Mux_v
    port map (
            O => \N__16669\,
            I => \N__16660\
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__16666\,
            I => \N__16660\
        );

    \I__3516\ : InMux
    port map (
            O => \N__16665\,
            I => \N__16657\
        );

    \I__3515\ : Odrv12
    port map (
            O => \N__16660\,
            I => measured_delay_tr_12
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__16657\,
            I => measured_delay_tr_12
        );

    \I__3513\ : InMux
    port map (
            O => \N__16652\,
            I => \N__16649\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__16649\,
            I => \N__16646\
        );

    \I__3511\ : Span4Mux_h
    port map (
            O => \N__16646\,
            I => \N__16642\
        );

    \I__3510\ : InMux
    port map (
            O => \N__16645\,
            I => \N__16639\
        );

    \I__3509\ : Span4Mux_h
    port map (
            O => \N__16642\,
            I => \N__16635\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__16639\,
            I => \N__16632\
        );

    \I__3507\ : InMux
    port map (
            O => \N__16638\,
            I => \N__16629\
        );

    \I__3506\ : Odrv4
    port map (
            O => \N__16635\,
            I => measured_delay_tr_11
        );

    \I__3505\ : Odrv12
    port map (
            O => \N__16632\,
            I => measured_delay_tr_11
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__16629\,
            I => measured_delay_tr_11
        );

    \I__3503\ : InMux
    port map (
            O => \N__16622\,
            I => \N__16619\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__16619\,
            I => \N__16615\
        );

    \I__3501\ : InMux
    port map (
            O => \N__16618\,
            I => \N__16612\
        );

    \I__3500\ : Span4Mux_h
    port map (
            O => \N__16615\,
            I => \N__16606\
        );

    \I__3499\ : LocalMux
    port map (
            O => \N__16612\,
            I => \N__16606\
        );

    \I__3498\ : CascadeMux
    port map (
            O => \N__16611\,
            I => \N__16603\
        );

    \I__3497\ : Span4Mux_h
    port map (
            O => \N__16606\,
            I => \N__16600\
        );

    \I__3496\ : InMux
    port map (
            O => \N__16603\,
            I => \N__16597\
        );

    \I__3495\ : Odrv4
    port map (
            O => \N__16600\,
            I => measured_delay_tr_13
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__16597\,
            I => measured_delay_tr_13
        );

    \I__3493\ : InMux
    port map (
            O => \N__16592\,
            I => \N__16589\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__16589\,
            I => \N__16585\
        );

    \I__3491\ : InMux
    port map (
            O => \N__16588\,
            I => \N__16582\
        );

    \I__3490\ : Span4Mux_h
    port map (
            O => \N__16585\,
            I => \N__16577\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__16582\,
            I => \N__16577\
        );

    \I__3488\ : Span4Mux_h
    port map (
            O => \N__16577\,
            I => \N__16573\
        );

    \I__3487\ : InMux
    port map (
            O => \N__16576\,
            I => \N__16570\
        );

    \I__3486\ : Odrv4
    port map (
            O => \N__16573\,
            I => measured_delay_tr_10
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__16570\,
            I => measured_delay_tr_10
        );

    \I__3484\ : CascadeMux
    port map (
            O => \N__16565\,
            I => \N__16561\
        );

    \I__3483\ : InMux
    port map (
            O => \N__16564\,
            I => \N__16558\
        );

    \I__3482\ : InMux
    port map (
            O => \N__16561\,
            I => \N__16555\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__16558\,
            I => \N__16552\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__16555\,
            I => \N__16549\
        );

    \I__3479\ : Span4Mux_h
    port map (
            O => \N__16552\,
            I => \N__16543\
        );

    \I__3478\ : Span4Mux_v
    port map (
            O => \N__16549\,
            I => \N__16543\
        );

    \I__3477\ : InMux
    port map (
            O => \N__16548\,
            I => \N__16540\
        );

    \I__3476\ : Span4Mux_h
    port map (
            O => \N__16543\,
            I => \N__16535\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__16540\,
            I => \N__16535\
        );

    \I__3474\ : Odrv4
    port map (
            O => \N__16535\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_0_6\
        );

    \I__3473\ : CascadeMux
    port map (
            O => \N__16532\,
            I => \N__16528\
        );

    \I__3472\ : InMux
    port map (
            O => \N__16531\,
            I => \N__16525\
        );

    \I__3471\ : InMux
    port map (
            O => \N__16528\,
            I => \N__16522\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__16525\,
            I => \N__16519\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__16522\,
            I => \N__16516\
        );

    \I__3468\ : Span4Mux_v
    port map (
            O => \N__16519\,
            I => \N__16510\
        );

    \I__3467\ : Span4Mux_h
    port map (
            O => \N__16516\,
            I => \N__16510\
        );

    \I__3466\ : InMux
    port map (
            O => \N__16515\,
            I => \N__16507\
        );

    \I__3465\ : Span4Mux_h
    port map (
            O => \N__16510\,
            I => \N__16504\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__16507\,
            I => \N__16501\
        );

    \I__3463\ : Odrv4
    port map (
            O => \N__16504\,
            I => measured_delay_tr_9
        );

    \I__3462\ : Odrv4
    port map (
            O => \N__16501\,
            I => measured_delay_tr_9
        );

    \I__3461\ : CascadeMux
    port map (
            O => \N__16496\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_0_6_cascade_\
        );

    \I__3460\ : InMux
    port map (
            O => \N__16493\,
            I => \N__16490\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__16490\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_9\
        );

    \I__3458\ : CascadeMux
    port map (
            O => \N__16487\,
            I => \N__16484\
        );

    \I__3457\ : InMux
    port map (
            O => \N__16484\,
            I => \N__16480\
        );

    \I__3456\ : CascadeMux
    port map (
            O => \N__16483\,
            I => \N__16477\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__16480\,
            I => \N__16474\
        );

    \I__3454\ : InMux
    port map (
            O => \N__16477\,
            I => \N__16471\
        );

    \I__3453\ : Span4Mux_v
    port map (
            O => \N__16474\,
            I => \N__16466\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__16471\,
            I => \N__16466\
        );

    \I__3451\ : Span4Mux_h
    port map (
            O => \N__16466\,
            I => \N__16463\
        );

    \I__3450\ : Odrv4
    port map (
            O => \N__16463\,
            I => measured_delay_tr_1
        );

    \I__3449\ : CascadeMux
    port map (
            O => \N__16460\,
            I => \N__16457\
        );

    \I__3448\ : InMux
    port map (
            O => \N__16457\,
            I => \N__16453\
        );

    \I__3447\ : InMux
    port map (
            O => \N__16456\,
            I => \N__16450\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__16453\,
            I => \N__16446\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__16450\,
            I => \N__16443\
        );

    \I__3444\ : InMux
    port map (
            O => \N__16449\,
            I => \N__16440\
        );

    \I__3443\ : Span4Mux_h
    port map (
            O => \N__16446\,
            I => \N__16437\
        );

    \I__3442\ : Span4Mux_h
    port map (
            O => \N__16443\,
            I => \N__16432\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__16440\,
            I => \N__16432\
        );

    \I__3440\ : Span4Mux_h
    port map (
            O => \N__16437\,
            I => \N__16429\
        );

    \I__3439\ : Span4Mux_h
    port map (
            O => \N__16432\,
            I => \N__16426\
        );

    \I__3438\ : Odrv4
    port map (
            O => \N__16429\,
            I => measured_delay_tr_2
        );

    \I__3437\ : Odrv4
    port map (
            O => \N__16426\,
            I => measured_delay_tr_2
        );

    \I__3436\ : CascadeMux
    port map (
            O => \N__16421\,
            I => \N__16417\
        );

    \I__3435\ : CascadeMux
    port map (
            O => \N__16420\,
            I => \N__16414\
        );

    \I__3434\ : InMux
    port map (
            O => \N__16417\,
            I => \N__16411\
        );

    \I__3433\ : InMux
    port map (
            O => \N__16414\,
            I => \N__16408\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__16411\,
            I => \N__16405\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__16408\,
            I => \N__16402\
        );

    \I__3430\ : Span4Mux_h
    port map (
            O => \N__16405\,
            I => \N__16398\
        );

    \I__3429\ : Span4Mux_h
    port map (
            O => \N__16402\,
            I => \N__16395\
        );

    \I__3428\ : InMux
    port map (
            O => \N__16401\,
            I => \N__16392\
        );

    \I__3427\ : Span4Mux_h
    port map (
            O => \N__16398\,
            I => \N__16389\
        );

    \I__3426\ : Span4Mux_h
    port map (
            O => \N__16395\,
            I => \N__16386\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__16392\,
            I => \N__16383\
        );

    \I__3424\ : Odrv4
    port map (
            O => \N__16389\,
            I => measured_delay_tr_3
        );

    \I__3423\ : Odrv4
    port map (
            O => \N__16386\,
            I => measured_delay_tr_3
        );

    \I__3422\ : Odrv4
    port map (
            O => \N__16383\,
            I => measured_delay_tr_3
        );

    \I__3421\ : CascadeMux
    port map (
            O => \N__16376\,
            I => \N__16371\
        );

    \I__3420\ : CascadeMux
    port map (
            O => \N__16375\,
            I => \N__16368\
        );

    \I__3419\ : InMux
    port map (
            O => \N__16374\,
            I => \N__16365\
        );

    \I__3418\ : InMux
    port map (
            O => \N__16371\,
            I => \N__16360\
        );

    \I__3417\ : InMux
    port map (
            O => \N__16368\,
            I => \N__16360\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__16365\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__16360\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__3414\ : InMux
    port map (
            O => \N__16355\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__3413\ : CascadeMux
    port map (
            O => \N__16352\,
            I => \N__16347\
        );

    \I__3412\ : CascadeMux
    port map (
            O => \N__16351\,
            I => \N__16344\
        );

    \I__3411\ : InMux
    port map (
            O => \N__16350\,
            I => \N__16341\
        );

    \I__3410\ : InMux
    port map (
            O => \N__16347\,
            I => \N__16336\
        );

    \I__3409\ : InMux
    port map (
            O => \N__16344\,
            I => \N__16336\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__16341\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__16336\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__3406\ : InMux
    port map (
            O => \N__16331\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__3405\ : InMux
    port map (
            O => \N__16328\,
            I => \N__16323\
        );

    \I__3404\ : InMux
    port map (
            O => \N__16327\,
            I => \N__16320\
        );

    \I__3403\ : InMux
    port map (
            O => \N__16326\,
            I => \N__16317\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__16323\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__16320\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__16317\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__3399\ : InMux
    port map (
            O => \N__16310\,
            I => \bfn_9_16_0_\
        );

    \I__3398\ : InMux
    port map (
            O => \N__16307\,
            I => \N__16302\
        );

    \I__3397\ : InMux
    port map (
            O => \N__16306\,
            I => \N__16299\
        );

    \I__3396\ : InMux
    port map (
            O => \N__16305\,
            I => \N__16296\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__16302\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__16299\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__16296\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__3392\ : InMux
    port map (
            O => \N__16289\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__3391\ : InMux
    port map (
            O => \N__16286\,
            I => \N__16282\
        );

    \I__3390\ : InMux
    port map (
            O => \N__16285\,
            I => \N__16279\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__16282\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__16279\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__3387\ : CascadeMux
    port map (
            O => \N__16274\,
            I => \N__16269\
        );

    \I__3386\ : CascadeMux
    port map (
            O => \N__16273\,
            I => \N__16266\
        );

    \I__3385\ : InMux
    port map (
            O => \N__16272\,
            I => \N__16263\
        );

    \I__3384\ : InMux
    port map (
            O => \N__16269\,
            I => \N__16258\
        );

    \I__3383\ : InMux
    port map (
            O => \N__16266\,
            I => \N__16258\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__16263\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__16258\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__3380\ : InMux
    port map (
            O => \N__16253\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__3379\ : InMux
    port map (
            O => \N__16250\,
            I => \N__16246\
        );

    \I__3378\ : InMux
    port map (
            O => \N__16249\,
            I => \N__16243\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__16246\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__16243\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__3375\ : CascadeMux
    port map (
            O => \N__16238\,
            I => \N__16233\
        );

    \I__3374\ : CascadeMux
    port map (
            O => \N__16237\,
            I => \N__16230\
        );

    \I__3373\ : InMux
    port map (
            O => \N__16236\,
            I => \N__16227\
        );

    \I__3372\ : InMux
    port map (
            O => \N__16233\,
            I => \N__16222\
        );

    \I__3371\ : InMux
    port map (
            O => \N__16230\,
            I => \N__16222\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__16227\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__16222\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__3368\ : InMux
    port map (
            O => \N__16217\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__3367\ : InMux
    port map (
            O => \N__16214\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__3366\ : CascadeMux
    port map (
            O => \N__16211\,
            I => \N__16206\
        );

    \I__3365\ : CascadeMux
    port map (
            O => \N__16210\,
            I => \N__16203\
        );

    \I__3364\ : InMux
    port map (
            O => \N__16209\,
            I => \N__16200\
        );

    \I__3363\ : InMux
    port map (
            O => \N__16206\,
            I => \N__16195\
        );

    \I__3362\ : InMux
    port map (
            O => \N__16203\,
            I => \N__16195\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__16200\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__16195\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__3359\ : InMux
    port map (
            O => \N__16190\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__3358\ : CascadeMux
    port map (
            O => \N__16187\,
            I => \N__16182\
        );

    \I__3357\ : CascadeMux
    port map (
            O => \N__16186\,
            I => \N__16179\
        );

    \I__3356\ : InMux
    port map (
            O => \N__16185\,
            I => \N__16176\
        );

    \I__3355\ : InMux
    port map (
            O => \N__16182\,
            I => \N__16171\
        );

    \I__3354\ : InMux
    port map (
            O => \N__16179\,
            I => \N__16171\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__16176\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__16171\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__3351\ : InMux
    port map (
            O => \N__16166\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__3350\ : InMux
    port map (
            O => \N__16163\,
            I => \N__16158\
        );

    \I__3349\ : InMux
    port map (
            O => \N__16162\,
            I => \N__16155\
        );

    \I__3348\ : InMux
    port map (
            O => \N__16161\,
            I => \N__16152\
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__16158\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__16155\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__16152\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__3344\ : InMux
    port map (
            O => \N__16145\,
            I => \bfn_9_15_0_\
        );

    \I__3343\ : InMux
    port map (
            O => \N__16142\,
            I => \N__16137\
        );

    \I__3342\ : InMux
    port map (
            O => \N__16141\,
            I => \N__16134\
        );

    \I__3341\ : InMux
    port map (
            O => \N__16140\,
            I => \N__16131\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__16137\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__16134\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__16131\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__3337\ : InMux
    port map (
            O => \N__16124\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__3336\ : CascadeMux
    port map (
            O => \N__16121\,
            I => \N__16116\
        );

    \I__3335\ : CascadeMux
    port map (
            O => \N__16120\,
            I => \N__16113\
        );

    \I__3334\ : InMux
    port map (
            O => \N__16119\,
            I => \N__16110\
        );

    \I__3333\ : InMux
    port map (
            O => \N__16116\,
            I => \N__16105\
        );

    \I__3332\ : InMux
    port map (
            O => \N__16113\,
            I => \N__16105\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__16110\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__16105\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__3329\ : InMux
    port map (
            O => \N__16100\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__3328\ : CascadeMux
    port map (
            O => \N__16097\,
            I => \N__16092\
        );

    \I__3327\ : CascadeMux
    port map (
            O => \N__16096\,
            I => \N__16089\
        );

    \I__3326\ : InMux
    port map (
            O => \N__16095\,
            I => \N__16086\
        );

    \I__3325\ : InMux
    port map (
            O => \N__16092\,
            I => \N__16081\
        );

    \I__3324\ : InMux
    port map (
            O => \N__16089\,
            I => \N__16081\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__16086\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__16081\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__3321\ : InMux
    port map (
            O => \N__16076\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__3320\ : InMux
    port map (
            O => \N__16073\,
            I => \N__16068\
        );

    \I__3319\ : InMux
    port map (
            O => \N__16072\,
            I => \N__16063\
        );

    \I__3318\ : InMux
    port map (
            O => \N__16071\,
            I => \N__16063\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__16068\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__3316\ : LocalMux
    port map (
            O => \N__16063\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__3315\ : InMux
    port map (
            O => \N__16058\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__3314\ : InMux
    port map (
            O => \N__16055\,
            I => \N__16050\
        );

    \I__3313\ : InMux
    port map (
            O => \N__16054\,
            I => \N__16045\
        );

    \I__3312\ : InMux
    port map (
            O => \N__16053\,
            I => \N__16045\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__16050\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__16045\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__3309\ : InMux
    port map (
            O => \N__16040\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__3308\ : InMux
    port map (
            O => \N__16037\,
            I => \N__16032\
        );

    \I__3307\ : InMux
    port map (
            O => \N__16036\,
            I => \N__16027\
        );

    \I__3306\ : InMux
    port map (
            O => \N__16035\,
            I => \N__16027\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__16032\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__16027\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__3303\ : InMux
    port map (
            O => \N__16022\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__3302\ : CascadeMux
    port map (
            O => \N__16019\,
            I => \N__16014\
        );

    \I__3301\ : CascadeMux
    port map (
            O => \N__16018\,
            I => \N__16011\
        );

    \I__3300\ : InMux
    port map (
            O => \N__16017\,
            I => \N__16008\
        );

    \I__3299\ : InMux
    port map (
            O => \N__16014\,
            I => \N__16003\
        );

    \I__3298\ : InMux
    port map (
            O => \N__16011\,
            I => \N__16003\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__16008\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__16003\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__3295\ : InMux
    port map (
            O => \N__15998\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__3294\ : CascadeMux
    port map (
            O => \N__15995\,
            I => \N__15990\
        );

    \I__3293\ : CascadeMux
    port map (
            O => \N__15994\,
            I => \N__15987\
        );

    \I__3292\ : InMux
    port map (
            O => \N__15993\,
            I => \N__15984\
        );

    \I__3291\ : InMux
    port map (
            O => \N__15990\,
            I => \N__15979\
        );

    \I__3290\ : InMux
    port map (
            O => \N__15987\,
            I => \N__15979\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__15984\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__15979\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__3287\ : InMux
    port map (
            O => \N__15974\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__3286\ : InMux
    port map (
            O => \N__15971\,
            I => \N__15966\
        );

    \I__3285\ : InMux
    port map (
            O => \N__15970\,
            I => \N__15963\
        );

    \I__3284\ : InMux
    port map (
            O => \N__15969\,
            I => \N__15960\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__15966\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__15963\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__15960\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__3280\ : InMux
    port map (
            O => \N__15953\,
            I => \bfn_9_14_0_\
        );

    \I__3279\ : InMux
    port map (
            O => \N__15950\,
            I => \N__15945\
        );

    \I__3278\ : InMux
    port map (
            O => \N__15949\,
            I => \N__15942\
        );

    \I__3277\ : InMux
    port map (
            O => \N__15948\,
            I => \N__15939\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__15945\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__15942\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__15939\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__3273\ : InMux
    port map (
            O => \N__15932\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__3272\ : CascadeMux
    port map (
            O => \N__15929\,
            I => \N__15924\
        );

    \I__3271\ : CascadeMux
    port map (
            O => \N__15928\,
            I => \N__15921\
        );

    \I__3270\ : InMux
    port map (
            O => \N__15927\,
            I => \N__15918\
        );

    \I__3269\ : InMux
    port map (
            O => \N__15924\,
            I => \N__15913\
        );

    \I__3268\ : InMux
    port map (
            O => \N__15921\,
            I => \N__15913\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__15918\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__15913\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__3265\ : InMux
    port map (
            O => \N__15908\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__3264\ : CascadeMux
    port map (
            O => \N__15905\,
            I => \N__15900\
        );

    \I__3263\ : CascadeMux
    port map (
            O => \N__15904\,
            I => \N__15897\
        );

    \I__3262\ : InMux
    port map (
            O => \N__15903\,
            I => \N__15894\
        );

    \I__3261\ : InMux
    port map (
            O => \N__15900\,
            I => \N__15889\
        );

    \I__3260\ : InMux
    port map (
            O => \N__15897\,
            I => \N__15889\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__15894\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__15889\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__3257\ : InMux
    port map (
            O => \N__15884\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__3256\ : InMux
    port map (
            O => \N__15881\,
            I => \N__15876\
        );

    \I__3255\ : InMux
    port map (
            O => \N__15880\,
            I => \N__15871\
        );

    \I__3254\ : InMux
    port map (
            O => \N__15879\,
            I => \N__15871\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__15876\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__15871\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__3251\ : InMux
    port map (
            O => \N__15866\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__3250\ : InMux
    port map (
            O => \N__15863\,
            I => \N__15858\
        );

    \I__3249\ : InMux
    port map (
            O => \N__15862\,
            I => \N__15853\
        );

    \I__3248\ : InMux
    port map (
            O => \N__15861\,
            I => \N__15853\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__15858\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__15853\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__3245\ : InMux
    port map (
            O => \N__15848\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__3244\ : InMux
    port map (
            O => \N__15845\,
            I => \N__15836\
        );

    \I__3243\ : InMux
    port map (
            O => \N__15844\,
            I => \N__15836\
        );

    \I__3242\ : InMux
    port map (
            O => \N__15843\,
            I => \N__15836\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__15836\,
            I => \delay_measurement_inst.N_243\
        );

    \I__3240\ : InMux
    port map (
            O => \N__15833\,
            I => \N__15816\
        );

    \I__3239\ : InMux
    port map (
            O => \N__15832\,
            I => \N__15816\
        );

    \I__3238\ : InMux
    port map (
            O => \N__15831\,
            I => \N__15816\
        );

    \I__3237\ : InMux
    port map (
            O => \N__15830\,
            I => \N__15816\
        );

    \I__3236\ : InMux
    port map (
            O => \N__15829\,
            I => \N__15816\
        );

    \I__3235\ : InMux
    port map (
            O => \N__15828\,
            I => \N__15813\
        );

    \I__3234\ : InMux
    port map (
            O => \N__15827\,
            I => \N__15810\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__15816\,
            I => \delay_measurement_inst.N_247\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__15813\,
            I => \delay_measurement_inst.N_247\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__15810\,
            I => \delay_measurement_inst.N_247\
        );

    \I__3230\ : InMux
    port map (
            O => \N__15803\,
            I => \N__15791\
        );

    \I__3229\ : InMux
    port map (
            O => \N__15802\,
            I => \N__15791\
        );

    \I__3228\ : InMux
    port map (
            O => \N__15801\,
            I => \N__15791\
        );

    \I__3227\ : InMux
    port map (
            O => \N__15800\,
            I => \N__15786\
        );

    \I__3226\ : InMux
    port map (
            O => \N__15799\,
            I => \N__15786\
        );

    \I__3225\ : InMux
    port map (
            O => \N__15798\,
            I => \N__15783\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__15791\,
            I => \delay_measurement_inst.N_216_1\
        );

    \I__3223\ : LocalMux
    port map (
            O => \N__15786\,
            I => \delay_measurement_inst.N_216_1\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__15783\,
            I => \delay_measurement_inst.N_216_1\
        );

    \I__3221\ : InMux
    port map (
            O => \N__15776\,
            I => \N__15773\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__15773\,
            I => \N__15768\
        );

    \I__3219\ : InMux
    port map (
            O => \N__15772\,
            I => \N__15765\
        );

    \I__3218\ : CascadeMux
    port map (
            O => \N__15771\,
            I => \N__15762\
        );

    \I__3217\ : Span4Mux_v
    port map (
            O => \N__15768\,
            I => \N__15759\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__15765\,
            I => \N__15756\
        );

    \I__3215\ : InMux
    port map (
            O => \N__15762\,
            I => \N__15753\
        );

    \I__3214\ : Span4Mux_v
    port map (
            O => \N__15759\,
            I => \N__15746\
        );

    \I__3213\ : Span4Mux_v
    port map (
            O => \N__15756\,
            I => \N__15746\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__15753\,
            I => \N__15746\
        );

    \I__3211\ : Span4Mux_h
    port map (
            O => \N__15746\,
            I => \N__15743\
        );

    \I__3210\ : Odrv4
    port map (
            O => \N__15743\,
            I => measured_delay_hc_13
        );

    \I__3209\ : CEMux
    port map (
            O => \N__15740\,
            I => \N__15736\
        );

    \I__3208\ : CEMux
    port map (
            O => \N__15739\,
            I => \N__15733\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__15736\,
            I => \N__15729\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__15733\,
            I => \N__15726\
        );

    \I__3205\ : CEMux
    port map (
            O => \N__15732\,
            I => \N__15723\
        );

    \I__3204\ : Span4Mux_v
    port map (
            O => \N__15729\,
            I => \N__15720\
        );

    \I__3203\ : Span4Mux_h
    port map (
            O => \N__15726\,
            I => \N__15717\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__15723\,
            I => \N__15714\
        );

    \I__3201\ : Odrv4
    port map (
            O => \N__15720\,
            I => \delay_measurement_inst.un3_elapsed_time_hc_0_i_0\
        );

    \I__3200\ : Odrv4
    port map (
            O => \N__15717\,
            I => \delay_measurement_inst.un3_elapsed_time_hc_0_i_0\
        );

    \I__3199\ : Odrv4
    port map (
            O => \N__15714\,
            I => \delay_measurement_inst.un3_elapsed_time_hc_0_i_0\
        );

    \I__3198\ : CascadeMux
    port map (
            O => \N__15707\,
            I => \N__15703\
        );

    \I__3197\ : InMux
    port map (
            O => \N__15706\,
            I => \N__15700\
        );

    \I__3196\ : InMux
    port map (
            O => \N__15703\,
            I => \N__15696\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__15700\,
            I => \N__15692\
        );

    \I__3194\ : InMux
    port map (
            O => \N__15699\,
            I => \N__15689\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__15696\,
            I => \N__15686\
        );

    \I__3192\ : InMux
    port map (
            O => \N__15695\,
            I => \N__15683\
        );

    \I__3191\ : Span4Mux_h
    port map (
            O => \N__15692\,
            I => \N__15678\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__15689\,
            I => \N__15678\
        );

    \I__3189\ : Odrv4
    port map (
            O => \N__15686\,
            I => \phase_controller_slave.stateZ0Z_1\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__15683\,
            I => \phase_controller_slave.stateZ0Z_1\
        );

    \I__3187\ : Odrv4
    port map (
            O => \N__15678\,
            I => \phase_controller_slave.stateZ0Z_1\
        );

    \I__3186\ : IoInMux
    port map (
            O => \N__15671\,
            I => \N__15668\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__15668\,
            I => \N__15665\
        );

    \I__3184\ : Odrv12
    port map (
            O => \N__15665\,
            I => s4_phy_c
        );

    \I__3183\ : InMux
    port map (
            O => \N__15662\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__3182\ : CascadeMux
    port map (
            O => \N__15659\,
            I => \N__15654\
        );

    \I__3181\ : CascadeMux
    port map (
            O => \N__15658\,
            I => \N__15651\
        );

    \I__3180\ : InMux
    port map (
            O => \N__15657\,
            I => \N__15648\
        );

    \I__3179\ : InMux
    port map (
            O => \N__15654\,
            I => \N__15643\
        );

    \I__3178\ : InMux
    port map (
            O => \N__15651\,
            I => \N__15643\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__15648\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__15643\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__3175\ : InMux
    port map (
            O => \N__15638\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__3174\ : CascadeMux
    port map (
            O => \N__15635\,
            I => \N__15630\
        );

    \I__3173\ : CascadeMux
    port map (
            O => \N__15634\,
            I => \N__15627\
        );

    \I__3172\ : InMux
    port map (
            O => \N__15633\,
            I => \N__15624\
        );

    \I__3171\ : InMux
    port map (
            O => \N__15630\,
            I => \N__15619\
        );

    \I__3170\ : InMux
    port map (
            O => \N__15627\,
            I => \N__15619\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__15624\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__15619\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__3167\ : InMux
    port map (
            O => \N__15614\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__3166\ : InMux
    port map (
            O => \N__15611\,
            I => \N__15606\
        );

    \I__3165\ : InMux
    port map (
            O => \N__15610\,
            I => \N__15601\
        );

    \I__3164\ : InMux
    port map (
            O => \N__15609\,
            I => \N__15601\
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__15606\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__15601\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__3161\ : InMux
    port map (
            O => \N__15596\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__3160\ : CascadeMux
    port map (
            O => \N__15593\,
            I => \delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_3_cascade_\
        );

    \I__3159\ : InMux
    port map (
            O => \N__15590\,
            I => \N__15584\
        );

    \I__3158\ : InMux
    port map (
            O => \N__15589\,
            I => \N__15584\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__15584\,
            I => \delay_measurement_inst.delay_hc_timer.N_232_4\
        );

    \I__3156\ : InMux
    port map (
            O => \N__15581\,
            I => \N__15578\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__15578\,
            I => \delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_2\
        );

    \I__3154\ : CascadeMux
    port map (
            O => \N__15575\,
            I => \delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_6_cascade_\
        );

    \I__3153\ : InMux
    port map (
            O => \N__15572\,
            I => \N__15569\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__15569\,
            I => \delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_0_7\
        );

    \I__3151\ : InMux
    port map (
            O => \N__15566\,
            I => \N__15563\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__15563\,
            I => \delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_7\
        );

    \I__3149\ : InMux
    port map (
            O => \N__15560\,
            I => \N__15554\
        );

    \I__3148\ : InMux
    port map (
            O => \N__15559\,
            I => \N__15554\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__15554\,
            I => \delay_measurement_inst.un3_elapsed_time_hc_0_i\
        );

    \I__3146\ : CascadeMux
    port map (
            O => \N__15551\,
            I => \delay_measurement_inst.un3_elapsed_time_hc_0_i_cascade_\
        );

    \I__3145\ : InMux
    port map (
            O => \N__15548\,
            I => \N__15545\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__15545\,
            I => \delay_measurement_inst.N_219\
        );

    \I__3143\ : CascadeMux
    port map (
            O => \N__15542\,
            I => \delay_measurement_inst.delay_hc_timer.N_237_cascade_\
        );

    \I__3142\ : CascadeMux
    port map (
            O => \N__15539\,
            I => \N__15534\
        );

    \I__3141\ : InMux
    port map (
            O => \N__15538\,
            I => \N__15524\
        );

    \I__3140\ : InMux
    port map (
            O => \N__15537\,
            I => \N__15524\
        );

    \I__3139\ : InMux
    port map (
            O => \N__15534\,
            I => \N__15517\
        );

    \I__3138\ : InMux
    port map (
            O => \N__15533\,
            I => \N__15517\
        );

    \I__3137\ : InMux
    port map (
            O => \N__15532\,
            I => \N__15517\
        );

    \I__3136\ : InMux
    port map (
            O => \N__15531\,
            I => \N__15512\
        );

    \I__3135\ : InMux
    port map (
            O => \N__15530\,
            I => \N__15512\
        );

    \I__3134\ : InMux
    port map (
            O => \N__15529\,
            I => \N__15509\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__15524\,
            I => \delay_measurement_inst.N_209\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__15517\,
            I => \delay_measurement_inst.N_209\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__15512\,
            I => \delay_measurement_inst.N_209\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__15509\,
            I => \delay_measurement_inst.N_209\
        );

    \I__3129\ : InMux
    port map (
            O => \N__15500\,
            I => \N__15495\
        );

    \I__3128\ : InMux
    port map (
            O => \N__15499\,
            I => \N__15492\
        );

    \I__3127\ : InMux
    port map (
            O => \N__15498\,
            I => \N__15489\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__15495\,
            I => \delay_measurement_inst.N_207\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__15492\,
            I => \delay_measurement_inst.N_207\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__15489\,
            I => \delay_measurement_inst.N_207\
        );

    \I__3123\ : CascadeMux
    port map (
            O => \N__15482\,
            I => \delay_measurement_inst.N_207_cascade_\
        );

    \I__3122\ : CascadeMux
    port map (
            O => \N__15479\,
            I => \N__15475\
        );

    \I__3121\ : CascadeMux
    port map (
            O => \N__15478\,
            I => \N__15472\
        );

    \I__3120\ : InMux
    port map (
            O => \N__15475\,
            I => \N__15463\
        );

    \I__3119\ : InMux
    port map (
            O => \N__15472\,
            I => \N__15460\
        );

    \I__3118\ : InMux
    port map (
            O => \N__15471\,
            I => \N__15440\
        );

    \I__3117\ : InMux
    port map (
            O => \N__15470\,
            I => \N__15440\
        );

    \I__3116\ : InMux
    port map (
            O => \N__15469\,
            I => \N__15440\
        );

    \I__3115\ : InMux
    port map (
            O => \N__15468\,
            I => \N__15440\
        );

    \I__3114\ : InMux
    port map (
            O => \N__15467\,
            I => \N__15440\
        );

    \I__3113\ : InMux
    port map (
            O => \N__15466\,
            I => \N__15437\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__15463\,
            I => \N__15429\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__15460\,
            I => \N__15426\
        );

    \I__3110\ : InMux
    port map (
            O => \N__15459\,
            I => \N__15421\
        );

    \I__3109\ : InMux
    port map (
            O => \N__15458\,
            I => \N__15421\
        );

    \I__3108\ : InMux
    port map (
            O => \N__15457\,
            I => \N__15405\
        );

    \I__3107\ : InMux
    port map (
            O => \N__15456\,
            I => \N__15405\
        );

    \I__3106\ : InMux
    port map (
            O => \N__15455\,
            I => \N__15405\
        );

    \I__3105\ : InMux
    port map (
            O => \N__15454\,
            I => \N__15405\
        );

    \I__3104\ : InMux
    port map (
            O => \N__15453\,
            I => \N__15405\
        );

    \I__3103\ : InMux
    port map (
            O => \N__15452\,
            I => \N__15405\
        );

    \I__3102\ : InMux
    port map (
            O => \N__15451\,
            I => \N__15405\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__15440\,
            I => \N__15402\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__15437\,
            I => \N__15399\
        );

    \I__3099\ : InMux
    port map (
            O => \N__15436\,
            I => \N__15395\
        );

    \I__3098\ : InMux
    port map (
            O => \N__15435\,
            I => \N__15392\
        );

    \I__3097\ : InMux
    port map (
            O => \N__15434\,
            I => \N__15385\
        );

    \I__3096\ : InMux
    port map (
            O => \N__15433\,
            I => \N__15385\
        );

    \I__3095\ : InMux
    port map (
            O => \N__15432\,
            I => \N__15385\
        );

    \I__3094\ : Span4Mux_h
    port map (
            O => \N__15429\,
            I => \N__15382\
        );

    \I__3093\ : Sp12to4
    port map (
            O => \N__15426\,
            I => \N__15377\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__15421\,
            I => \N__15377\
        );

    \I__3091\ : InMux
    port map (
            O => \N__15420\,
            I => \N__15374\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__15405\,
            I => \N__15367\
        );

    \I__3089\ : Span4Mux_h
    port map (
            O => \N__15402\,
            I => \N__15367\
        );

    \I__3088\ : Span4Mux_h
    port map (
            O => \N__15399\,
            I => \N__15367\
        );

    \I__3087\ : InMux
    port map (
            O => \N__15398\,
            I => \N__15364\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__15395\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__15392\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__15385\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__3083\ : Odrv4
    port map (
            O => \N__15382\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__3082\ : Odrv12
    port map (
            O => \N__15377\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__15374\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__3080\ : Odrv4
    port map (
            O => \N__15367\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__15364\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__3078\ : CascadeMux
    port map (
            O => \N__15347\,
            I => \N__15338\
        );

    \I__3077\ : CascadeMux
    port map (
            O => \N__15346\,
            I => \N__15331\
        );

    \I__3076\ : CascadeMux
    port map (
            O => \N__15345\,
            I => \N__15327\
        );

    \I__3075\ : CascadeMux
    port map (
            O => \N__15344\,
            I => \N__15324\
        );

    \I__3074\ : CascadeMux
    port map (
            O => \N__15343\,
            I => \N__15321\
        );

    \I__3073\ : CascadeMux
    port map (
            O => \N__15342\,
            I => \N__15313\
        );

    \I__3072\ : CascadeMux
    port map (
            O => \N__15341\,
            I => \N__15310\
        );

    \I__3071\ : InMux
    port map (
            O => \N__15338\,
            I => \N__15307\
        );

    \I__3070\ : CascadeMux
    port map (
            O => \N__15337\,
            I => \N__15300\
        );

    \I__3069\ : CascadeMux
    port map (
            O => \N__15336\,
            I => \N__15297\
        );

    \I__3068\ : CascadeMux
    port map (
            O => \N__15335\,
            I => \N__15294\
        );

    \I__3067\ : CascadeMux
    port map (
            O => \N__15334\,
            I => \N__15291\
        );

    \I__3066\ : InMux
    port map (
            O => \N__15331\,
            I => \N__15286\
        );

    \I__3065\ : InMux
    port map (
            O => \N__15330\,
            I => \N__15286\
        );

    \I__3064\ : InMux
    port map (
            O => \N__15327\,
            I => \N__15282\
        );

    \I__3063\ : InMux
    port map (
            O => \N__15324\,
            I => \N__15275\
        );

    \I__3062\ : InMux
    port map (
            O => \N__15321\,
            I => \N__15275\
        );

    \I__3061\ : InMux
    port map (
            O => \N__15320\,
            I => \N__15275\
        );

    \I__3060\ : InMux
    port map (
            O => \N__15319\,
            I => \N__15262\
        );

    \I__3059\ : InMux
    port map (
            O => \N__15318\,
            I => \N__15262\
        );

    \I__3058\ : InMux
    port map (
            O => \N__15317\,
            I => \N__15262\
        );

    \I__3057\ : InMux
    port map (
            O => \N__15316\,
            I => \N__15262\
        );

    \I__3056\ : InMux
    port map (
            O => \N__15313\,
            I => \N__15262\
        );

    \I__3055\ : InMux
    port map (
            O => \N__15310\,
            I => \N__15262\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__15307\,
            I => \N__15259\
        );

    \I__3053\ : InMux
    port map (
            O => \N__15306\,
            I => \N__15242\
        );

    \I__3052\ : InMux
    port map (
            O => \N__15305\,
            I => \N__15242\
        );

    \I__3051\ : InMux
    port map (
            O => \N__15304\,
            I => \N__15242\
        );

    \I__3050\ : InMux
    port map (
            O => \N__15303\,
            I => \N__15242\
        );

    \I__3049\ : InMux
    port map (
            O => \N__15300\,
            I => \N__15242\
        );

    \I__3048\ : InMux
    port map (
            O => \N__15297\,
            I => \N__15242\
        );

    \I__3047\ : InMux
    port map (
            O => \N__15294\,
            I => \N__15242\
        );

    \I__3046\ : InMux
    port map (
            O => \N__15291\,
            I => \N__15242\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__15286\,
            I => \N__15239\
        );

    \I__3044\ : InMux
    port map (
            O => \N__15285\,
            I => \N__15236\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__15282\,
            I => \N__15230\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__15275\,
            I => \N__15230\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__15262\,
            I => \N__15227\
        );

    \I__3040\ : Span4Mux_v
    port map (
            O => \N__15259\,
            I => \N__15222\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__15242\,
            I => \N__15222\
        );

    \I__3038\ : Span4Mux_h
    port map (
            O => \N__15239\,
            I => \N__15218\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__15236\,
            I => \N__15215\
        );

    \I__3036\ : InMux
    port map (
            O => \N__15235\,
            I => \N__15212\
        );

    \I__3035\ : Span4Mux_v
    port map (
            O => \N__15230\,
            I => \N__15209\
        );

    \I__3034\ : Span4Mux_v
    port map (
            O => \N__15227\,
            I => \N__15204\
        );

    \I__3033\ : Span4Mux_h
    port map (
            O => \N__15222\,
            I => \N__15204\
        );

    \I__3032\ : InMux
    port map (
            O => \N__15221\,
            I => \N__15201\
        );

    \I__3031\ : Span4Mux_v
    port map (
            O => \N__15218\,
            I => \N__15196\
        );

    \I__3030\ : Span4Mux_h
    port map (
            O => \N__15215\,
            I => \N__15196\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__15212\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__3028\ : Odrv4
    port map (
            O => \N__15209\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__3027\ : Odrv4
    port map (
            O => \N__15204\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__15201\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__3025\ : Odrv4
    port map (
            O => \N__15196\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__3024\ : InMux
    port map (
            O => \N__15185\,
            I => \N__15181\
        );

    \I__3023\ : InMux
    port map (
            O => \N__15184\,
            I => \N__15178\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__15181\,
            I => \N__15172\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__15178\,
            I => \N__15172\
        );

    \I__3020\ : InMux
    port map (
            O => \N__15177\,
            I => \N__15169\
        );

    \I__3019\ : Span4Mux_h
    port map (
            O => \N__15172\,
            I => \N__15164\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__15169\,
            I => \N__15161\
        );

    \I__3017\ : InMux
    port map (
            O => \N__15168\,
            I => \N__15156\
        );

    \I__3016\ : InMux
    port map (
            O => \N__15167\,
            I => \N__15156\
        );

    \I__3015\ : Odrv4
    port map (
            O => \N__15164\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__3014\ : Odrv4
    port map (
            O => \N__15161\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__15156\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__3012\ : CascadeMux
    port map (
            O => \N__15149\,
            I => \N__15137\
        );

    \I__3011\ : InMux
    port map (
            O => \N__15148\,
            I => \N__15124\
        );

    \I__3010\ : InMux
    port map (
            O => \N__15147\,
            I => \N__15124\
        );

    \I__3009\ : InMux
    port map (
            O => \N__15146\,
            I => \N__15111\
        );

    \I__3008\ : InMux
    port map (
            O => \N__15145\,
            I => \N__15111\
        );

    \I__3007\ : InMux
    port map (
            O => \N__15144\,
            I => \N__15111\
        );

    \I__3006\ : InMux
    port map (
            O => \N__15143\,
            I => \N__15111\
        );

    \I__3005\ : InMux
    port map (
            O => \N__15142\,
            I => \N__15111\
        );

    \I__3004\ : InMux
    port map (
            O => \N__15141\,
            I => \N__15111\
        );

    \I__3003\ : InMux
    port map (
            O => \N__15140\,
            I => \N__15108\
        );

    \I__3002\ : InMux
    port map (
            O => \N__15137\,
            I => \N__15100\
        );

    \I__3001\ : InMux
    port map (
            O => \N__15136\,
            I => \N__15083\
        );

    \I__3000\ : InMux
    port map (
            O => \N__15135\,
            I => \N__15083\
        );

    \I__2999\ : InMux
    port map (
            O => \N__15134\,
            I => \N__15083\
        );

    \I__2998\ : InMux
    port map (
            O => \N__15133\,
            I => \N__15083\
        );

    \I__2997\ : InMux
    port map (
            O => \N__15132\,
            I => \N__15083\
        );

    \I__2996\ : InMux
    port map (
            O => \N__15131\,
            I => \N__15083\
        );

    \I__2995\ : InMux
    port map (
            O => \N__15130\,
            I => \N__15083\
        );

    \I__2994\ : InMux
    port map (
            O => \N__15129\,
            I => \N__15083\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__15124\,
            I => \N__15078\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__15111\,
            I => \N__15078\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__15108\,
            I => \N__15075\
        );

    \I__2990\ : InMux
    port map (
            O => \N__15107\,
            I => \N__15071\
        );

    \I__2989\ : InMux
    port map (
            O => \N__15106\,
            I => \N__15068\
        );

    \I__2988\ : InMux
    port map (
            O => \N__15105\,
            I => \N__15063\
        );

    \I__2987\ : InMux
    port map (
            O => \N__15104\,
            I => \N__15063\
        );

    \I__2986\ : InMux
    port map (
            O => \N__15103\,
            I => \N__15060\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__15100\,
            I => \N__15051\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__15083\,
            I => \N__15051\
        );

    \I__2983\ : Span4Mux_h
    port map (
            O => \N__15078\,
            I => \N__15051\
        );

    \I__2982\ : Span4Mux_h
    port map (
            O => \N__15075\,
            I => \N__15051\
        );

    \I__2981\ : InMux
    port map (
            O => \N__15074\,
            I => \N__15048\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__15071\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__15068\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__15063\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__15060\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__2976\ : Odrv4
    port map (
            O => \N__15051\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__15048\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__2974\ : CascadeMux
    port map (
            O => \N__15035\,
            I => \N__15031\
        );

    \I__2973\ : CascadeMux
    port map (
            O => \N__15034\,
            I => \N__15028\
        );

    \I__2972\ : InMux
    port map (
            O => \N__15031\,
            I => \N__15025\
        );

    \I__2971\ : InMux
    port map (
            O => \N__15028\,
            I => \N__15022\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__15025\,
            I => \delay_measurement_inst.elapsed_time_hc_1\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__15022\,
            I => \delay_measurement_inst.elapsed_time_hc_1\
        );

    \I__2968\ : CascadeMux
    port map (
            O => \N__15017\,
            I => \N__15014\
        );

    \I__2967\ : InMux
    port map (
            O => \N__15014\,
            I => \N__15011\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__15011\,
            I => \delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_0_4\
        );

    \I__2965\ : InMux
    port map (
            O => \N__15008\,
            I => \N__15005\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__15005\,
            I => \delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_0_3\
        );

    \I__2963\ : InMux
    port map (
            O => \N__15002\,
            I => \N__14997\
        );

    \I__2962\ : InMux
    port map (
            O => \N__15001\,
            I => \N__14992\
        );

    \I__2961\ : InMux
    port map (
            O => \N__15000\,
            I => \N__14992\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__14997\,
            I => \delay_measurement_inst.elapsed_time_hc_2\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__14992\,
            I => \delay_measurement_inst.elapsed_time_hc_2\
        );

    \I__2958\ : InMux
    port map (
            O => \N__14987\,
            I => \N__14984\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__14984\,
            I => \N__14980\
        );

    \I__2956\ : InMux
    port map (
            O => \N__14983\,
            I => \N__14977\
        );

    \I__2955\ : Span4Mux_h
    port map (
            O => \N__14980\,
            I => \N__14974\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__14977\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__2953\ : Odrv4
    port map (
            O => \N__14974\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__2952\ : InMux
    port map (
            O => \N__14969\,
            I => \N__14966\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__14966\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16\
        );

    \I__2950\ : InMux
    port map (
            O => \N__14963\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14\
        );

    \I__2949\ : InMux
    port map (
            O => \N__14960\,
            I => \N__14956\
        );

    \I__2948\ : InMux
    port map (
            O => \N__14959\,
            I => \N__14953\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__14956\,
            I => \N__14950\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__14953\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__2945\ : Odrv4
    port map (
            O => \N__14950\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__2944\ : InMux
    port map (
            O => \N__14945\,
            I => \N__14942\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__14942\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17\
        );

    \I__2942\ : InMux
    port map (
            O => \N__14939\,
            I => \bfn_8_19_0_\
        );

    \I__2941\ : InMux
    port map (
            O => \N__14936\,
            I => \N__14932\
        );

    \I__2940\ : InMux
    port map (
            O => \N__14935\,
            I => \N__14929\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__14932\,
            I => \N__14926\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__14929\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__2937\ : Odrv4
    port map (
            O => \N__14926\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__2936\ : InMux
    port map (
            O => \N__14921\,
            I => \N__14918\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__14918\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18\
        );

    \I__2934\ : InMux
    port map (
            O => \N__14915\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16\
        );

    \I__2933\ : InMux
    port map (
            O => \N__14912\,
            I => \N__14908\
        );

    \I__2932\ : InMux
    port map (
            O => \N__14911\,
            I => \N__14905\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__14908\,
            I => \N__14902\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__14905\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__2929\ : Odrv4
    port map (
            O => \N__14902\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__2928\ : InMux
    port map (
            O => \N__14897\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17\
        );

    \I__2927\ : InMux
    port map (
            O => \N__14894\,
            I => \N__14891\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__14891\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19\
        );

    \I__2925\ : InMux
    port map (
            O => \N__14888\,
            I => \N__14884\
        );

    \I__2924\ : InMux
    port map (
            O => \N__14887\,
            I => \N__14881\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__14884\,
            I => \N__14876\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__14881\,
            I => \N__14873\
        );

    \I__2921\ : InMux
    port map (
            O => \N__14880\,
            I => \N__14868\
        );

    \I__2920\ : InMux
    port map (
            O => \N__14879\,
            I => \N__14868\
        );

    \I__2919\ : Span4Mux_h
    port map (
            O => \N__14876\,
            I => \N__14865\
        );

    \I__2918\ : Span4Mux_h
    port map (
            O => \N__14873\,
            I => \N__14862\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__14868\,
            I => \N__14859\
        );

    \I__2916\ : Odrv4
    port map (
            O => \N__14865\,
            I => \phase_controller_inst1.stoper_tr.N_55\
        );

    \I__2915\ : Odrv4
    port map (
            O => \N__14862\,
            I => \phase_controller_inst1.stoper_tr.N_55\
        );

    \I__2914\ : Odrv12
    port map (
            O => \N__14859\,
            I => \phase_controller_inst1.stoper_tr.N_55\
        );

    \I__2913\ : InMux
    port map (
            O => \N__14852\,
            I => \N__14849\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__14849\,
            I => \N__14843\
        );

    \I__2911\ : InMux
    port map (
            O => \N__14848\,
            I => \N__14836\
        );

    \I__2910\ : InMux
    port map (
            O => \N__14847\,
            I => \N__14836\
        );

    \I__2909\ : InMux
    port map (
            O => \N__14846\,
            I => \N__14836\
        );

    \I__2908\ : Span4Mux_v
    port map (
            O => \N__14843\,
            I => \N__14831\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__14836\,
            I => \N__14831\
        );

    \I__2906\ : Odrv4
    port map (
            O => \N__14831\,
            I => \phase_controller_slave.stoper_tr.time_passed11\
        );

    \I__2905\ : InMux
    port map (
            O => \N__14828\,
            I => \N__14816\
        );

    \I__2904\ : InMux
    port map (
            O => \N__14827\,
            I => \N__14816\
        );

    \I__2903\ : InMux
    port map (
            O => \N__14826\,
            I => \N__14816\
        );

    \I__2902\ : InMux
    port map (
            O => \N__14825\,
            I => \N__14807\
        );

    \I__2901\ : InMux
    port map (
            O => \N__14824\,
            I => \N__14807\
        );

    \I__2900\ : InMux
    port map (
            O => \N__14823\,
            I => \N__14807\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__14816\,
            I => \N__14804\
        );

    \I__2898\ : CascadeMux
    port map (
            O => \N__14815\,
            I => \N__14801\
        );

    \I__2897\ : CascadeMux
    port map (
            O => \N__14814\,
            I => \N__14795\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__14807\,
            I => \N__14791\
        );

    \I__2895\ : Span4Mux_v
    port map (
            O => \N__14804\,
            I => \N__14788\
        );

    \I__2894\ : InMux
    port map (
            O => \N__14801\,
            I => \N__14775\
        );

    \I__2893\ : InMux
    port map (
            O => \N__14800\,
            I => \N__14775\
        );

    \I__2892\ : InMux
    port map (
            O => \N__14799\,
            I => \N__14775\
        );

    \I__2891\ : InMux
    port map (
            O => \N__14798\,
            I => \N__14775\
        );

    \I__2890\ : InMux
    port map (
            O => \N__14795\,
            I => \N__14775\
        );

    \I__2889\ : InMux
    port map (
            O => \N__14794\,
            I => \N__14775\
        );

    \I__2888\ : Span4Mux_v
    port map (
            O => \N__14791\,
            I => \N__14772\
        );

    \I__2887\ : Span4Mux_h
    port map (
            O => \N__14788\,
            I => \N__14769\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__14775\,
            I => \N__14766\
        );

    \I__2885\ : Odrv4
    port map (
            O => \N__14772\,
            I => \phase_controller_inst1.stoper_tr.N_50\
        );

    \I__2884\ : Odrv4
    port map (
            O => \N__14769\,
            I => \phase_controller_inst1.stoper_tr.N_50\
        );

    \I__2883\ : Odrv12
    port map (
            O => \N__14766\,
            I => \phase_controller_inst1.stoper_tr.N_50\
        );

    \I__2882\ : InMux
    port map (
            O => \N__14759\,
            I => \N__14751\
        );

    \I__2881\ : InMux
    port map (
            O => \N__14758\,
            I => \N__14751\
        );

    \I__2880\ : InMux
    port map (
            O => \N__14757\,
            I => \N__14746\
        );

    \I__2879\ : InMux
    port map (
            O => \N__14756\,
            I => \N__14746\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__14751\,
            I => \N__14742\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__14746\,
            I => \N__14739\
        );

    \I__2876\ : InMux
    port map (
            O => \N__14745\,
            I => \N__14736\
        );

    \I__2875\ : Span4Mux_v
    port map (
            O => \N__14742\,
            I => \N__14729\
        );

    \I__2874\ : Span4Mux_v
    port map (
            O => \N__14739\,
            I => \N__14729\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__14736\,
            I => \N__14729\
        );

    \I__2872\ : Odrv4
    port map (
            O => \N__14729\,
            I => \phase_controller_inst1.stoper_tr.N_32\
        );

    \I__2871\ : CascadeMux
    port map (
            O => \N__14726\,
            I => \phase_controller_inst1.stoper_tr.N_32_cascade_\
        );

    \I__2870\ : InMux
    port map (
            O => \N__14723\,
            I => \N__14709\
        );

    \I__2869\ : InMux
    port map (
            O => \N__14722\,
            I => \N__14709\
        );

    \I__2868\ : InMux
    port map (
            O => \N__14721\,
            I => \N__14709\
        );

    \I__2867\ : InMux
    port map (
            O => \N__14720\,
            I => \N__14698\
        );

    \I__2866\ : InMux
    port map (
            O => \N__14719\,
            I => \N__14698\
        );

    \I__2865\ : InMux
    port map (
            O => \N__14718\,
            I => \N__14698\
        );

    \I__2864\ : InMux
    port map (
            O => \N__14717\,
            I => \N__14698\
        );

    \I__2863\ : InMux
    port map (
            O => \N__14716\,
            I => \N__14698\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__14709\,
            I => \N__14687\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__14698\,
            I => \N__14684\
        );

    \I__2860\ : InMux
    port map (
            O => \N__14697\,
            I => \N__14667\
        );

    \I__2859\ : InMux
    port map (
            O => \N__14696\,
            I => \N__14667\
        );

    \I__2858\ : InMux
    port map (
            O => \N__14695\,
            I => \N__14667\
        );

    \I__2857\ : InMux
    port map (
            O => \N__14694\,
            I => \N__14667\
        );

    \I__2856\ : InMux
    port map (
            O => \N__14693\,
            I => \N__14667\
        );

    \I__2855\ : InMux
    port map (
            O => \N__14692\,
            I => \N__14667\
        );

    \I__2854\ : InMux
    port map (
            O => \N__14691\,
            I => \N__14667\
        );

    \I__2853\ : InMux
    port map (
            O => \N__14690\,
            I => \N__14667\
        );

    \I__2852\ : Span4Mux_h
    port map (
            O => \N__14687\,
            I => \N__14664\
        );

    \I__2851\ : Span4Mux_h
    port map (
            O => \N__14684\,
            I => \N__14661\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__14667\,
            I => \N__14658\
        );

    \I__2849\ : Odrv4
    port map (
            O => \N__14664\,
            I => \phase_controller_inst1.stoper_tr.N_33\
        );

    \I__2848\ : Odrv4
    port map (
            O => \N__14661\,
            I => \phase_controller_inst1.stoper_tr.N_33\
        );

    \I__2847\ : Odrv12
    port map (
            O => \N__14658\,
            I => \phase_controller_inst1.stoper_tr.N_33\
        );

    \I__2846\ : InMux
    port map (
            O => \N__14651\,
            I => \N__14647\
        );

    \I__2845\ : InMux
    port map (
            O => \N__14650\,
            I => \N__14644\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__14647\,
            I => \N__14641\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__14644\,
            I => \N__14636\
        );

    \I__2842\ : Span4Mux_h
    port map (
            O => \N__14641\,
            I => \N__14636\
        );

    \I__2841\ : Odrv4
    port map (
            O => \N__14636\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__2840\ : CascadeMux
    port map (
            O => \N__14633\,
            I => \N__14630\
        );

    \I__2839\ : InMux
    port map (
            O => \N__14630\,
            I => \N__14627\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__14627\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8\
        );

    \I__2837\ : InMux
    port map (
            O => \N__14624\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6\
        );

    \I__2836\ : InMux
    port map (
            O => \N__14621\,
            I => \N__14617\
        );

    \I__2835\ : InMux
    port map (
            O => \N__14620\,
            I => \N__14614\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__14617\,
            I => \N__14611\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__14614\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__2832\ : Odrv4
    port map (
            O => \N__14611\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__2831\ : InMux
    port map (
            O => \N__14606\,
            I => \N__14603\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__14603\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9\
        );

    \I__2829\ : InMux
    port map (
            O => \N__14600\,
            I => \bfn_8_18_0_\
        );

    \I__2828\ : InMux
    port map (
            O => \N__14597\,
            I => \N__14593\
        );

    \I__2827\ : InMux
    port map (
            O => \N__14596\,
            I => \N__14590\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__14593\,
            I => \N__14587\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__14590\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__2824\ : Odrv4
    port map (
            O => \N__14587\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__2823\ : CascadeMux
    port map (
            O => \N__14582\,
            I => \N__14579\
        );

    \I__2822\ : InMux
    port map (
            O => \N__14579\,
            I => \N__14576\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__14576\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10\
        );

    \I__2820\ : InMux
    port map (
            O => \N__14573\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8\
        );

    \I__2819\ : InMux
    port map (
            O => \N__14570\,
            I => \N__14566\
        );

    \I__2818\ : InMux
    port map (
            O => \N__14569\,
            I => \N__14563\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__14566\,
            I => \N__14560\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__14563\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__2815\ : Odrv4
    port map (
            O => \N__14560\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__2814\ : InMux
    port map (
            O => \N__14555\,
            I => \N__14552\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__14552\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11\
        );

    \I__2812\ : InMux
    port map (
            O => \N__14549\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9\
        );

    \I__2811\ : InMux
    port map (
            O => \N__14546\,
            I => \N__14543\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__14543\,
            I => \N__14539\
        );

    \I__2809\ : InMux
    port map (
            O => \N__14542\,
            I => \N__14536\
        );

    \I__2808\ : Span4Mux_h
    port map (
            O => \N__14539\,
            I => \N__14533\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__14536\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__2806\ : Odrv4
    port map (
            O => \N__14533\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__2805\ : CascadeMux
    port map (
            O => \N__14528\,
            I => \N__14525\
        );

    \I__2804\ : InMux
    port map (
            O => \N__14525\,
            I => \N__14522\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__14522\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12\
        );

    \I__2802\ : InMux
    port map (
            O => \N__14519\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10\
        );

    \I__2801\ : InMux
    port map (
            O => \N__14516\,
            I => \N__14512\
        );

    \I__2800\ : InMux
    port map (
            O => \N__14515\,
            I => \N__14509\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__14512\,
            I => \N__14506\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__14509\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__2797\ : Odrv4
    port map (
            O => \N__14506\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__2796\ : InMux
    port map (
            O => \N__14501\,
            I => \N__14498\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__14498\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13\
        );

    \I__2794\ : InMux
    port map (
            O => \N__14495\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11\
        );

    \I__2793\ : InMux
    port map (
            O => \N__14492\,
            I => \N__14488\
        );

    \I__2792\ : InMux
    port map (
            O => \N__14491\,
            I => \N__14485\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__14488\,
            I => \N__14482\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__14485\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__2789\ : Odrv4
    port map (
            O => \N__14482\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__2788\ : CascadeMux
    port map (
            O => \N__14477\,
            I => \N__14474\
        );

    \I__2787\ : InMux
    port map (
            O => \N__14474\,
            I => \N__14471\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__14471\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14\
        );

    \I__2785\ : InMux
    port map (
            O => \N__14468\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12\
        );

    \I__2784\ : InMux
    port map (
            O => \N__14465\,
            I => \N__14461\
        );

    \I__2783\ : InMux
    port map (
            O => \N__14464\,
            I => \N__14458\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__14461\,
            I => \N__14455\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__14458\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__2780\ : Odrv4
    port map (
            O => \N__14455\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__2779\ : InMux
    port map (
            O => \N__14450\,
            I => \N__14447\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__14447\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15\
        );

    \I__2777\ : InMux
    port map (
            O => \N__14444\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13\
        );

    \I__2776\ : InMux
    port map (
            O => \N__14441\,
            I => \N__14437\
        );

    \I__2775\ : InMux
    port map (
            O => \N__14440\,
            I => \N__14434\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__14437\,
            I => \N__14430\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__14434\,
            I => \N__14427\
        );

    \I__2772\ : InMux
    port map (
            O => \N__14433\,
            I => \N__14424\
        );

    \I__2771\ : Odrv4
    port map (
            O => \N__14430\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__2770\ : Odrv12
    port map (
            O => \N__14427\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__14424\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__2768\ : CascadeMux
    port map (
            O => \N__14417\,
            I => \N__14414\
        );

    \I__2767\ : InMux
    port map (
            O => \N__14414\,
            I => \N__14411\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__14411\,
            I => \N__14408\
        );

    \I__2765\ : Span4Mux_h
    port map (
            O => \N__14408\,
            I => \N__14405\
        );

    \I__2764\ : Odrv4
    port map (
            O => \N__14405\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\
        );

    \I__2763\ : InMux
    port map (
            O => \N__14402\,
            I => \N__14399\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__14399\,
            I => \N__14395\
        );

    \I__2761\ : InMux
    port map (
            O => \N__14398\,
            I => \N__14392\
        );

    \I__2760\ : Odrv12
    port map (
            O => \N__14395\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__14392\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__2758\ : InMux
    port map (
            O => \N__14387\,
            I => \N__14384\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__14384\,
            I => \N__14381\
        );

    \I__2756\ : Span4Mux_h
    port map (
            O => \N__14381\,
            I => \N__14378\
        );

    \I__2755\ : Odrv4
    port map (
            O => \N__14378\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2\
        );

    \I__2754\ : InMux
    port map (
            O => \N__14375\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0\
        );

    \I__2753\ : InMux
    port map (
            O => \N__14372\,
            I => \N__14369\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__14369\,
            I => \N__14365\
        );

    \I__2751\ : InMux
    port map (
            O => \N__14368\,
            I => \N__14362\
        );

    \I__2750\ : Odrv12
    port map (
            O => \N__14365\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__14362\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__2748\ : CascadeMux
    port map (
            O => \N__14357\,
            I => \N__14354\
        );

    \I__2747\ : InMux
    port map (
            O => \N__14354\,
            I => \N__14351\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__14351\,
            I => \N__14348\
        );

    \I__2745\ : Span4Mux_h
    port map (
            O => \N__14348\,
            I => \N__14345\
        );

    \I__2744\ : Odrv4
    port map (
            O => \N__14345\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6\
        );

    \I__2743\ : CascadeMux
    port map (
            O => \N__14342\,
            I => \N__14339\
        );

    \I__2742\ : InMux
    port map (
            O => \N__14339\,
            I => \N__14336\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__14336\,
            I => \N__14333\
        );

    \I__2740\ : Odrv12
    port map (
            O => \N__14333\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3\
        );

    \I__2739\ : InMux
    port map (
            O => \N__14330\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1\
        );

    \I__2738\ : CascadeMux
    port map (
            O => \N__14327\,
            I => \N__14324\
        );

    \I__2737\ : InMux
    port map (
            O => \N__14324\,
            I => \N__14321\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__14321\,
            I => \N__14317\
        );

    \I__2735\ : InMux
    port map (
            O => \N__14320\,
            I => \N__14314\
        );

    \I__2734\ : Odrv12
    port map (
            O => \N__14317\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__14314\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__2732\ : InMux
    port map (
            O => \N__14309\,
            I => \N__14306\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__14306\,
            I => \N__14303\
        );

    \I__2730\ : Span4Mux_h
    port map (
            O => \N__14303\,
            I => \N__14300\
        );

    \I__2729\ : Odrv4
    port map (
            O => \N__14300\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4\
        );

    \I__2728\ : InMux
    port map (
            O => \N__14297\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2\
        );

    \I__2727\ : CascadeMux
    port map (
            O => \N__14294\,
            I => \N__14291\
        );

    \I__2726\ : InMux
    port map (
            O => \N__14291\,
            I => \N__14288\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__14288\,
            I => \N__14284\
        );

    \I__2724\ : InMux
    port map (
            O => \N__14287\,
            I => \N__14281\
        );

    \I__2723\ : Odrv12
    port map (
            O => \N__14284\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__14281\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__2721\ : CascadeMux
    port map (
            O => \N__14276\,
            I => \N__14273\
        );

    \I__2720\ : InMux
    port map (
            O => \N__14273\,
            I => \N__14270\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__14270\,
            I => \N__14267\
        );

    \I__2718\ : Span4Mux_h
    port map (
            O => \N__14267\,
            I => \N__14264\
        );

    \I__2717\ : Odrv4
    port map (
            O => \N__14264\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5\
        );

    \I__2716\ : InMux
    port map (
            O => \N__14261\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3\
        );

    \I__2715\ : InMux
    port map (
            O => \N__14258\,
            I => \N__14255\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__14255\,
            I => \N__14251\
        );

    \I__2713\ : InMux
    port map (
            O => \N__14254\,
            I => \N__14248\
        );

    \I__2712\ : Odrv12
    port map (
            O => \N__14251\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__14248\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__2710\ : CascadeMux
    port map (
            O => \N__14243\,
            I => \N__14240\
        );

    \I__2709\ : InMux
    port map (
            O => \N__14240\,
            I => \N__14237\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__14237\,
            I => \N__14234\
        );

    \I__2707\ : Span4Mux_h
    port map (
            O => \N__14234\,
            I => \N__14231\
        );

    \I__2706\ : Odrv4
    port map (
            O => \N__14231\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6\
        );

    \I__2705\ : InMux
    port map (
            O => \N__14228\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4\
        );

    \I__2704\ : InMux
    port map (
            O => \N__14225\,
            I => \N__14221\
        );

    \I__2703\ : InMux
    port map (
            O => \N__14224\,
            I => \N__14218\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__14221\,
            I => \N__14215\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__14218\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__2700\ : Odrv4
    port map (
            O => \N__14215\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__2699\ : InMux
    port map (
            O => \N__14210\,
            I => \N__14207\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__14207\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7\
        );

    \I__2697\ : InMux
    port map (
            O => \N__14204\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5\
        );

    \I__2696\ : InMux
    port map (
            O => \N__14201\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_20\
        );

    \I__2695\ : InMux
    port map (
            O => \N__14198\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_21\
        );

    \I__2694\ : InMux
    port map (
            O => \N__14195\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_22\
        );

    \I__2693\ : InMux
    port map (
            O => \N__14192\,
            I => \bfn_8_16_0_\
        );

    \I__2692\ : InMux
    port map (
            O => \N__14189\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_24\
        );

    \I__2691\ : InMux
    port map (
            O => \N__14186\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_25\
        );

    \I__2690\ : InMux
    port map (
            O => \N__14183\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_26\
        );

    \I__2689\ : InMux
    port map (
            O => \N__14180\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_27\
        );

    \I__2688\ : InMux
    port map (
            O => \N__14177\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_28\
        );

    \I__2687\ : CEMux
    port map (
            O => \N__14174\,
            I => \N__14162\
        );

    \I__2686\ : CEMux
    port map (
            O => \N__14173\,
            I => \N__14162\
        );

    \I__2685\ : CEMux
    port map (
            O => \N__14172\,
            I => \N__14162\
        );

    \I__2684\ : CEMux
    port map (
            O => \N__14171\,
            I => \N__14162\
        );

    \I__2683\ : GlobalMux
    port map (
            O => \N__14162\,
            I => \N__14159\
        );

    \I__2682\ : gio2CtrlBuf
    port map (
            O => \N__14159\,
            I => \delay_measurement_inst.delay_tr_timer.N_256_i_g\
        );

    \I__2681\ : InMux
    port map (
            O => \N__14156\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_10\
        );

    \I__2680\ : InMux
    port map (
            O => \N__14153\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_11\
        );

    \I__2679\ : InMux
    port map (
            O => \N__14150\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_12\
        );

    \I__2678\ : InMux
    port map (
            O => \N__14147\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_13\
        );

    \I__2677\ : InMux
    port map (
            O => \N__14144\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_14\
        );

    \I__2676\ : InMux
    port map (
            O => \N__14141\,
            I => \bfn_8_15_0_\
        );

    \I__2675\ : InMux
    port map (
            O => \N__14138\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_16\
        );

    \I__2674\ : InMux
    port map (
            O => \N__14135\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_17\
        );

    \I__2673\ : InMux
    port map (
            O => \N__14132\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_18\
        );

    \I__2672\ : InMux
    port map (
            O => \N__14129\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_19\
        );

    \I__2671\ : InMux
    port map (
            O => \N__14126\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_1\
        );

    \I__2670\ : InMux
    port map (
            O => \N__14123\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_2\
        );

    \I__2669\ : InMux
    port map (
            O => \N__14120\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_3\
        );

    \I__2668\ : InMux
    port map (
            O => \N__14117\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_4\
        );

    \I__2667\ : InMux
    port map (
            O => \N__14114\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_5\
        );

    \I__2666\ : InMux
    port map (
            O => \N__14111\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_6\
        );

    \I__2665\ : InMux
    port map (
            O => \N__14108\,
            I => \bfn_8_14_0_\
        );

    \I__2664\ : InMux
    port map (
            O => \N__14105\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_8\
        );

    \I__2663\ : InMux
    port map (
            O => \N__14102\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_9\
        );

    \I__2662\ : InMux
    port map (
            O => \N__14099\,
            I => \N__14096\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__14096\,
            I => \N__14092\
        );

    \I__2660\ : InMux
    port map (
            O => \N__14095\,
            I => \N__14089\
        );

    \I__2659\ : Span4Mux_h
    port map (
            O => \N__14092\,
            I => \N__14085\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__14089\,
            I => \N__14082\
        );

    \I__2657\ : InMux
    port map (
            O => \N__14088\,
            I => \N__14079\
        );

    \I__2656\ : Span4Mux_v
    port map (
            O => \N__14085\,
            I => \N__14076\
        );

    \I__2655\ : Span4Mux_v
    port map (
            O => \N__14082\,
            I => \N__14071\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__14079\,
            I => \N__14071\
        );

    \I__2653\ : Odrv4
    port map (
            O => \N__14076\,
            I => measured_delay_hc_6
        );

    \I__2652\ : Odrv4
    port map (
            O => \N__14071\,
            I => measured_delay_hc_6
        );

    \I__2651\ : InMux
    port map (
            O => \N__14066\,
            I => \N__14063\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__14063\,
            I => \N__14058\
        );

    \I__2649\ : InMux
    port map (
            O => \N__14062\,
            I => \N__14055\
        );

    \I__2648\ : InMux
    port map (
            O => \N__14061\,
            I => \N__14051\
        );

    \I__2647\ : Span4Mux_v
    port map (
            O => \N__14058\,
            I => \N__14048\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__14055\,
            I => \N__14045\
        );

    \I__2645\ : InMux
    port map (
            O => \N__14054\,
            I => \N__14042\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__14051\,
            I => \N__14039\
        );

    \I__2643\ : Span4Mux_v
    port map (
            O => \N__14048\,
            I => \N__14032\
        );

    \I__2642\ : Span4Mux_v
    port map (
            O => \N__14045\,
            I => \N__14032\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__14042\,
            I => \N__14032\
        );

    \I__2640\ : Span4Mux_h
    port map (
            O => \N__14039\,
            I => \N__14029\
        );

    \I__2639\ : Odrv4
    port map (
            O => \N__14032\,
            I => measured_delay_hc_17
        );

    \I__2638\ : Odrv4
    port map (
            O => \N__14029\,
            I => measured_delay_hc_17
        );

    \I__2637\ : InMux
    port map (
            O => \N__14024\,
            I => \N__14021\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__14021\,
            I => \N__14016\
        );

    \I__2635\ : InMux
    port map (
            O => \N__14020\,
            I => \N__14012\
        );

    \I__2634\ : InMux
    port map (
            O => \N__14019\,
            I => \N__14009\
        );

    \I__2633\ : Span4Mux_h
    port map (
            O => \N__14016\,
            I => \N__14006\
        );

    \I__2632\ : InMux
    port map (
            O => \N__14015\,
            I => \N__14003\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__14012\,
            I => \N__14000\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__14009\,
            I => \N__13997\
        );

    \I__2629\ : Span4Mux_v
    port map (
            O => \N__14006\,
            I => \N__13994\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__14003\,
            I => \N__13991\
        );

    \I__2627\ : Span4Mux_h
    port map (
            O => \N__14000\,
            I => \N__13986\
        );

    \I__2626\ : Span4Mux_h
    port map (
            O => \N__13997\,
            I => \N__13986\
        );

    \I__2625\ : Odrv4
    port map (
            O => \N__13994\,
            I => measured_delay_hc_16
        );

    \I__2624\ : Odrv4
    port map (
            O => \N__13991\,
            I => measured_delay_hc_16
        );

    \I__2623\ : Odrv4
    port map (
            O => \N__13986\,
            I => measured_delay_hc_16
        );

    \I__2622\ : InMux
    port map (
            O => \N__13979\,
            I => \N__13976\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__13976\,
            I => \N__13970\
        );

    \I__2620\ : InMux
    port map (
            O => \N__13975\,
            I => \N__13967\
        );

    \I__2619\ : InMux
    port map (
            O => \N__13974\,
            I => \N__13961\
        );

    \I__2618\ : InMux
    port map (
            O => \N__13973\,
            I => \N__13961\
        );

    \I__2617\ : Span4Mux_v
    port map (
            O => \N__13970\,
            I => \N__13958\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__13967\,
            I => \N__13955\
        );

    \I__2615\ : InMux
    port map (
            O => \N__13966\,
            I => \N__13952\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__13961\,
            I => \N__13949\
        );

    \I__2613\ : Span4Mux_v
    port map (
            O => \N__13958\,
            I => \N__13942\
        );

    \I__2612\ : Span4Mux_v
    port map (
            O => \N__13955\,
            I => \N__13942\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__13952\,
            I => \N__13942\
        );

    \I__2610\ : Span4Mux_h
    port map (
            O => \N__13949\,
            I => \N__13939\
        );

    \I__2609\ : Odrv4
    port map (
            O => \N__13942\,
            I => measured_delay_hc_14
        );

    \I__2608\ : Odrv4
    port map (
            O => \N__13939\,
            I => measured_delay_hc_14
        );

    \I__2607\ : InMux
    port map (
            O => \N__13934\,
            I => \N__13930\
        );

    \I__2606\ : InMux
    port map (
            O => \N__13933\,
            I => \N__13927\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__13930\,
            I => \N__13923\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__13927\,
            I => \N__13919\
        );

    \I__2603\ : InMux
    port map (
            O => \N__13926\,
            I => \N__13916\
        );

    \I__2602\ : Span4Mux_h
    port map (
            O => \N__13923\,
            I => \N__13913\
        );

    \I__2601\ : InMux
    port map (
            O => \N__13922\,
            I => \N__13910\
        );

    \I__2600\ : Span4Mux_h
    port map (
            O => \N__13919\,
            I => \N__13907\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__13916\,
            I => \N__13904\
        );

    \I__2598\ : Span4Mux_v
    port map (
            O => \N__13913\,
            I => \N__13901\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__13910\,
            I => \N__13898\
        );

    \I__2596\ : Span4Mux_v
    port map (
            O => \N__13907\,
            I => \N__13893\
        );

    \I__2595\ : Span4Mux_h
    port map (
            O => \N__13904\,
            I => \N__13893\
        );

    \I__2594\ : Span4Mux_v
    port map (
            O => \N__13901\,
            I => \N__13888\
        );

    \I__2593\ : Span4Mux_h
    port map (
            O => \N__13898\,
            I => \N__13888\
        );

    \I__2592\ : Odrv4
    port map (
            O => \N__13893\,
            I => measured_delay_hc_18
        );

    \I__2591\ : Odrv4
    port map (
            O => \N__13888\,
            I => measured_delay_hc_18
        );

    \I__2590\ : InMux
    port map (
            O => \N__13883\,
            I => \N__13878\
        );

    \I__2589\ : InMux
    port map (
            O => \N__13882\,
            I => \N__13875\
        );

    \I__2588\ : InMux
    port map (
            O => \N__13881\,
            I => \N__13872\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__13878\,
            I => \N__13868\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__13875\,
            I => \N__13863\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__13872\,
            I => \N__13863\
        );

    \I__2584\ : InMux
    port map (
            O => \N__13871\,
            I => \N__13860\
        );

    \I__2583\ : Span12Mux_v
    port map (
            O => \N__13868\,
            I => \N__13857\
        );

    \I__2582\ : Span4Mux_v
    port map (
            O => \N__13863\,
            I => \N__13854\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__13860\,
            I => measured_delay_hc_7
        );

    \I__2580\ : Odrv12
    port map (
            O => \N__13857\,
            I => measured_delay_hc_7
        );

    \I__2579\ : Odrv4
    port map (
            O => \N__13854\,
            I => measured_delay_hc_7
        );

    \I__2578\ : InMux
    port map (
            O => \N__13847\,
            I => \N__13843\
        );

    \I__2577\ : InMux
    port map (
            O => \N__13846\,
            I => \N__13839\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__13843\,
            I => \N__13835\
        );

    \I__2575\ : InMux
    port map (
            O => \N__13842\,
            I => \N__13832\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__13839\,
            I => \N__13829\
        );

    \I__2573\ : InMux
    port map (
            O => \N__13838\,
            I => \N__13826\
        );

    \I__2572\ : Span12Mux_s7_h
    port map (
            O => \N__13835\,
            I => \N__13823\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__13832\,
            I => \N__13820\
        );

    \I__2570\ : Span4Mux_h
    port map (
            O => \N__13829\,
            I => \N__13817\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__13826\,
            I => measured_delay_hc_8
        );

    \I__2568\ : Odrv12
    port map (
            O => \N__13823\,
            I => measured_delay_hc_8
        );

    \I__2567\ : Odrv4
    port map (
            O => \N__13820\,
            I => measured_delay_hc_8
        );

    \I__2566\ : Odrv4
    port map (
            O => \N__13817\,
            I => measured_delay_hc_8
        );

    \I__2565\ : InMux
    port map (
            O => \N__13808\,
            I => \bfn_8_13_0_\
        );

    \I__2564\ : InMux
    port map (
            O => \N__13805\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_0\
        );

    \I__2563\ : InMux
    port map (
            O => \N__13802\,
            I => \N__13799\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__13799\,
            I => \N__13795\
        );

    \I__2561\ : InMux
    port map (
            O => \N__13798\,
            I => \N__13792\
        );

    \I__2560\ : Span4Mux_v
    port map (
            O => \N__13795\,
            I => \N__13788\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__13792\,
            I => \N__13785\
        );

    \I__2558\ : InMux
    port map (
            O => \N__13791\,
            I => \N__13782\
        );

    \I__2557\ : Span4Mux_v
    port map (
            O => \N__13788\,
            I => \N__13775\
        );

    \I__2556\ : Span4Mux_v
    port map (
            O => \N__13785\,
            I => \N__13775\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__13782\,
            I => \N__13775\
        );

    \I__2554\ : Odrv4
    port map (
            O => \N__13775\,
            I => measured_delay_hc_11
        );

    \I__2553\ : InMux
    port map (
            O => \N__13772\,
            I => \N__13769\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__13769\,
            I => \N__13765\
        );

    \I__2551\ : InMux
    port map (
            O => \N__13768\,
            I => \N__13762\
        );

    \I__2550\ : Span4Mux_v
    port map (
            O => \N__13765\,
            I => \N__13758\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__13762\,
            I => \N__13755\
        );

    \I__2548\ : InMux
    port map (
            O => \N__13761\,
            I => \N__13752\
        );

    \I__2547\ : Span4Mux_v
    port map (
            O => \N__13758\,
            I => \N__13745\
        );

    \I__2546\ : Span4Mux_v
    port map (
            O => \N__13755\,
            I => \N__13745\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__13752\,
            I => \N__13745\
        );

    \I__2544\ : Odrv4
    port map (
            O => \N__13745\,
            I => measured_delay_hc_12
        );

    \I__2543\ : CascadeMux
    port map (
            O => \N__13742\,
            I => \N__13738\
        );

    \I__2542\ : CascadeMux
    port map (
            O => \N__13741\,
            I => \N__13735\
        );

    \I__2541\ : InMux
    port map (
            O => \N__13738\,
            I => \N__13732\
        );

    \I__2540\ : InMux
    port map (
            O => \N__13735\,
            I => \N__13729\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__13732\,
            I => \N__13726\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__13729\,
            I => \N__13722\
        );

    \I__2537\ : Span4Mux_v
    port map (
            O => \N__13726\,
            I => \N__13719\
        );

    \I__2536\ : InMux
    port map (
            O => \N__13725\,
            I => \N__13716\
        );

    \I__2535\ : Span4Mux_h
    port map (
            O => \N__13722\,
            I => \N__13713\
        );

    \I__2534\ : Span4Mux_v
    port map (
            O => \N__13719\,
            I => \N__13708\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__13716\,
            I => \N__13708\
        );

    \I__2532\ : Odrv4
    port map (
            O => \N__13713\,
            I => measured_delay_hc_3
        );

    \I__2531\ : Odrv4
    port map (
            O => \N__13708\,
            I => measured_delay_hc_3
        );

    \I__2530\ : InMux
    port map (
            O => \N__13703\,
            I => \N__13700\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__13700\,
            I => \N__13696\
        );

    \I__2528\ : InMux
    port map (
            O => \N__13699\,
            I => \N__13693\
        );

    \I__2527\ : Span4Mux_v
    port map (
            O => \N__13696\,
            I => \N__13689\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__13693\,
            I => \N__13686\
        );

    \I__2525\ : InMux
    port map (
            O => \N__13692\,
            I => \N__13683\
        );

    \I__2524\ : Span4Mux_v
    port map (
            O => \N__13689\,
            I => \N__13676\
        );

    \I__2523\ : Span4Mux_v
    port map (
            O => \N__13686\,
            I => \N__13676\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__13683\,
            I => \N__13676\
        );

    \I__2521\ : Odrv4
    port map (
            O => \N__13676\,
            I => measured_delay_hc_4
        );

    \I__2520\ : CascadeMux
    port map (
            O => \N__13673\,
            I => \N__13666\
        );

    \I__2519\ : InMux
    port map (
            O => \N__13672\,
            I => \N__13655\
        );

    \I__2518\ : InMux
    port map (
            O => \N__13671\,
            I => \N__13655\
        );

    \I__2517\ : InMux
    port map (
            O => \N__13670\,
            I => \N__13655\
        );

    \I__2516\ : InMux
    port map (
            O => \N__13669\,
            I => \N__13655\
        );

    \I__2515\ : InMux
    port map (
            O => \N__13666\,
            I => \N__13655\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__13655\,
            I => \delay_measurement_inst.delay_hc_reg_3_0_a2_0_6\
        );

    \I__2513\ : CascadeMux
    port map (
            O => \N__13652\,
            I => \N__13649\
        );

    \I__2512\ : InMux
    port map (
            O => \N__13649\,
            I => \N__13645\
        );

    \I__2511\ : CascadeMux
    port map (
            O => \N__13648\,
            I => \N__13642\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__13645\,
            I => \N__13639\
        );

    \I__2509\ : InMux
    port map (
            O => \N__13642\,
            I => \N__13636\
        );

    \I__2508\ : Span4Mux_h
    port map (
            O => \N__13639\,
            I => \N__13633\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__13636\,
            I => \N__13630\
        );

    \I__2506\ : Span4Mux_v
    port map (
            O => \N__13633\,
            I => \N__13627\
        );

    \I__2505\ : Span4Mux_h
    port map (
            O => \N__13630\,
            I => \N__13624\
        );

    \I__2504\ : Odrv4
    port map (
            O => \N__13627\,
            I => measured_delay_hc_1
        );

    \I__2503\ : Odrv4
    port map (
            O => \N__13624\,
            I => measured_delay_hc_1
        );

    \I__2502\ : InMux
    port map (
            O => \N__13619\,
            I => \N__13615\
        );

    \I__2501\ : InMux
    port map (
            O => \N__13618\,
            I => \N__13612\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__13615\,
            I => \N__13608\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__13612\,
            I => \N__13605\
        );

    \I__2498\ : InMux
    port map (
            O => \N__13611\,
            I => \N__13602\
        );

    \I__2497\ : Span12Mux_v
    port map (
            O => \N__13608\,
            I => \N__13599\
        );

    \I__2496\ : Span4Mux_v
    port map (
            O => \N__13605\,
            I => \N__13594\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__13602\,
            I => \N__13594\
        );

    \I__2494\ : Odrv12
    port map (
            O => \N__13599\,
            I => measured_delay_hc_10
        );

    \I__2493\ : Odrv4
    port map (
            O => \N__13594\,
            I => measured_delay_hc_10
        );

    \I__2492\ : InMux
    port map (
            O => \N__13589\,
            I => \N__13586\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__13586\,
            I => \N__13581\
        );

    \I__2490\ : InMux
    port map (
            O => \N__13585\,
            I => \N__13578\
        );

    \I__2489\ : InMux
    port map (
            O => \N__13584\,
            I => \N__13575\
        );

    \I__2488\ : Span4Mux_v
    port map (
            O => \N__13581\,
            I => \N__13572\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__13578\,
            I => \N__13569\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__13575\,
            I => \N__13566\
        );

    \I__2485\ : Span4Mux_v
    port map (
            O => \N__13572\,
            I => \N__13559\
        );

    \I__2484\ : Span4Mux_v
    port map (
            O => \N__13569\,
            I => \N__13559\
        );

    \I__2483\ : Span4Mux_v
    port map (
            O => \N__13566\,
            I => \N__13559\
        );

    \I__2482\ : Odrv4
    port map (
            O => \N__13559\,
            I => measured_delay_hc_9
        );

    \I__2481\ : InMux
    port map (
            O => \N__13556\,
            I => \N__13543\
        );

    \I__2480\ : InMux
    port map (
            O => \N__13555\,
            I => \N__13543\
        );

    \I__2479\ : InMux
    port map (
            O => \N__13554\,
            I => \N__13543\
        );

    \I__2478\ : CascadeMux
    port map (
            O => \N__13553\,
            I => \N__13537\
        );

    \I__2477\ : InMux
    port map (
            O => \N__13552\,
            I => \N__13530\
        );

    \I__2476\ : InMux
    port map (
            O => \N__13551\,
            I => \N__13530\
        );

    \I__2475\ : InMux
    port map (
            O => \N__13550\,
            I => \N__13530\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__13543\,
            I => \N__13527\
        );

    \I__2473\ : InMux
    port map (
            O => \N__13542\,
            I => \N__13522\
        );

    \I__2472\ : InMux
    port map (
            O => \N__13541\,
            I => \N__13522\
        );

    \I__2471\ : InMux
    port map (
            O => \N__13540\,
            I => \N__13517\
        );

    \I__2470\ : InMux
    port map (
            O => \N__13537\,
            I => \N__13517\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__13530\,
            I => \N__13514\
        );

    \I__2468\ : Span4Mux_v
    port map (
            O => \N__13527\,
            I => \N__13507\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__13522\,
            I => \N__13507\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__13517\,
            I => \N__13507\
        );

    \I__2465\ : Span4Mux_v
    port map (
            O => \N__13514\,
            I => \N__13502\
        );

    \I__2464\ : Span4Mux_v
    port map (
            O => \N__13507\,
            I => \N__13502\
        );

    \I__2463\ : Odrv4
    port map (
            O => \N__13502\,
            I => measured_delay_hc_15
        );

    \I__2462\ : CascadeMux
    port map (
            O => \N__13499\,
            I => \N__13495\
        );

    \I__2461\ : InMux
    port map (
            O => \N__13498\,
            I => \N__13492\
        );

    \I__2460\ : InMux
    port map (
            O => \N__13495\,
            I => \N__13487\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__13492\,
            I => \N__13484\
        );

    \I__2458\ : InMux
    port map (
            O => \N__13491\,
            I => \N__13481\
        );

    \I__2457\ : CascadeMux
    port map (
            O => \N__13490\,
            I => \N__13478\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__13487\,
            I => \N__13475\
        );

    \I__2455\ : Span4Mux_v
    port map (
            O => \N__13484\,
            I => \N__13472\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__13481\,
            I => \N__13469\
        );

    \I__2453\ : InMux
    port map (
            O => \N__13478\,
            I => \N__13466\
        );

    \I__2452\ : Span4Mux_h
    port map (
            O => \N__13475\,
            I => \N__13463\
        );

    \I__2451\ : Span4Mux_v
    port map (
            O => \N__13472\,
            I => \N__13458\
        );

    \I__2450\ : Span4Mux_v
    port map (
            O => \N__13469\,
            I => \N__13458\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__13466\,
            I => \N__13455\
        );

    \I__2448\ : Span4Mux_h
    port map (
            O => \N__13463\,
            I => \N__13452\
        );

    \I__2447\ : Odrv4
    port map (
            O => \N__13458\,
            I => measured_delay_hc_19
        );

    \I__2446\ : Odrv12
    port map (
            O => \N__13455\,
            I => measured_delay_hc_19
        );

    \I__2445\ : Odrv4
    port map (
            O => \N__13452\,
            I => measured_delay_hc_19
        );

    \I__2444\ : CascadeMux
    port map (
            O => \N__13445\,
            I => \N__13442\
        );

    \I__2443\ : InMux
    port map (
            O => \N__13442\,
            I => \N__13439\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__13439\,
            I => \N__13436\
        );

    \I__2441\ : Span4Mux_h
    port map (
            O => \N__13436\,
            I => \N__13433\
        );

    \I__2440\ : Odrv4
    port map (
            O => \N__13433\,
            I => \phase_controller_slave.stoper_tr.time_passed_1_sqmuxa\
        );

    \I__2439\ : InMux
    port map (
            O => \N__13430\,
            I => \N__13427\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__13427\,
            I => \N__13424\
        );

    \I__2437\ : Odrv12
    port map (
            O => \N__13424\,
            I => \il_min_comp2_D1\
        );

    \I__2436\ : CascadeMux
    port map (
            O => \N__13421\,
            I => \N__13418\
        );

    \I__2435\ : InMux
    port map (
            O => \N__13418\,
            I => \N__13413\
        );

    \I__2434\ : InMux
    port map (
            O => \N__13417\,
            I => \N__13410\
        );

    \I__2433\ : InMux
    port map (
            O => \N__13416\,
            I => \N__13407\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__13413\,
            I => \N__13404\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__13410\,
            I => \N__13401\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__13407\,
            I => \N__13398\
        );

    \I__2429\ : Span4Mux_v
    port map (
            O => \N__13404\,
            I => \N__13395\
        );

    \I__2428\ : Span4Mux_h
    port map (
            O => \N__13401\,
            I => \N__13392\
        );

    \I__2427\ : Span4Mux_h
    port map (
            O => \N__13398\,
            I => \N__13389\
        );

    \I__2426\ : Odrv4
    port map (
            O => \N__13395\,
            I => \il_min_comp2_D2\
        );

    \I__2425\ : Odrv4
    port map (
            O => \N__13392\,
            I => \il_min_comp2_D2\
        );

    \I__2424\ : Odrv4
    port map (
            O => \N__13389\,
            I => \il_min_comp2_D2\
        );

    \I__2423\ : InMux
    port map (
            O => \N__13382\,
            I => \N__13379\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__13379\,
            I => \N__13374\
        );

    \I__2421\ : InMux
    port map (
            O => \N__13378\,
            I => \N__13371\
        );

    \I__2420\ : InMux
    port map (
            O => \N__13377\,
            I => \N__13368\
        );

    \I__2419\ : Span4Mux_h
    port map (
            O => \N__13374\,
            I => \N__13365\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__13371\,
            I => \N__13362\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__13368\,
            I => \N__13359\
        );

    \I__2416\ : Span4Mux_v
    port map (
            O => \N__13365\,
            I => \N__13356\
        );

    \I__2415\ : Span4Mux_h
    port map (
            O => \N__13362\,
            I => \N__13353\
        );

    \I__2414\ : Span4Mux_h
    port map (
            O => \N__13359\,
            I => \N__13350\
        );

    \I__2413\ : Odrv4
    port map (
            O => \N__13356\,
            I => measured_delay_hc_5
        );

    \I__2412\ : Odrv4
    port map (
            O => \N__13353\,
            I => measured_delay_hc_5
        );

    \I__2411\ : Odrv4
    port map (
            O => \N__13350\,
            I => measured_delay_hc_5
        );

    \I__2410\ : InMux
    port map (
            O => \N__13343\,
            I => \N__13340\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__13340\,
            I => \N__13336\
        );

    \I__2408\ : InMux
    port map (
            O => \N__13339\,
            I => \N__13333\
        );

    \I__2407\ : Span4Mux_h
    port map (
            O => \N__13336\,
            I => \N__13329\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__13333\,
            I => \N__13326\
        );

    \I__2405\ : InMux
    port map (
            O => \N__13332\,
            I => \N__13323\
        );

    \I__2404\ : Span4Mux_v
    port map (
            O => \N__13329\,
            I => \N__13320\
        );

    \I__2403\ : Span4Mux_h
    port map (
            O => \N__13326\,
            I => \N__13317\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__13323\,
            I => \N__13314\
        );

    \I__2401\ : Odrv4
    port map (
            O => \N__13320\,
            I => measured_delay_hc_2
        );

    \I__2400\ : Odrv4
    port map (
            O => \N__13317\,
            I => measured_delay_hc_2
        );

    \I__2399\ : Odrv12
    port map (
            O => \N__13314\,
            I => measured_delay_hc_2
        );

    \I__2398\ : CascadeMux
    port map (
            O => \N__13307\,
            I => \N__13303\
        );

    \I__2397\ : InMux
    port map (
            O => \N__13306\,
            I => \N__13297\
        );

    \I__2396\ : InMux
    port map (
            O => \N__13303\,
            I => \N__13297\
        );

    \I__2395\ : InMux
    port map (
            O => \N__13302\,
            I => \N__13294\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__13297\,
            I => \phase_controller_slave.stateZ0Z_2\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__13294\,
            I => \phase_controller_slave.stateZ0Z_2\
        );

    \I__2392\ : InMux
    port map (
            O => \N__13289\,
            I => \N__13283\
        );

    \I__2391\ : InMux
    port map (
            O => \N__13288\,
            I => \N__13283\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__13283\,
            I => \N__13278\
        );

    \I__2389\ : InMux
    port map (
            O => \N__13282\,
            I => \N__13275\
        );

    \I__2388\ : InMux
    port map (
            O => \N__13281\,
            I => \N__13272\
        );

    \I__2387\ : Span4Mux_h
    port map (
            O => \N__13278\,
            I => \N__13267\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__13275\,
            I => \N__13267\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__13272\,
            I => \phase_controller_slave.hc_time_passed\
        );

    \I__2384\ : Odrv4
    port map (
            O => \N__13267\,
            I => \phase_controller_slave.hc_time_passed\
        );

    \I__2383\ : CascadeMux
    port map (
            O => \N__13262\,
            I => \N__13259\
        );

    \I__2382\ : InMux
    port map (
            O => \N__13259\,
            I => \N__13256\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__13256\,
            I => \N__13253\
        );

    \I__2380\ : Odrv4
    port map (
            O => \N__13253\,
            I => \phase_controller_slave.start_timer_hc_RNOZ0Z_0\
        );

    \I__2379\ : InMux
    port map (
            O => \N__13250\,
            I => \N__13247\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__13247\,
            I => \N__13244\
        );

    \I__2377\ : Span4Mux_v
    port map (
            O => \N__13244\,
            I => \N__13241\
        );

    \I__2376\ : Span4Mux_v
    port map (
            O => \N__13241\,
            I => \N__13238\
        );

    \I__2375\ : Odrv4
    port map (
            O => \N__13238\,
            I => il_max_comp1_c
        );

    \I__2374\ : InMux
    port map (
            O => \N__13235\,
            I => \N__13232\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__13232\,
            I => \N__13229\
        );

    \I__2372\ : Span12Mux_v
    port map (
            O => \N__13229\,
            I => \N__13226\
        );

    \I__2371\ : Odrv12
    port map (
            O => \N__13226\,
            I => il_min_comp2_c
        );

    \I__2370\ : InMux
    port map (
            O => \N__13223\,
            I => \N__13220\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__13220\,
            I => \il_max_comp1_D1\
        );

    \I__2368\ : InMux
    port map (
            O => \N__13217\,
            I => \N__13213\
        );

    \I__2367\ : InMux
    port map (
            O => \N__13216\,
            I => \N__13210\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__13213\,
            I => \N__13205\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__13210\,
            I => \N__13205\
        );

    \I__2364\ : Span4Mux_h
    port map (
            O => \N__13205\,
            I => \N__13201\
        );

    \I__2363\ : InMux
    port map (
            O => \N__13204\,
            I => \N__13198\
        );

    \I__2362\ : Odrv4
    port map (
            O => \N__13201\,
            I => \il_max_comp1_D2\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__13198\,
            I => \il_max_comp1_D2\
        );

    \I__2360\ : InMux
    port map (
            O => \N__13193\,
            I => \N__13190\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__13190\,
            I => \N__13187\
        );

    \I__2358\ : Odrv12
    port map (
            O => \N__13187\,
            I => \phase_controller_inst1.start_timer_hc_0_sqmuxa\
        );

    \I__2357\ : InMux
    port map (
            O => \N__13184\,
            I => \N__13181\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__13181\,
            I => \N__13178\
        );

    \I__2355\ : Span4Mux_v
    port map (
            O => \N__13178\,
            I => \N__13175\
        );

    \I__2354\ : Sp12to4
    port map (
            O => \N__13175\,
            I => \N__13172\
        );

    \I__2353\ : Span12Mux_h
    port map (
            O => \N__13172\,
            I => \N__13169\
        );

    \I__2352\ : Odrv12
    port map (
            O => \N__13169\,
            I => il_min_comp1_c
        );

    \I__2351\ : InMux
    port map (
            O => \N__13166\,
            I => \N__13163\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__13163\,
            I => \il_min_comp1_D1\
        );

    \I__2349\ : InMux
    port map (
            O => \N__13160\,
            I => \N__13154\
        );

    \I__2348\ : InMux
    port map (
            O => \N__13159\,
            I => \N__13154\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__13154\,
            I => \N__13151\
        );

    \I__2346\ : Span4Mux_h
    port map (
            O => \N__13151\,
            I => \N__13147\
        );

    \I__2345\ : InMux
    port map (
            O => \N__13150\,
            I => \N__13144\
        );

    \I__2344\ : Odrv4
    port map (
            O => \N__13147\,
            I => \il_min_comp1_D2\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__13144\,
            I => \il_min_comp1_D2\
        );

    \I__2342\ : InMux
    port map (
            O => \N__13139\,
            I => \N__13133\
        );

    \I__2341\ : InMux
    port map (
            O => \N__13138\,
            I => \N__13133\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__13133\,
            I => \N__13130\
        );

    \I__2339\ : Odrv4
    port map (
            O => \N__13130\,
            I => \phase_controller_inst1.T01_0_sqmuxa\
        );

    \I__2338\ : InMux
    port map (
            O => \N__13127\,
            I => \N__13122\
        );

    \I__2337\ : InMux
    port map (
            O => \N__13126\,
            I => \N__13119\
        );

    \I__2336\ : InMux
    port map (
            O => \N__13125\,
            I => \N__13116\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__13122\,
            I => \N__13113\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__13119\,
            I => \phase_controller_slave.tr_time_passed\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__13116\,
            I => \phase_controller_slave.tr_time_passed\
        );

    \I__2332\ : Odrv4
    port map (
            O => \N__13113\,
            I => \phase_controller_slave.tr_time_passed\
        );

    \I__2331\ : InMux
    port map (
            O => \N__13106\,
            I => \N__13102\
        );

    \I__2330\ : InMux
    port map (
            O => \N__13105\,
            I => \N__13099\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__13102\,
            I => \phase_controller_slave.stateZ0Z_0\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__13099\,
            I => \phase_controller_slave.stateZ0Z_0\
        );

    \I__2327\ : InMux
    port map (
            O => \N__13094\,
            I => \N__13088\
        );

    \I__2326\ : InMux
    port map (
            O => \N__13093\,
            I => \N__13088\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__13088\,
            I => \phase_controller_slave.state_RNIVDE2Z0Z_0\
        );

    \I__2324\ : InMux
    port map (
            O => \N__13085\,
            I => \N__13078\
        );

    \I__2323\ : InMux
    port map (
            O => \N__13084\,
            I => \N__13078\
        );

    \I__2322\ : CascadeMux
    port map (
            O => \N__13083\,
            I => \N__13075\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__13078\,
            I => \N__13072\
        );

    \I__2320\ : InMux
    port map (
            O => \N__13075\,
            I => \N__13068\
        );

    \I__2319\ : Span4Mux_s3_v
    port map (
            O => \N__13072\,
            I => \N__13065\
        );

    \I__2318\ : InMux
    port map (
            O => \N__13071\,
            I => \N__13062\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__13068\,
            I => \N__13059\
        );

    \I__2316\ : Span4Mux_h
    port map (
            O => \N__13065\,
            I => \N__13052\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__13062\,
            I => \N__13052\
        );

    \I__2314\ : Span4Mux_v
    port map (
            O => \N__13059\,
            I => \N__13049\
        );

    \I__2313\ : InMux
    port map (
            O => \N__13058\,
            I => \N__13046\
        );

    \I__2312\ : InMux
    port map (
            O => \N__13057\,
            I => \N__13043\
        );

    \I__2311\ : Sp12to4
    port map (
            O => \N__13052\,
            I => \N__13040\
        );

    \I__2310\ : Span4Mux_v
    port map (
            O => \N__13049\,
            I => \N__13035\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__13046\,
            I => \N__13035\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__13043\,
            I => \N__13032\
        );

    \I__2307\ : Span12Mux_v
    port map (
            O => \N__13040\,
            I => \N__13025\
        );

    \I__2306\ : Sp12to4
    port map (
            O => \N__13035\,
            I => \N__13025\
        );

    \I__2305\ : Sp12to4
    port map (
            O => \N__13032\,
            I => \N__13025\
        );

    \I__2304\ : Span12Mux_v
    port map (
            O => \N__13025\,
            I => \N__13022\
        );

    \I__2303\ : Span12Mux_h
    port map (
            O => \N__13022\,
            I => \N__13019\
        );

    \I__2302\ : Odrv12
    port map (
            O => \N__13019\,
            I => start_stop_c
        );

    \I__2301\ : CascadeMux
    port map (
            O => \N__13016\,
            I => \N__13011\
        );

    \I__2300\ : InMux
    port map (
            O => \N__13015\,
            I => \N__13008\
        );

    \I__2299\ : InMux
    port map (
            O => \N__13014\,
            I => \N__13005\
        );

    \I__2298\ : InMux
    port map (
            O => \N__13011\,
            I => \N__13002\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__13008\,
            I => \N__12997\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__13005\,
            I => \N__12997\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__13002\,
            I => shift_flag_start
        );

    \I__2294\ : Odrv12
    port map (
            O => \N__12997\,
            I => shift_flag_start
        );

    \I__2293\ : InMux
    port map (
            O => \N__12992\,
            I => \N__12989\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__12989\,
            I => \N__12986\
        );

    \I__2291\ : Span12Mux_v
    port map (
            O => \N__12986\,
            I => \N__12983\
        );

    \I__2290\ : Span12Mux_v
    port map (
            O => \N__12983\,
            I => \N__12980\
        );

    \I__2289\ : Odrv12
    port map (
            O => \N__12980\,
            I => il_max_comp2_c
        );

    \I__2288\ : InMux
    port map (
            O => \N__12977\,
            I => \N__12974\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__12974\,
            I => \il_max_comp2_D1\
        );

    \I__2286\ : InMux
    port map (
            O => \N__12971\,
            I => \N__12968\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__12968\,
            I => \N__12965\
        );

    \I__2284\ : Odrv4
    port map (
            O => \N__12965\,
            I => \phase_controller_slave.state_RNO_0Z0Z_3\
        );

    \I__2283\ : InMux
    port map (
            O => \N__12962\,
            I => \N__12955\
        );

    \I__2282\ : InMux
    port map (
            O => \N__12961\,
            I => \N__12955\
        );

    \I__2281\ : InMux
    port map (
            O => \N__12960\,
            I => \N__12952\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__12955\,
            I => \il_max_comp2_D2\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__12952\,
            I => \il_max_comp2_D2\
        );

    \I__2278\ : InMux
    port map (
            O => \N__12947\,
            I => \N__12944\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__12944\,
            I => \phase_controller_slave.start_timer_hc_0_sqmuxa\
        );

    \I__2276\ : CascadeMux
    port map (
            O => \N__12941\,
            I => \N__12937\
        );

    \I__2275\ : InMux
    port map (
            O => \N__12940\,
            I => \N__12931\
        );

    \I__2274\ : InMux
    port map (
            O => \N__12937\,
            I => \N__12931\
        );

    \I__2273\ : CascadeMux
    port map (
            O => \N__12936\,
            I => \N__12928\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__12931\,
            I => \N__12924\
        );

    \I__2271\ : InMux
    port map (
            O => \N__12928\,
            I => \N__12919\
        );

    \I__2270\ : InMux
    port map (
            O => \N__12927\,
            I => \N__12919\
        );

    \I__2269\ : Odrv4
    port map (
            O => \N__12924\,
            I => \phase_controller_slave.stateZ0Z_4\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__12919\,
            I => \phase_controller_slave.stateZ0Z_4\
        );

    \I__2267\ : CascadeMux
    port map (
            O => \N__12914\,
            I => \N__12899\
        );

    \I__2266\ : CascadeMux
    port map (
            O => \N__12913\,
            I => \N__12896\
        );

    \I__2265\ : CascadeMux
    port map (
            O => \N__12912\,
            I => \N__12893\
        );

    \I__2264\ : CascadeMux
    port map (
            O => \N__12911\,
            I => \N__12889\
        );

    \I__2263\ : CascadeMux
    port map (
            O => \N__12910\,
            I => \N__12885\
        );

    \I__2262\ : CascadeMux
    port map (
            O => \N__12909\,
            I => \N__12882\
        );

    \I__2261\ : CascadeMux
    port map (
            O => \N__12908\,
            I => \N__12875\
        );

    \I__2260\ : CascadeMux
    port map (
            O => \N__12907\,
            I => \N__12872\
        );

    \I__2259\ : CascadeMux
    port map (
            O => \N__12906\,
            I => \N__12869\
        );

    \I__2258\ : CascadeMux
    port map (
            O => \N__12905\,
            I => \N__12866\
        );

    \I__2257\ : CascadeMux
    port map (
            O => \N__12904\,
            I => \N__12863\
        );

    \I__2256\ : CascadeMux
    port map (
            O => \N__12903\,
            I => \N__12858\
        );

    \I__2255\ : CascadeMux
    port map (
            O => \N__12902\,
            I => \N__12855\
        );

    \I__2254\ : InMux
    port map (
            O => \N__12899\,
            I => \N__12844\
        );

    \I__2253\ : InMux
    port map (
            O => \N__12896\,
            I => \N__12844\
        );

    \I__2252\ : InMux
    port map (
            O => \N__12893\,
            I => \N__12844\
        );

    \I__2251\ : InMux
    port map (
            O => \N__12892\,
            I => \N__12844\
        );

    \I__2250\ : InMux
    port map (
            O => \N__12889\,
            I => \N__12835\
        );

    \I__2249\ : InMux
    port map (
            O => \N__12888\,
            I => \N__12835\
        );

    \I__2248\ : InMux
    port map (
            O => \N__12885\,
            I => \N__12835\
        );

    \I__2247\ : InMux
    port map (
            O => \N__12882\,
            I => \N__12835\
        );

    \I__2246\ : InMux
    port map (
            O => \N__12881\,
            I => \N__12818\
        );

    \I__2245\ : InMux
    port map (
            O => \N__12880\,
            I => \N__12818\
        );

    \I__2244\ : InMux
    port map (
            O => \N__12879\,
            I => \N__12818\
        );

    \I__2243\ : InMux
    port map (
            O => \N__12878\,
            I => \N__12818\
        );

    \I__2242\ : InMux
    port map (
            O => \N__12875\,
            I => \N__12818\
        );

    \I__2241\ : InMux
    port map (
            O => \N__12872\,
            I => \N__12818\
        );

    \I__2240\ : InMux
    port map (
            O => \N__12869\,
            I => \N__12818\
        );

    \I__2239\ : InMux
    port map (
            O => \N__12866\,
            I => \N__12818\
        );

    \I__2238\ : InMux
    port map (
            O => \N__12863\,
            I => \N__12813\
        );

    \I__2237\ : InMux
    port map (
            O => \N__12862\,
            I => \N__12813\
        );

    \I__2236\ : InMux
    port map (
            O => \N__12861\,
            I => \N__12810\
        );

    \I__2235\ : InMux
    port map (
            O => \N__12858\,
            I => \N__12803\
        );

    \I__2234\ : InMux
    port map (
            O => \N__12855\,
            I => \N__12803\
        );

    \I__2233\ : InMux
    port map (
            O => \N__12854\,
            I => \N__12803\
        );

    \I__2232\ : InMux
    port map (
            O => \N__12853\,
            I => \N__12800\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__12844\,
            I => \N__12794\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__12835\,
            I => \N__12794\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__12818\,
            I => \N__12791\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__12813\,
            I => \N__12786\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__12810\,
            I => \N__12786\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__12803\,
            I => \N__12783\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__12800\,
            I => \N__12780\
        );

    \I__2224\ : InMux
    port map (
            O => \N__12799\,
            I => \N__12777\
        );

    \I__2223\ : Span4Mux_h
    port map (
            O => \N__12794\,
            I => \N__12774\
        );

    \I__2222\ : Span4Mux_h
    port map (
            O => \N__12791\,
            I => \N__12769\
        );

    \I__2221\ : Span4Mux_h
    port map (
            O => \N__12786\,
            I => \N__12769\
        );

    \I__2220\ : Span4Mux_h
    port map (
            O => \N__12783\,
            I => \N__12764\
        );

    \I__2219\ : Span4Mux_h
    port map (
            O => \N__12780\,
            I => \N__12764\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__12777\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__2217\ : Odrv4
    port map (
            O => \N__12774\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__2216\ : Odrv4
    port map (
            O => \N__12769\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__2215\ : Odrv4
    port map (
            O => \N__12764\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__2214\ : InMux
    port map (
            O => \N__12755\,
            I => \N__12752\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__12752\,
            I => \N__12749\
        );

    \I__2212\ : Odrv4
    port map (
            O => \N__12749\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_14\
        );

    \I__2211\ : InMux
    port map (
            O => \N__12746\,
            I => \N__12743\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__12743\,
            I => \N__12740\
        );

    \I__2209\ : Odrv4
    port map (
            O => \N__12740\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_15\
        );

    \I__2208\ : InMux
    port map (
            O => \N__12737\,
            I => \N__12728\
        );

    \I__2207\ : InMux
    port map (
            O => \N__12736\,
            I => \N__12728\
        );

    \I__2206\ : InMux
    port map (
            O => \N__12735\,
            I => \N__12728\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__12728\,
            I => \N__12718\
        );

    \I__2204\ : InMux
    port map (
            O => \N__12727\,
            I => \N__12707\
        );

    \I__2203\ : InMux
    port map (
            O => \N__12726\,
            I => \N__12707\
        );

    \I__2202\ : InMux
    port map (
            O => \N__12725\,
            I => \N__12707\
        );

    \I__2201\ : InMux
    port map (
            O => \N__12724\,
            I => \N__12707\
        );

    \I__2200\ : InMux
    port map (
            O => \N__12723\,
            I => \N__12707\
        );

    \I__2199\ : InMux
    port map (
            O => \N__12722\,
            I => \N__12702\
        );

    \I__2198\ : InMux
    port map (
            O => \N__12721\,
            I => \N__12702\
        );

    \I__2197\ : Odrv4
    port map (
            O => \N__12718\,
            I => \phase_controller_inst1.stoper_tr.N_38\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__12707\,
            I => \phase_controller_inst1.stoper_tr.N_38\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__12702\,
            I => \phase_controller_inst1.stoper_tr.N_38\
        );

    \I__2194\ : InMux
    port map (
            O => \N__12695\,
            I => \N__12692\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__12692\,
            I => \N__12689\
        );

    \I__2192\ : Odrv4
    port map (
            O => \N__12689\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_13\
        );

    \I__2191\ : InMux
    port map (
            O => \N__12686\,
            I => \N__12683\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__12683\,
            I => \N__12680\
        );

    \I__2189\ : Odrv4
    port map (
            O => \N__12680\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_18\
        );

    \I__2188\ : InMux
    port map (
            O => \N__12677\,
            I => \N__12674\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__12674\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_17\
        );

    \I__2186\ : CEMux
    port map (
            O => \N__12671\,
            I => \N__12668\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__12668\,
            I => \N__12663\
        );

    \I__2184\ : CEMux
    port map (
            O => \N__12667\,
            I => \N__12660\
        );

    \I__2183\ : CEMux
    port map (
            O => \N__12666\,
            I => \N__12657\
        );

    \I__2182\ : Span4Mux_v
    port map (
            O => \N__12663\,
            I => \N__12652\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__12660\,
            I => \N__12652\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__12657\,
            I => \N__12649\
        );

    \I__2179\ : Span4Mux_v
    port map (
            O => \N__12652\,
            I => \N__12646\
        );

    \I__2178\ : Span4Mux_h
    port map (
            O => \N__12649\,
            I => \N__12641\
        );

    \I__2177\ : Span4Mux_v
    port map (
            O => \N__12646\,
            I => \N__12641\
        );

    \I__2176\ : Odrv4
    port map (
            O => \N__12641\,
            I => \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__2175\ : InMux
    port map (
            O => \N__12638\,
            I => \N__12635\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__12635\,
            I => \phase_controller_slave.start_timer_tr_0_sqmuxa\
        );

    \I__2173\ : CascadeMux
    port map (
            O => \N__12632\,
            I => \N__12629\
        );

    \I__2172\ : InMux
    port map (
            O => \N__12629\,
            I => \N__12626\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__12626\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_19\
        );

    \I__2170\ : InMux
    port map (
            O => \N__12623\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__2169\ : CascadeMux
    port map (
            O => \N__12620\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO_cascade_\
        );

    \I__2168\ : InMux
    port map (
            O => \N__12617\,
            I => \N__12614\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__12614\,
            I => \N__12611\
        );

    \I__2166\ : Odrv4
    port map (
            O => \N__12611\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0\
        );

    \I__2165\ : InMux
    port map (
            O => \N__12608\,
            I => \N__12605\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__12605\,
            I => \N__12602\
        );

    \I__2163\ : Odrv4
    port map (
            O => \N__12602\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_16\
        );

    \I__2162\ : InMux
    port map (
            O => \N__12599\,
            I => \N__12596\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__12596\,
            I => \N__12593\
        );

    \I__2160\ : Odrv4
    port map (
            O => \N__12593\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_10\
        );

    \I__2159\ : InMux
    port map (
            O => \N__12590\,
            I => \N__12587\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__12587\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_19\
        );

    \I__2157\ : InMux
    port map (
            O => \N__12584\,
            I => \N__12581\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__12581\,
            I => \N__12578\
        );

    \I__2155\ : Odrv4
    port map (
            O => \N__12578\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_11\
        );

    \I__2154\ : CascadeMux
    port map (
            O => \N__12575\,
            I => \N__12572\
        );

    \I__2153\ : InMux
    port map (
            O => \N__12572\,
            I => \N__12569\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__12569\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_11\
        );

    \I__2151\ : InMux
    port map (
            O => \N__12566\,
            I => \N__12563\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__12563\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_12\
        );

    \I__2149\ : CascadeMux
    port map (
            O => \N__12560\,
            I => \N__12557\
        );

    \I__2148\ : InMux
    port map (
            O => \N__12557\,
            I => \N__12554\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__12554\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_12\
        );

    \I__2146\ : CascadeMux
    port map (
            O => \N__12551\,
            I => \N__12548\
        );

    \I__2145\ : InMux
    port map (
            O => \N__12548\,
            I => \N__12545\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__12545\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_13\
        );

    \I__2143\ : CascadeMux
    port map (
            O => \N__12542\,
            I => \N__12539\
        );

    \I__2142\ : InMux
    port map (
            O => \N__12539\,
            I => \N__12536\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__12536\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_14\
        );

    \I__2140\ : CascadeMux
    port map (
            O => \N__12533\,
            I => \N__12530\
        );

    \I__2139\ : InMux
    port map (
            O => \N__12530\,
            I => \N__12527\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__12527\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_15\
        );

    \I__2137\ : CascadeMux
    port map (
            O => \N__12524\,
            I => \N__12521\
        );

    \I__2136\ : InMux
    port map (
            O => \N__12521\,
            I => \N__12518\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__12518\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_16\
        );

    \I__2134\ : CascadeMux
    port map (
            O => \N__12515\,
            I => \N__12512\
        );

    \I__2133\ : InMux
    port map (
            O => \N__12512\,
            I => \N__12509\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__12509\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_17\
        );

    \I__2131\ : CascadeMux
    port map (
            O => \N__12506\,
            I => \N__12503\
        );

    \I__2130\ : InMux
    port map (
            O => \N__12503\,
            I => \N__12500\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__12500\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_18\
        );

    \I__2128\ : InMux
    port map (
            O => \N__12497\,
            I => \N__12494\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__12494\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_3\
        );

    \I__2126\ : CascadeMux
    port map (
            O => \N__12491\,
            I => \N__12488\
        );

    \I__2125\ : InMux
    port map (
            O => \N__12488\,
            I => \N__12485\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__12485\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_3\
        );

    \I__2123\ : InMux
    port map (
            O => \N__12482\,
            I => \N__12479\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__12479\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_4\
        );

    \I__2121\ : CascadeMux
    port map (
            O => \N__12476\,
            I => \N__12473\
        );

    \I__2120\ : InMux
    port map (
            O => \N__12473\,
            I => \N__12470\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__12470\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_4\
        );

    \I__2118\ : InMux
    port map (
            O => \N__12467\,
            I => \N__12464\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__12464\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_5\
        );

    \I__2116\ : CascadeMux
    port map (
            O => \N__12461\,
            I => \N__12458\
        );

    \I__2115\ : InMux
    port map (
            O => \N__12458\,
            I => \N__12455\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__12455\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_5\
        );

    \I__2113\ : InMux
    port map (
            O => \N__12452\,
            I => \N__12449\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__12449\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_6\
        );

    \I__2111\ : CascadeMux
    port map (
            O => \N__12446\,
            I => \N__12443\
        );

    \I__2110\ : InMux
    port map (
            O => \N__12443\,
            I => \N__12440\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__12440\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_6\
        );

    \I__2108\ : InMux
    port map (
            O => \N__12437\,
            I => \N__12434\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__12434\,
            I => \N__12431\
        );

    \I__2106\ : Odrv4
    port map (
            O => \N__12431\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_7\
        );

    \I__2105\ : CascadeMux
    port map (
            O => \N__12428\,
            I => \N__12425\
        );

    \I__2104\ : InMux
    port map (
            O => \N__12425\,
            I => \N__12422\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__12422\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_7\
        );

    \I__2102\ : InMux
    port map (
            O => \N__12419\,
            I => \N__12416\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__12416\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_8\
        );

    \I__2100\ : CascadeMux
    port map (
            O => \N__12413\,
            I => \N__12410\
        );

    \I__2099\ : InMux
    port map (
            O => \N__12410\,
            I => \N__12407\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__12407\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_8\
        );

    \I__2097\ : InMux
    port map (
            O => \N__12404\,
            I => \N__12401\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__12401\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_9\
        );

    \I__2095\ : CascadeMux
    port map (
            O => \N__12398\,
            I => \N__12395\
        );

    \I__2094\ : InMux
    port map (
            O => \N__12395\,
            I => \N__12392\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__12392\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_9\
        );

    \I__2092\ : CascadeMux
    port map (
            O => \N__12389\,
            I => \N__12386\
        );

    \I__2091\ : InMux
    port map (
            O => \N__12386\,
            I => \N__12383\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__12383\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_10\
        );

    \I__2089\ : InMux
    port map (
            O => \N__12380\,
            I => \N__12375\
        );

    \I__2088\ : InMux
    port map (
            O => \N__12379\,
            I => \N__12372\
        );

    \I__2087\ : InMux
    port map (
            O => \N__12378\,
            I => \N__12369\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__12375\,
            I => \N__12364\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__12372\,
            I => \N__12364\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__12369\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__2083\ : Odrv4
    port map (
            O => \N__12364\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__2082\ : InMux
    port map (
            O => \N__12359\,
            I => \N__12355\
        );

    \I__2081\ : InMux
    port map (
            O => \N__12358\,
            I => \N__12352\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__12355\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__12352\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__2078\ : InMux
    port map (
            O => \N__12347\,
            I => \N__12341\
        );

    \I__2077\ : InMux
    port map (
            O => \N__12346\,
            I => \N__12341\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__12341\,
            I => \N__12336\
        );

    \I__2075\ : InMux
    port map (
            O => \N__12340\,
            I => \N__12333\
        );

    \I__2074\ : InMux
    port map (
            O => \N__12339\,
            I => \N__12330\
        );

    \I__2073\ : Odrv4
    port map (
            O => \N__12336\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__12333\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__12330\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__2070\ : InMux
    port map (
            O => \N__12323\,
            I => \N__12318\
        );

    \I__2069\ : InMux
    port map (
            O => \N__12322\,
            I => \N__12315\
        );

    \I__2068\ : InMux
    port map (
            O => \N__12321\,
            I => \N__12311\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__12318\,
            I => \N__12308\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__12315\,
            I => \N__12305\
        );

    \I__2065\ : InMux
    port map (
            O => \N__12314\,
            I => \N__12302\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__12311\,
            I => \N__12295\
        );

    \I__2063\ : Span4Mux_v
    port map (
            O => \N__12308\,
            I => \N__12295\
        );

    \I__2062\ : Span4Mux_h
    port map (
            O => \N__12305\,
            I => \N__12295\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__12302\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__2060\ : Odrv4
    port map (
            O => \N__12295\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__2059\ : CascadeMux
    port map (
            O => \N__12290\,
            I => \N__12287\
        );

    \I__2058\ : InMux
    port map (
            O => \N__12287\,
            I => \N__12281\
        );

    \I__2057\ : InMux
    port map (
            O => \N__12286\,
            I => \N__12278\
        );

    \I__2056\ : InMux
    port map (
            O => \N__12285\,
            I => \N__12272\
        );

    \I__2055\ : InMux
    port map (
            O => \N__12284\,
            I => \N__12272\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__12281\,
            I => \N__12267\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__12278\,
            I => \N__12267\
        );

    \I__2052\ : InMux
    port map (
            O => \N__12277\,
            I => \N__12264\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__12272\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__2050\ : Odrv4
    port map (
            O => \N__12267\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__12264\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__2048\ : InMux
    port map (
            O => \N__12257\,
            I => \N__12253\
        );

    \I__2047\ : InMux
    port map (
            O => \N__12256\,
            I => \N__12250\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__12253\,
            I => \phase_controller_inst1.N_107\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__12250\,
            I => \phase_controller_inst1.N_107\
        );

    \I__2044\ : CascadeMux
    port map (
            O => \N__12245\,
            I => \N__12238\
        );

    \I__2043\ : CascadeMux
    port map (
            O => \N__12244\,
            I => \N__12235\
        );

    \I__2042\ : CascadeMux
    port map (
            O => \N__12243\,
            I => \N__12232\
        );

    \I__2041\ : CascadeMux
    port map (
            O => \N__12242\,
            I => \N__12217\
        );

    \I__2040\ : CascadeMux
    port map (
            O => \N__12241\,
            I => \N__12214\
        );

    \I__2039\ : InMux
    port map (
            O => \N__12238\,
            I => \N__12199\
        );

    \I__2038\ : InMux
    port map (
            O => \N__12235\,
            I => \N__12199\
        );

    \I__2037\ : InMux
    port map (
            O => \N__12232\,
            I => \N__12199\
        );

    \I__2036\ : InMux
    port map (
            O => \N__12231\,
            I => \N__12199\
        );

    \I__2035\ : InMux
    port map (
            O => \N__12230\,
            I => \N__12199\
        );

    \I__2034\ : InMux
    port map (
            O => \N__12229\,
            I => \N__12199\
        );

    \I__2033\ : InMux
    port map (
            O => \N__12228\,
            I => \N__12199\
        );

    \I__2032\ : CascadeMux
    port map (
            O => \N__12227\,
            I => \N__12196\
        );

    \I__2031\ : CascadeMux
    port map (
            O => \N__12226\,
            I => \N__12193\
        );

    \I__2030\ : CascadeMux
    port map (
            O => \N__12225\,
            I => \N__12190\
        );

    \I__2029\ : CascadeMux
    port map (
            O => \N__12224\,
            I => \N__12187\
        );

    \I__2028\ : CascadeMux
    port map (
            O => \N__12223\,
            I => \N__12180\
        );

    \I__2027\ : CascadeMux
    port map (
            O => \N__12222\,
            I => \N__12177\
        );

    \I__2026\ : CascadeMux
    port map (
            O => \N__12221\,
            I => \N__12174\
        );

    \I__2025\ : CascadeMux
    port map (
            O => \N__12220\,
            I => \N__12171\
        );

    \I__2024\ : InMux
    port map (
            O => \N__12217\,
            I => \N__12164\
        );

    \I__2023\ : InMux
    port map (
            O => \N__12214\,
            I => \N__12164\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__12199\,
            I => \N__12161\
        );

    \I__2021\ : InMux
    port map (
            O => \N__12196\,
            I => \N__12144\
        );

    \I__2020\ : InMux
    port map (
            O => \N__12193\,
            I => \N__12144\
        );

    \I__2019\ : InMux
    port map (
            O => \N__12190\,
            I => \N__12144\
        );

    \I__2018\ : InMux
    port map (
            O => \N__12187\,
            I => \N__12144\
        );

    \I__2017\ : InMux
    port map (
            O => \N__12186\,
            I => \N__12144\
        );

    \I__2016\ : InMux
    port map (
            O => \N__12185\,
            I => \N__12144\
        );

    \I__2015\ : InMux
    port map (
            O => \N__12184\,
            I => \N__12144\
        );

    \I__2014\ : InMux
    port map (
            O => \N__12183\,
            I => \N__12144\
        );

    \I__2013\ : InMux
    port map (
            O => \N__12180\,
            I => \N__12137\
        );

    \I__2012\ : InMux
    port map (
            O => \N__12177\,
            I => \N__12137\
        );

    \I__2011\ : InMux
    port map (
            O => \N__12174\,
            I => \N__12137\
        );

    \I__2010\ : InMux
    port map (
            O => \N__12171\,
            I => \N__12134\
        );

    \I__2009\ : InMux
    port map (
            O => \N__12170\,
            I => \N__12131\
        );

    \I__2008\ : InMux
    port map (
            O => \N__12169\,
            I => \N__12128\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__12164\,
            I => \N__12124\
        );

    \I__2006\ : Sp12to4
    port map (
            O => \N__12161\,
            I => \N__12115\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__12144\,
            I => \N__12115\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__12137\,
            I => \N__12115\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__12134\,
            I => \N__12115\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__12131\,
            I => \N__12110\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__12128\,
            I => \N__12110\
        );

    \I__2000\ : InMux
    port map (
            O => \N__12127\,
            I => \N__12107\
        );

    \I__1999\ : Span4Mux_h
    port map (
            O => \N__12124\,
            I => \N__12104\
        );

    \I__1998\ : Span12Mux_v
    port map (
            O => \N__12115\,
            I => \N__12101\
        );

    \I__1997\ : Span4Mux_h
    port map (
            O => \N__12110\,
            I => \N__12098\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__12107\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__1995\ : Odrv4
    port map (
            O => \N__12104\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__1994\ : Odrv12
    port map (
            O => \N__12101\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__1993\ : Odrv4
    port map (
            O => \N__12098\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__1992\ : InMux
    port map (
            O => \N__12089\,
            I => \N__12086\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__12086\,
            I => \N__12083\
        );

    \I__1990\ : Odrv4
    port map (
            O => \N__12083\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_1\
        );

    \I__1989\ : CascadeMux
    port map (
            O => \N__12080\,
            I => \N__12077\
        );

    \I__1988\ : InMux
    port map (
            O => \N__12077\,
            I => \N__12074\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__12074\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_1\
        );

    \I__1986\ : InMux
    port map (
            O => \N__12071\,
            I => \N__12068\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__12068\,
            I => \N__12065\
        );

    \I__1984\ : Span4Mux_h
    port map (
            O => \N__12065\,
            I => \N__12062\
        );

    \I__1983\ : Odrv4
    port map (
            O => \N__12062\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_2\
        );

    \I__1982\ : CascadeMux
    port map (
            O => \N__12059\,
            I => \N__12056\
        );

    \I__1981\ : InMux
    port map (
            O => \N__12056\,
            I => \N__12053\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__12053\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_2\
        );

    \I__1979\ : InMux
    port map (
            O => \N__12050\,
            I => \N__12047\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__12047\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_18\
        );

    \I__1977\ : CEMux
    port map (
            O => \N__12044\,
            I => \N__12039\
        );

    \I__1976\ : CEMux
    port map (
            O => \N__12043\,
            I => \N__12036\
        );

    \I__1975\ : CEMux
    port map (
            O => \N__12042\,
            I => \N__12032\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__12039\,
            I => \N__12027\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__12036\,
            I => \N__12027\
        );

    \I__1972\ : CEMux
    port map (
            O => \N__12035\,
            I => \N__12024\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__12032\,
            I => \N__12021\
        );

    \I__1970\ : Span4Mux_v
    port map (
            O => \N__12027\,
            I => \N__12016\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__12024\,
            I => \N__12016\
        );

    \I__1968\ : Span4Mux_h
    port map (
            O => \N__12021\,
            I => \N__12013\
        );

    \I__1967\ : Span4Mux_v
    port map (
            O => \N__12016\,
            I => \N__12010\
        );

    \I__1966\ : Span4Mux_s3_h
    port map (
            O => \N__12013\,
            I => \N__12007\
        );

    \I__1965\ : Span4Mux_s0_v
    port map (
            O => \N__12010\,
            I => \N__12004\
        );

    \I__1964\ : Odrv4
    port map (
            O => \N__12007\,
            I => \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__1963\ : Odrv4
    port map (
            O => \N__12004\,
            I => \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__1962\ : InMux
    port map (
            O => \N__11999\,
            I => \N__11996\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__11996\,
            I => \N__11993\
        );

    \I__1960\ : Span4Mux_h
    port map (
            O => \N__11993\,
            I => \N__11988\
        );

    \I__1959\ : InMux
    port map (
            O => \N__11992\,
            I => \N__11985\
        );

    \I__1958\ : InMux
    port map (
            O => \N__11991\,
            I => \N__11982\
        );

    \I__1957\ : Odrv4
    port map (
            O => \N__11988\,
            I => \phase_controller_slave.stoper_hc.time_passed11\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__11985\,
            I => \phase_controller_slave.stoper_hc.time_passed11\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__11982\,
            I => \phase_controller_slave.stoper_hc.time_passed11\
        );

    \I__1954\ : CascadeMux
    port map (
            O => \N__11975\,
            I => \N__11972\
        );

    \I__1953\ : InMux
    port map (
            O => \N__11972\,
            I => \N__11969\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__11969\,
            I => \phase_controller_slave.stoper_hc.time_passed_1_sqmuxa\
        );

    \I__1951\ : InMux
    port map (
            O => \N__11966\,
            I => \N__11959\
        );

    \I__1950\ : InMux
    port map (
            O => \N__11965\,
            I => \N__11954\
        );

    \I__1949\ : InMux
    port map (
            O => \N__11964\,
            I => \N__11954\
        );

    \I__1948\ : InMux
    port map (
            O => \N__11963\,
            I => \N__11949\
        );

    \I__1947\ : InMux
    port map (
            O => \N__11962\,
            I => \N__11949\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__11959\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__11954\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__11949\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__1943\ : CascadeMux
    port map (
            O => \N__11942\,
            I => \N__11929\
        );

    \I__1942\ : CascadeMux
    port map (
            O => \N__11941\,
            I => \N__11925\
        );

    \I__1941\ : CascadeMux
    port map (
            O => \N__11940\,
            I => \N__11922\
        );

    \I__1940\ : CascadeMux
    port map (
            O => \N__11939\,
            I => \N__11919\
        );

    \I__1939\ : CascadeMux
    port map (
            O => \N__11938\,
            I => \N__11916\
        );

    \I__1938\ : CascadeMux
    port map (
            O => \N__11937\,
            I => \N__11908\
        );

    \I__1937\ : CascadeMux
    port map (
            O => \N__11936\,
            I => \N__11905\
        );

    \I__1936\ : CascadeMux
    port map (
            O => \N__11935\,
            I => \N__11898\
        );

    \I__1935\ : CascadeMux
    port map (
            O => \N__11934\,
            I => \N__11895\
        );

    \I__1934\ : CascadeMux
    port map (
            O => \N__11933\,
            I => \N__11892\
        );

    \I__1933\ : CascadeMux
    port map (
            O => \N__11932\,
            I => \N__11889\
        );

    \I__1932\ : InMux
    port map (
            O => \N__11929\,
            I => \N__11883\
        );

    \I__1931\ : InMux
    port map (
            O => \N__11928\,
            I => \N__11883\
        );

    \I__1930\ : InMux
    port map (
            O => \N__11925\,
            I => \N__11866\
        );

    \I__1929\ : InMux
    port map (
            O => \N__11922\,
            I => \N__11866\
        );

    \I__1928\ : InMux
    port map (
            O => \N__11919\,
            I => \N__11866\
        );

    \I__1927\ : InMux
    port map (
            O => \N__11916\,
            I => \N__11866\
        );

    \I__1926\ : InMux
    port map (
            O => \N__11915\,
            I => \N__11866\
        );

    \I__1925\ : InMux
    port map (
            O => \N__11914\,
            I => \N__11866\
        );

    \I__1924\ : InMux
    port map (
            O => \N__11913\,
            I => \N__11866\
        );

    \I__1923\ : InMux
    port map (
            O => \N__11912\,
            I => \N__11861\
        );

    \I__1922\ : InMux
    port map (
            O => \N__11911\,
            I => \N__11861\
        );

    \I__1921\ : InMux
    port map (
            O => \N__11908\,
            I => \N__11856\
        );

    \I__1920\ : InMux
    port map (
            O => \N__11905\,
            I => \N__11856\
        );

    \I__1919\ : InMux
    port map (
            O => \N__11904\,
            I => \N__11839\
        );

    \I__1918\ : InMux
    port map (
            O => \N__11903\,
            I => \N__11839\
        );

    \I__1917\ : InMux
    port map (
            O => \N__11902\,
            I => \N__11839\
        );

    \I__1916\ : InMux
    port map (
            O => \N__11901\,
            I => \N__11839\
        );

    \I__1915\ : InMux
    port map (
            O => \N__11898\,
            I => \N__11839\
        );

    \I__1914\ : InMux
    port map (
            O => \N__11895\,
            I => \N__11839\
        );

    \I__1913\ : InMux
    port map (
            O => \N__11892\,
            I => \N__11839\
        );

    \I__1912\ : InMux
    port map (
            O => \N__11889\,
            I => \N__11839\
        );

    \I__1911\ : CascadeMux
    port map (
            O => \N__11888\,
            I => \N__11836\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__11883\,
            I => \N__11833\
        );

    \I__1909\ : InMux
    port map (
            O => \N__11882\,
            I => \N__11828\
        );

    \I__1908\ : InMux
    port map (
            O => \N__11881\,
            I => \N__11828\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__11866\,
            I => \N__11825\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__11861\,
            I => \N__11820\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__11856\,
            I => \N__11820\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__11839\,
            I => \N__11817\
        );

    \I__1903\ : InMux
    port map (
            O => \N__11836\,
            I => \N__11814\
        );

    \I__1902\ : Span4Mux_v
    port map (
            O => \N__11833\,
            I => \N__11809\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__11828\,
            I => \N__11809\
        );

    \I__1900\ : Span4Mux_h
    port map (
            O => \N__11825\,
            I => \N__11806\
        );

    \I__1899\ : Span4Mux_h
    port map (
            O => \N__11820\,
            I => \N__11803\
        );

    \I__1898\ : Span4Mux_h
    port map (
            O => \N__11817\,
            I => \N__11800\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__11814\,
            I => \N__11795\
        );

    \I__1896\ : Span4Mux_v
    port map (
            O => \N__11809\,
            I => \N__11795\
        );

    \I__1895\ : Odrv4
    port map (
            O => \N__11806\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__1894\ : Odrv4
    port map (
            O => \N__11803\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__1893\ : Odrv4
    port map (
            O => \N__11800\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__1892\ : Odrv4
    port map (
            O => \N__11795\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__1891\ : InMux
    port map (
            O => \N__11786\,
            I => \N__11783\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__11783\,
            I => \N__11780\
        );

    \I__1889\ : Odrv4
    port map (
            O => \N__11780\,
            I => \phase_controller_inst1.N_110\
        );

    \I__1888\ : InMux
    port map (
            O => \N__11777\,
            I => \N__11774\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__11774\,
            I => \phase_controller_inst1.N_112\
        );

    \I__1886\ : InMux
    port map (
            O => \N__11771\,
            I => \N__11768\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__11768\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_13\
        );

    \I__1884\ : InMux
    port map (
            O => \N__11765\,
            I => \N__11762\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__11762\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_10\
        );

    \I__1882\ : InMux
    port map (
            O => \N__11759\,
            I => \N__11756\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__11756\,
            I => \N__11753\
        );

    \I__1880\ : Odrv4
    port map (
            O => \N__11753\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_12\
        );

    \I__1879\ : InMux
    port map (
            O => \N__11750\,
            I => \N__11746\
        );

    \I__1878\ : InMux
    port map (
            O => \N__11749\,
            I => \N__11743\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__11746\,
            I => \N__11739\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__11743\,
            I => \N__11736\
        );

    \I__1875\ : InMux
    port map (
            O => \N__11742\,
            I => \N__11733\
        );

    \I__1874\ : Odrv12
    port map (
            O => \N__11739\,
            I => \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_0Z0Z_6\
        );

    \I__1873\ : Odrv4
    port map (
            O => \N__11736\,
            I => \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_0Z0Z_6\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__11733\,
            I => \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_0Z0Z_6\
        );

    \I__1871\ : InMux
    port map (
            O => \N__11726\,
            I => \N__11723\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__11723\,
            I => \N__11720\
        );

    \I__1869\ : Span12Mux_s5_v
    port map (
            O => \N__11720\,
            I => \N__11717\
        );

    \I__1868\ : Odrv12
    port map (
            O => \N__11717\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_9\
        );

    \I__1867\ : CascadeMux
    port map (
            O => \N__11714\,
            I => \N__11709\
        );

    \I__1866\ : CascadeMux
    port map (
            O => \N__11713\,
            I => \N__11703\
        );

    \I__1865\ : InMux
    port map (
            O => \N__11712\,
            I => \N__11696\
        );

    \I__1864\ : InMux
    port map (
            O => \N__11709\,
            I => \N__11687\
        );

    \I__1863\ : InMux
    port map (
            O => \N__11708\,
            I => \N__11687\
        );

    \I__1862\ : InMux
    port map (
            O => \N__11707\,
            I => \N__11687\
        );

    \I__1861\ : InMux
    port map (
            O => \N__11706\,
            I => \N__11687\
        );

    \I__1860\ : InMux
    port map (
            O => \N__11703\,
            I => \N__11676\
        );

    \I__1859\ : InMux
    port map (
            O => \N__11702\,
            I => \N__11676\
        );

    \I__1858\ : InMux
    port map (
            O => \N__11701\,
            I => \N__11676\
        );

    \I__1857\ : InMux
    port map (
            O => \N__11700\,
            I => \N__11676\
        );

    \I__1856\ : InMux
    port map (
            O => \N__11699\,
            I => \N__11676\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__11696\,
            I => \N__11671\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__11687\,
            I => \N__11671\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__11676\,
            I => \N__11668\
        );

    \I__1852\ : Odrv12
    port map (
            O => \N__11671\,
            I => \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_o2Z0Z_9\
        );

    \I__1851\ : Odrv4
    port map (
            O => \N__11668\,
            I => \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_o2Z0Z_9\
        );

    \I__1850\ : InMux
    port map (
            O => \N__11663\,
            I => \N__11660\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__11660\,
            I => \N__11657\
        );

    \I__1848\ : Span4Mux_v
    port map (
            O => \N__11657\,
            I => \N__11654\
        );

    \I__1847\ : Odrv4
    port map (
            O => \N__11654\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_11\
        );

    \I__1846\ : InMux
    port map (
            O => \N__11651\,
            I => \N__11645\
        );

    \I__1845\ : InMux
    port map (
            O => \N__11650\,
            I => \N__11645\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__11645\,
            I => \N__11640\
        );

    \I__1843\ : InMux
    port map (
            O => \N__11644\,
            I => \N__11635\
        );

    \I__1842\ : InMux
    port map (
            O => \N__11643\,
            I => \N__11635\
        );

    \I__1841\ : Sp12to4
    port map (
            O => \N__11640\,
            I => \N__11631\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__11635\,
            I => \N__11628\
        );

    \I__1839\ : InMux
    port map (
            O => \N__11634\,
            I => \N__11625\
        );

    \I__1838\ : Odrv12
    port map (
            O => \N__11631\,
            I => \phase_controller_inst1.stoper_hc.target_time_6_i_o2Z0Z_15\
        );

    \I__1837\ : Odrv12
    port map (
            O => \N__11628\,
            I => \phase_controller_inst1.stoper_hc.target_time_6_i_o2Z0Z_15\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__11625\,
            I => \phase_controller_inst1.stoper_hc.target_time_6_i_o2Z0Z_15\
        );

    \I__1835\ : InMux
    port map (
            O => \N__11618\,
            I => \N__11615\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__11615\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_14\
        );

    \I__1833\ : InMux
    port map (
            O => \N__11612\,
            I => \N__11609\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__11609\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_16\
        );

    \I__1831\ : InMux
    port map (
            O => \N__11606\,
            I => \N__11603\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__11603\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_19\
        );

    \I__1829\ : InMux
    port map (
            O => \N__11600\,
            I => \N__11597\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__11597\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_17\
        );

    \I__1827\ : InMux
    port map (
            O => \N__11594\,
            I => \N__11591\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__11591\,
            I => \N__11588\
        );

    \I__1825\ : Span4Mux_h
    port map (
            O => \N__11588\,
            I => \N__11585\
        );

    \I__1824\ : Odrv4
    port map (
            O => \N__11585\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_5\
        );

    \I__1823\ : InMux
    port map (
            O => \N__11582\,
            I => \N__11579\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__11579\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_1\
        );

    \I__1821\ : InMux
    port map (
            O => \N__11576\,
            I => \N__11573\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__11573\,
            I => \N__11570\
        );

    \I__1819\ : Span4Mux_h
    port map (
            O => \N__11570\,
            I => \N__11567\
        );

    \I__1818\ : Odrv4
    port map (
            O => \N__11567\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_7\
        );

    \I__1817\ : InMux
    port map (
            O => \N__11564\,
            I => \N__11561\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__11561\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_6\
        );

    \I__1815\ : InMux
    port map (
            O => \N__11558\,
            I => \N__11550\
        );

    \I__1814\ : InMux
    port map (
            O => \N__11557\,
            I => \N__11550\
        );

    \I__1813\ : InMux
    port map (
            O => \N__11556\,
            I => \N__11545\
        );

    \I__1812\ : InMux
    port map (
            O => \N__11555\,
            I => \N__11545\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__11550\,
            I => \N__11542\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__11545\,
            I => \N__11539\
        );

    \I__1809\ : Odrv12
    port map (
            O => \N__11542\,
            I => \phase_controller_inst1.stoper_hc.N_122\
        );

    \I__1808\ : Odrv4
    port map (
            O => \N__11539\,
            I => \phase_controller_inst1.stoper_hc.N_122\
        );

    \I__1807\ : CascadeMux
    port map (
            O => \N__11534\,
            I => \N__11531\
        );

    \I__1806\ : InMux
    port map (
            O => \N__11531\,
            I => \N__11528\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__11528\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_2\
        );

    \I__1804\ : InMux
    port map (
            O => \N__11525\,
            I => \N__11522\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__11522\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_4\
        );

    \I__1802\ : InMux
    port map (
            O => \N__11519\,
            I => \N__11501\
        );

    \I__1801\ : InMux
    port map (
            O => \N__11518\,
            I => \N__11501\
        );

    \I__1800\ : InMux
    port map (
            O => \N__11517\,
            I => \N__11501\
        );

    \I__1799\ : InMux
    port map (
            O => \N__11516\,
            I => \N__11501\
        );

    \I__1798\ : InMux
    port map (
            O => \N__11515\,
            I => \N__11501\
        );

    \I__1797\ : InMux
    port map (
            O => \N__11514\,
            I => \N__11501\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__11501\,
            I => \N__11498\
        );

    \I__1795\ : Span4Mux_v
    port map (
            O => \N__11498\,
            I => \N__11495\
        );

    \I__1794\ : Span4Mux_v
    port map (
            O => \N__11495\,
            I => \N__11486\
        );

    \I__1793\ : InMux
    port map (
            O => \N__11494\,
            I => \N__11473\
        );

    \I__1792\ : InMux
    port map (
            O => \N__11493\,
            I => \N__11473\
        );

    \I__1791\ : InMux
    port map (
            O => \N__11492\,
            I => \N__11473\
        );

    \I__1790\ : InMux
    port map (
            O => \N__11491\,
            I => \N__11473\
        );

    \I__1789\ : InMux
    port map (
            O => \N__11490\,
            I => \N__11473\
        );

    \I__1788\ : InMux
    port map (
            O => \N__11489\,
            I => \N__11473\
        );

    \I__1787\ : Odrv4
    port map (
            O => \N__11486\,
            I => \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a3_0Z0Z_6\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__11473\,
            I => \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a3_0Z0Z_6\
        );

    \I__1785\ : InMux
    port map (
            O => \N__11468\,
            I => \N__11464\
        );

    \I__1784\ : InMux
    port map (
            O => \N__11467\,
            I => \N__11461\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__11464\,
            I => \N__11458\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__11461\,
            I => \N__11455\
        );

    \I__1781\ : Odrv12
    port map (
            O => \N__11458\,
            I => \phase_controller_inst1.stoper_hc.N_144\
        );

    \I__1780\ : Odrv4
    port map (
            O => \N__11455\,
            I => \phase_controller_inst1.stoper_hc.N_144\
        );

    \I__1779\ : InMux
    port map (
            O => \N__11450\,
            I => \N__11447\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__11447\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_3\
        );

    \I__1777\ : CascadeMux
    port map (
            O => \N__11444\,
            I => \N__11435\
        );

    \I__1776\ : InMux
    port map (
            O => \N__11443\,
            I => \N__11429\
        );

    \I__1775\ : InMux
    port map (
            O => \N__11442\,
            I => \N__11429\
        );

    \I__1774\ : InMux
    port map (
            O => \N__11441\,
            I => \N__11416\
        );

    \I__1773\ : InMux
    port map (
            O => \N__11440\,
            I => \N__11416\
        );

    \I__1772\ : InMux
    port map (
            O => \N__11439\,
            I => \N__11416\
        );

    \I__1771\ : InMux
    port map (
            O => \N__11438\,
            I => \N__11416\
        );

    \I__1770\ : InMux
    port map (
            O => \N__11435\,
            I => \N__11416\
        );

    \I__1769\ : InMux
    port map (
            O => \N__11434\,
            I => \N__11416\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__11429\,
            I => \N__11409\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__11416\,
            I => \N__11409\
        );

    \I__1766\ : CascadeMux
    port map (
            O => \N__11415\,
            I => \N__11405\
        );

    \I__1765\ : CascadeMux
    port map (
            O => \N__11414\,
            I => \N__11398\
        );

    \I__1764\ : Span4Mux_v
    port map (
            O => \N__11409\,
            I => \N__11394\
        );

    \I__1763\ : InMux
    port map (
            O => \N__11408\,
            I => \N__11377\
        );

    \I__1762\ : InMux
    port map (
            O => \N__11405\,
            I => \N__11377\
        );

    \I__1761\ : InMux
    port map (
            O => \N__11404\,
            I => \N__11377\
        );

    \I__1760\ : InMux
    port map (
            O => \N__11403\,
            I => \N__11377\
        );

    \I__1759\ : InMux
    port map (
            O => \N__11402\,
            I => \N__11377\
        );

    \I__1758\ : InMux
    port map (
            O => \N__11401\,
            I => \N__11377\
        );

    \I__1757\ : InMux
    port map (
            O => \N__11398\,
            I => \N__11377\
        );

    \I__1756\ : InMux
    port map (
            O => \N__11397\,
            I => \N__11377\
        );

    \I__1755\ : Span4Mux_v
    port map (
            O => \N__11394\,
            I => \N__11372\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__11377\,
            I => \N__11372\
        );

    \I__1753\ : Odrv4
    port map (
            O => \N__11372\,
            I => \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_o2Z0Z_6\
        );

    \I__1752\ : InMux
    port map (
            O => \N__11369\,
            I => \N__11366\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__11366\,
            I => \N__11363\
        );

    \I__1750\ : Odrv4
    port map (
            O => \N__11363\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_8\
        );

    \I__1749\ : InMux
    port map (
            O => \N__11360\,
            I => \N__11357\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__11357\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_15\
        );

    \I__1747\ : InMux
    port map (
            O => \N__11354\,
            I => \N__11351\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__11351\,
            I => \phase_controller_inst1.stoper_hc.target_time_6_f0_0_a2_4Z0Z_3\
        );

    \I__1745\ : CascadeMux
    port map (
            O => \N__11348\,
            I => \phase_controller_inst1.stoper_hc.target_time_6_f0_0_a2_3Z0Z_3_cascade_\
        );

    \I__1744\ : CascadeMux
    port map (
            O => \N__11345\,
            I => \phase_controller_inst1.stoper_hc.N_144_cascade_\
        );

    \I__1743\ : CascadeMux
    port map (
            O => \N__11342\,
            I => \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_0Z0Z_6_cascade_\
        );

    \I__1742\ : InMux
    port map (
            O => \N__11339\,
            I => \N__11336\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__11336\,
            I => \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2Z0Z_9\
        );

    \I__1740\ : CascadeMux
    port map (
            O => \N__11333\,
            I => \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2Z0Z_9_cascade_\
        );

    \I__1739\ : CascadeMux
    port map (
            O => \N__11330\,
            I => \phase_controller_inst1.stoper_hc.target_time_6_i_o2Z0Z_15_cascade_\
        );

    \I__1738\ : InMux
    port map (
            O => \N__11327\,
            I => \N__11324\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__11324\,
            I => \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_1Z0Z_6\
        );

    \I__1736\ : CascadeMux
    port map (
            O => \N__11321\,
            I => \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_1Z0Z_6_cascade_\
        );

    \I__1735\ : InMux
    port map (
            O => \N__11318\,
            I => \N__11315\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__11315\,
            I => \N__11312\
        );

    \I__1733\ : Odrv4
    port map (
            O => \N__11312\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\
        );

    \I__1732\ : InMux
    port map (
            O => \N__11309\,
            I => \N__11306\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__11306\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\
        );

    \I__1730\ : InMux
    port map (
            O => \N__11303\,
            I => \N__11300\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__11300\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\
        );

    \I__1728\ : InMux
    port map (
            O => \N__11297\,
            I => \N__11294\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__11294\,
            I => \N__11291\
        );

    \I__1726\ : Odrv4
    port map (
            O => \N__11291\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\
        );

    \I__1725\ : InMux
    port map (
            O => \N__11288\,
            I => \N__11285\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__11285\,
            I => \N__11282\
        );

    \I__1723\ : Odrv4
    port map (
            O => \N__11282\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\
        );

    \I__1722\ : InMux
    port map (
            O => \N__11279\,
            I => \N__11276\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__11276\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\
        );

    \I__1720\ : CEMux
    port map (
            O => \N__11273\,
            I => \N__11270\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__11270\,
            I => \N__11266\
        );

    \I__1718\ : CEMux
    port map (
            O => \N__11269\,
            I => \N__11263\
        );

    \I__1717\ : Span4Mux_v
    port map (
            O => \N__11266\,
            I => \N__11259\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__11263\,
            I => \N__11256\
        );

    \I__1715\ : CEMux
    port map (
            O => \N__11262\,
            I => \N__11253\
        );

    \I__1714\ : Span4Mux_h
    port map (
            O => \N__11259\,
            I => \N__11250\
        );

    \I__1713\ : Span4Mux_h
    port map (
            O => \N__11256\,
            I => \N__11247\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__11253\,
            I => \N__11244\
        );

    \I__1711\ : Odrv4
    port map (
            O => \N__11250\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__1710\ : Odrv4
    port map (
            O => \N__11247\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__1709\ : Odrv12
    port map (
            O => \N__11244\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__1708\ : InMux
    port map (
            O => \N__11237\,
            I => \N__11234\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__11234\,
            I => \N__11231\
        );

    \I__1706\ : Odrv4
    port map (
            O => \N__11231\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\
        );

    \I__1705\ : InMux
    port map (
            O => \N__11228\,
            I => \N__11225\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__11225\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\
        );

    \I__1703\ : InMux
    port map (
            O => \N__11222\,
            I => \N__11219\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__11219\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\
        );

    \I__1701\ : InMux
    port map (
            O => \N__11216\,
            I => \N__11213\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__11213\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\
        );

    \I__1699\ : InMux
    port map (
            O => \N__11210\,
            I => \N__11207\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__11207\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\
        );

    \I__1697\ : InMux
    port map (
            O => \N__11204\,
            I => \N__11201\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__11201\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\
        );

    \I__1695\ : InMux
    port map (
            O => \N__11198\,
            I => \N__11195\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__11195\,
            I => \N__11192\
        );

    \I__1693\ : Odrv4
    port map (
            O => \N__11192\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\
        );

    \I__1692\ : InMux
    port map (
            O => \N__11189\,
            I => \N__11186\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__11186\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\
        );

    \I__1690\ : InMux
    port map (
            O => \N__11183\,
            I => \N__11180\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__11180\,
            I => \N__11177\
        );

    \I__1688\ : Odrv4
    port map (
            O => \N__11177\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\
        );

    \I__1687\ : InMux
    port map (
            O => \N__11174\,
            I => \N__11171\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__11171\,
            I => \N__11168\
        );

    \I__1685\ : Odrv4
    port map (
            O => \N__11168\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\
        );

    \I__1684\ : InMux
    port map (
            O => \N__11165\,
            I => \N__11162\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__11162\,
            I => \N__11159\
        );

    \I__1682\ : Odrv4
    port map (
            O => \N__11159\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\
        );

    \I__1681\ : InMux
    port map (
            O => \N__11156\,
            I => \N__11153\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__11153\,
            I => \N__11150\
        );

    \I__1679\ : Odrv4
    port map (
            O => \N__11150\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\
        );

    \I__1678\ : CEMux
    port map (
            O => \N__11147\,
            I => \N__11142\
        );

    \I__1677\ : CEMux
    port map (
            O => \N__11146\,
            I => \N__11139\
        );

    \I__1676\ : CEMux
    port map (
            O => \N__11145\,
            I => \N__11136\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__11142\,
            I => \N__11133\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__11139\,
            I => \N__11130\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__11136\,
            I => \N__11127\
        );

    \I__1672\ : Span4Mux_v
    port map (
            O => \N__11133\,
            I => \N__11120\
        );

    \I__1671\ : Span4Mux_v
    port map (
            O => \N__11130\,
            I => \N__11120\
        );

    \I__1670\ : Span4Mux_h
    port map (
            O => \N__11127\,
            I => \N__11120\
        );

    \I__1669\ : Odrv4
    port map (
            O => \N__11120\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__1668\ : InMux
    port map (
            O => \N__11117\,
            I => \N__11110\
        );

    \I__1667\ : InMux
    port map (
            O => \N__11116\,
            I => \N__11110\
        );

    \I__1666\ : InMux
    port map (
            O => \N__11115\,
            I => \N__11107\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__11110\,
            I => \N__11104\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__11107\,
            I => \N__11101\
        );

    \I__1663\ : Span4Mux_v
    port map (
            O => \N__11104\,
            I => \N__11098\
        );

    \I__1662\ : Odrv4
    port map (
            O => \N__11101\,
            I => \phase_controller_inst1.stoper_tr.time_passed11\
        );

    \I__1661\ : Odrv4
    port map (
            O => \N__11098\,
            I => \phase_controller_inst1.stoper_tr.time_passed11\
        );

    \I__1660\ : CascadeMux
    port map (
            O => \N__11093\,
            I => \N__11090\
        );

    \I__1659\ : InMux
    port map (
            O => \N__11090\,
            I => \N__11087\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__11087\,
            I => \N__11084\
        );

    \I__1657\ : Odrv4
    port map (
            O => \N__11084\,
            I => \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa\
        );

    \I__1656\ : InMux
    port map (
            O => \N__11081\,
            I => \N__11077\
        );

    \I__1655\ : InMux
    port map (
            O => \N__11080\,
            I => \N__11072\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__11077\,
            I => \N__11068\
        );

    \I__1653\ : InMux
    port map (
            O => \N__11076\,
            I => \N__11063\
        );

    \I__1652\ : InMux
    port map (
            O => \N__11075\,
            I => \N__11063\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__11072\,
            I => \N__11060\
        );

    \I__1650\ : InMux
    port map (
            O => \N__11071\,
            I => \N__11057\
        );

    \I__1649\ : Span4Mux_h
    port map (
            O => \N__11068\,
            I => \N__11050\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__11063\,
            I => \N__11050\
        );

    \I__1647\ : Span4Mux_s3_h
    port map (
            O => \N__11060\,
            I => \N__11050\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__11057\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__1645\ : Odrv4
    port map (
            O => \N__11050\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__1644\ : InMux
    port map (
            O => \N__11045\,
            I => \N__11038\
        );

    \I__1643\ : InMux
    port map (
            O => \N__11044\,
            I => \N__11033\
        );

    \I__1642\ : InMux
    port map (
            O => \N__11043\,
            I => \N__11033\
        );

    \I__1641\ : InMux
    port map (
            O => \N__11042\,
            I => \N__11028\
        );

    \I__1640\ : InMux
    port map (
            O => \N__11041\,
            I => \N__11028\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__11038\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__11033\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__11028\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__1636\ : CascadeMux
    port map (
            O => \N__11021\,
            I => \N__11018\
        );

    \I__1635\ : InMux
    port map (
            O => \N__11018\,
            I => \N__11015\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__11015\,
            I => \N__11012\
        );

    \I__1633\ : Odrv4
    port map (
            O => \N__11012\,
            I => \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa\
        );

    \I__1632\ : InMux
    port map (
            O => \N__11009\,
            I => \N__11006\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__11006\,
            I => \N__11001\
        );

    \I__1630\ : InMux
    port map (
            O => \N__11005\,
            I => \N__10998\
        );

    \I__1629\ : InMux
    port map (
            O => \N__11004\,
            I => \N__10995\
        );

    \I__1628\ : Odrv4
    port map (
            O => \N__11001\,
            I => \phase_controller_inst1.stoper_hc.time_passed11\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__10998\,
            I => \phase_controller_inst1.stoper_hc.time_passed11\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__10995\,
            I => \phase_controller_inst1.stoper_hc.time_passed11\
        );

    \I__1625\ : InMux
    port map (
            O => \N__10988\,
            I => \N__10985\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__10985\,
            I => \N__10982\
        );

    \I__1623\ : Odrv4
    port map (
            O => \N__10982\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\
        );

    \I__1622\ : InMux
    port map (
            O => \N__10979\,
            I => \N__10976\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__10976\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\
        );

    \I__1620\ : InMux
    port map (
            O => \N__10973\,
            I => \N__10970\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__10970\,
            I => \N__10967\
        );

    \I__1618\ : Odrv4
    port map (
            O => \N__10967\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\
        );

    \I__1617\ : InMux
    port map (
            O => \N__10964\,
            I => \N__10961\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__10961\,
            I => \N__10958\
        );

    \I__1615\ : Odrv4
    port map (
            O => \N__10958\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\
        );

    \I__1614\ : InMux
    port map (
            O => \N__10955\,
            I => \N__10952\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__10952\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\
        );

    \I__1612\ : InMux
    port map (
            O => \N__10949\,
            I => \N__10946\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__10946\,
            I => \N__10943\
        );

    \I__1610\ : Odrv4
    port map (
            O => \N__10943\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\
        );

    \I__1609\ : InMux
    port map (
            O => \N__10940\,
            I => \N__10937\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__10937\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\
        );

    \I__1607\ : InMux
    port map (
            O => \N__10934\,
            I => \N__10931\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__10931\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\
        );

    \I__1605\ : InMux
    port map (
            O => \N__10928\,
            I => \N__10925\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__10925\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\
        );

    \I__1603\ : InMux
    port map (
            O => \N__10922\,
            I => \N__10919\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__10919\,
            I => \N__10916\
        );

    \I__1601\ : Odrv4
    port map (
            O => \N__10916\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\
        );

    \I__1600\ : InMux
    port map (
            O => \N__10913\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__1599\ : CascadeMux
    port map (
            O => \N__10910\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_\
        );

    \I__1598\ : CascadeMux
    port map (
            O => \N__10907\,
            I => \N__10904\
        );

    \I__1597\ : InMux
    port map (
            O => \N__10904\,
            I => \N__10901\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__10901\,
            I => \N__10898\
        );

    \I__1595\ : Span4Mux_s3_h
    port map (
            O => \N__10898\,
            I => \N__10895\
        );

    \I__1594\ : Odrv4
    port map (
            O => \N__10895\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\
        );

    \I__1593\ : CascadeMux
    port map (
            O => \N__10892\,
            I => \N__10876\
        );

    \I__1592\ : InMux
    port map (
            O => \N__10891\,
            I => \N__10853\
        );

    \I__1591\ : InMux
    port map (
            O => \N__10890\,
            I => \N__10853\
        );

    \I__1590\ : InMux
    port map (
            O => \N__10889\,
            I => \N__10853\
        );

    \I__1589\ : InMux
    port map (
            O => \N__10888\,
            I => \N__10853\
        );

    \I__1588\ : InMux
    port map (
            O => \N__10887\,
            I => \N__10853\
        );

    \I__1587\ : InMux
    port map (
            O => \N__10886\,
            I => \N__10853\
        );

    \I__1586\ : InMux
    port map (
            O => \N__10885\,
            I => \N__10853\
        );

    \I__1585\ : InMux
    port map (
            O => \N__10884\,
            I => \N__10853\
        );

    \I__1584\ : InMux
    port map (
            O => \N__10883\,
            I => \N__10846\
        );

    \I__1583\ : InMux
    port map (
            O => \N__10882\,
            I => \N__10846\
        );

    \I__1582\ : InMux
    port map (
            O => \N__10881\,
            I => \N__10846\
        );

    \I__1581\ : CascadeMux
    port map (
            O => \N__10880\,
            I => \N__10843\
        );

    \I__1580\ : InMux
    port map (
            O => \N__10879\,
            I => \N__10825\
        );

    \I__1579\ : InMux
    port map (
            O => \N__10876\,
            I => \N__10825\
        );

    \I__1578\ : InMux
    port map (
            O => \N__10875\,
            I => \N__10825\
        );

    \I__1577\ : InMux
    port map (
            O => \N__10874\,
            I => \N__10825\
        );

    \I__1576\ : InMux
    port map (
            O => \N__10873\,
            I => \N__10825\
        );

    \I__1575\ : InMux
    port map (
            O => \N__10872\,
            I => \N__10825\
        );

    \I__1574\ : InMux
    port map (
            O => \N__10871\,
            I => \N__10825\
        );

    \I__1573\ : InMux
    port map (
            O => \N__10870\,
            I => \N__10825\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__10853\,
            I => \N__10822\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__10846\,
            I => \N__10819\
        );

    \I__1570\ : InMux
    port map (
            O => \N__10843\,
            I => \N__10811\
        );

    \I__1569\ : InMux
    port map (
            O => \N__10842\,
            I => \N__10811\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__10825\,
            I => \N__10806\
        );

    \I__1567\ : Span4Mux_h
    port map (
            O => \N__10822\,
            I => \N__10806\
        );

    \I__1566\ : Span4Mux_v
    port map (
            O => \N__10819\,
            I => \N__10803\
        );

    \I__1565\ : InMux
    port map (
            O => \N__10818\,
            I => \N__10800\
        );

    \I__1564\ : InMux
    port map (
            O => \N__10817\,
            I => \N__10797\
        );

    \I__1563\ : InMux
    port map (
            O => \N__10816\,
            I => \N__10794\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__10811\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__1561\ : Odrv4
    port map (
            O => \N__10806\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__1560\ : Odrv4
    port map (
            O => \N__10803\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__10800\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__10797\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__10794\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__1556\ : InMux
    port map (
            O => \N__10781\,
            I => \N__10746\
        );

    \I__1555\ : InMux
    port map (
            O => \N__10780\,
            I => \N__10746\
        );

    \I__1554\ : InMux
    port map (
            O => \N__10779\,
            I => \N__10746\
        );

    \I__1553\ : InMux
    port map (
            O => \N__10778\,
            I => \N__10746\
        );

    \I__1552\ : InMux
    port map (
            O => \N__10777\,
            I => \N__10746\
        );

    \I__1551\ : InMux
    port map (
            O => \N__10776\,
            I => \N__10746\
        );

    \I__1550\ : InMux
    port map (
            O => \N__10775\,
            I => \N__10746\
        );

    \I__1549\ : InMux
    port map (
            O => \N__10774\,
            I => \N__10746\
        );

    \I__1548\ : InMux
    port map (
            O => \N__10773\,
            I => \N__10729\
        );

    \I__1547\ : InMux
    port map (
            O => \N__10772\,
            I => \N__10729\
        );

    \I__1546\ : InMux
    port map (
            O => \N__10771\,
            I => \N__10729\
        );

    \I__1545\ : InMux
    port map (
            O => \N__10770\,
            I => \N__10729\
        );

    \I__1544\ : InMux
    port map (
            O => \N__10769\,
            I => \N__10729\
        );

    \I__1543\ : InMux
    port map (
            O => \N__10768\,
            I => \N__10729\
        );

    \I__1542\ : InMux
    port map (
            O => \N__10767\,
            I => \N__10729\
        );

    \I__1541\ : InMux
    port map (
            O => \N__10766\,
            I => \N__10729\
        );

    \I__1540\ : InMux
    port map (
            O => \N__10765\,
            I => \N__10722\
        );

    \I__1539\ : InMux
    port map (
            O => \N__10764\,
            I => \N__10722\
        );

    \I__1538\ : InMux
    port map (
            O => \N__10763\,
            I => \N__10722\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__10746\,
            I => \N__10715\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__10729\,
            I => \N__10715\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__10722\,
            I => \N__10712\
        );

    \I__1534\ : InMux
    port map (
            O => \N__10721\,
            I => \N__10704\
        );

    \I__1533\ : InMux
    port map (
            O => \N__10720\,
            I => \N__10704\
        );

    \I__1532\ : Span4Mux_v
    port map (
            O => \N__10715\,
            I => \N__10699\
        );

    \I__1531\ : Span4Mux_v
    port map (
            O => \N__10712\,
            I => \N__10699\
        );

    \I__1530\ : InMux
    port map (
            O => \N__10711\,
            I => \N__10696\
        );

    \I__1529\ : InMux
    port map (
            O => \N__10710\,
            I => \N__10693\
        );

    \I__1528\ : InMux
    port map (
            O => \N__10709\,
            I => \N__10690\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__10704\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__1526\ : Odrv4
    port map (
            O => \N__10699\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__10696\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__10693\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__10690\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__1522\ : InMux
    port map (
            O => \N__10679\,
            I => \N__10676\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__10676\,
            I => \N__10673\
        );

    \I__1520\ : Glb2LocalMux
    port map (
            O => \N__10673\,
            I => \N__10670\
        );

    \I__1519\ : GlobalMux
    port map (
            O => \N__10670\,
            I => clk_12mhz
        );

    \I__1518\ : IoInMux
    port map (
            O => \N__10667\,
            I => \N__10664\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__10664\,
            I => \N__10661\
        );

    \I__1516\ : Span4Mux_s0_v
    port map (
            O => \N__10661\,
            I => \N__10658\
        );

    \I__1515\ : Span4Mux_h
    port map (
            O => \N__10658\,
            I => \N__10655\
        );

    \I__1514\ : Odrv4
    port map (
            O => \N__10655\,
            I => \GB_BUFFER_clk_12mhz_THRU_CO\
        );

    \I__1513\ : InMux
    port map (
            O => \N__10652\,
            I => \N__10649\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__10649\,
            I => \N__10646\
        );

    \I__1511\ : Odrv4
    port map (
            O => \N__10646\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\
        );

    \I__1510\ : InMux
    port map (
            O => \N__10643\,
            I => \N__10640\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__10640\,
            I => \N__10637\
        );

    \I__1508\ : Odrv4
    port map (
            O => \N__10637\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\
        );

    \I__1507\ : InMux
    port map (
            O => \N__10634\,
            I => \N__10631\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__10631\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\
        );

    \I__1505\ : InMux
    port map (
            O => \N__10628\,
            I => \N__10625\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__10625\,
            I => \N__10622\
        );

    \I__1503\ : Odrv4
    port map (
            O => \N__10622\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\
        );

    \I__1502\ : InMux
    port map (
            O => \N__10619\,
            I => \N__10615\
        );

    \I__1501\ : InMux
    port map (
            O => \N__10618\,
            I => \N__10612\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__10615\,
            I => \N__10609\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__10612\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__1498\ : Odrv4
    port map (
            O => \N__10609\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__1497\ : CascadeMux
    port map (
            O => \N__10604\,
            I => \N__10601\
        );

    \I__1496\ : InMux
    port map (
            O => \N__10601\,
            I => \N__10598\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__10598\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_13\
        );

    \I__1494\ : InMux
    port map (
            O => \N__10595\,
            I => \N__10591\
        );

    \I__1493\ : InMux
    port map (
            O => \N__10594\,
            I => \N__10588\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__10591\,
            I => \N__10585\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__10588\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__1490\ : Odrv4
    port map (
            O => \N__10585\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__1489\ : CascadeMux
    port map (
            O => \N__10580\,
            I => \N__10577\
        );

    \I__1488\ : InMux
    port map (
            O => \N__10577\,
            I => \N__10574\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__10574\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_14\
        );

    \I__1486\ : InMux
    port map (
            O => \N__10571\,
            I => \N__10567\
        );

    \I__1485\ : InMux
    port map (
            O => \N__10570\,
            I => \N__10564\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__10567\,
            I => \N__10561\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__10564\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__1482\ : Odrv12
    port map (
            O => \N__10561\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__1481\ : CascadeMux
    port map (
            O => \N__10556\,
            I => \N__10553\
        );

    \I__1480\ : InMux
    port map (
            O => \N__10553\,
            I => \N__10550\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__10550\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_15\
        );

    \I__1478\ : InMux
    port map (
            O => \N__10547\,
            I => \N__10543\
        );

    \I__1477\ : InMux
    port map (
            O => \N__10546\,
            I => \N__10540\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__10543\,
            I => \N__10537\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__10540\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__1474\ : Odrv12
    port map (
            O => \N__10537\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__1473\ : CascadeMux
    port map (
            O => \N__10532\,
            I => \N__10529\
        );

    \I__1472\ : InMux
    port map (
            O => \N__10529\,
            I => \N__10526\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__10526\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_16\
        );

    \I__1470\ : InMux
    port map (
            O => \N__10523\,
            I => \N__10519\
        );

    \I__1469\ : InMux
    port map (
            O => \N__10522\,
            I => \N__10516\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__10519\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__10516\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__1466\ : CascadeMux
    port map (
            O => \N__10511\,
            I => \N__10508\
        );

    \I__1465\ : InMux
    port map (
            O => \N__10508\,
            I => \N__10505\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__10505\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_17\
        );

    \I__1463\ : InMux
    port map (
            O => \N__10502\,
            I => \N__10498\
        );

    \I__1462\ : InMux
    port map (
            O => \N__10501\,
            I => \N__10495\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__10498\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__10495\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__1459\ : CascadeMux
    port map (
            O => \N__10490\,
            I => \N__10487\
        );

    \I__1458\ : InMux
    port map (
            O => \N__10487\,
            I => \N__10484\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__10484\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_18\
        );

    \I__1456\ : InMux
    port map (
            O => \N__10481\,
            I => \N__10477\
        );

    \I__1455\ : InMux
    port map (
            O => \N__10480\,
            I => \N__10474\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__10477\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__10474\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__1452\ : CascadeMux
    port map (
            O => \N__10469\,
            I => \N__10466\
        );

    \I__1451\ : InMux
    port map (
            O => \N__10466\,
            I => \N__10463\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__10463\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_19\
        );

    \I__1449\ : InMux
    port map (
            O => \N__10460\,
            I => \N__10456\
        );

    \I__1448\ : InMux
    port map (
            O => \N__10459\,
            I => \N__10453\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__10456\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__10453\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__1445\ : CascadeMux
    port map (
            O => \N__10448\,
            I => \N__10445\
        );

    \I__1444\ : InMux
    port map (
            O => \N__10445\,
            I => \N__10442\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__10442\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_5\
        );

    \I__1442\ : InMux
    port map (
            O => \N__10439\,
            I => \N__10435\
        );

    \I__1441\ : InMux
    port map (
            O => \N__10438\,
            I => \N__10432\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__10435\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__10432\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__1438\ : CascadeMux
    port map (
            O => \N__10427\,
            I => \N__10424\
        );

    \I__1437\ : InMux
    port map (
            O => \N__10424\,
            I => \N__10421\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__10421\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_6\
        );

    \I__1435\ : InMux
    port map (
            O => \N__10418\,
            I => \N__10414\
        );

    \I__1434\ : InMux
    port map (
            O => \N__10417\,
            I => \N__10411\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__10414\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__10411\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__1431\ : CascadeMux
    port map (
            O => \N__10406\,
            I => \N__10403\
        );

    \I__1430\ : InMux
    port map (
            O => \N__10403\,
            I => \N__10400\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__10400\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_7\
        );

    \I__1428\ : InMux
    port map (
            O => \N__10397\,
            I => \N__10393\
        );

    \I__1427\ : InMux
    port map (
            O => \N__10396\,
            I => \N__10390\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__10393\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__10390\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__1424\ : CascadeMux
    port map (
            O => \N__10385\,
            I => \N__10382\
        );

    \I__1423\ : InMux
    port map (
            O => \N__10382\,
            I => \N__10379\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__10379\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_8\
        );

    \I__1421\ : InMux
    port map (
            O => \N__10376\,
            I => \N__10373\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__10373\,
            I => \N__10369\
        );

    \I__1419\ : InMux
    port map (
            O => \N__10372\,
            I => \N__10366\
        );

    \I__1418\ : Odrv4
    port map (
            O => \N__10369\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__10366\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__1416\ : CascadeMux
    port map (
            O => \N__10361\,
            I => \N__10358\
        );

    \I__1415\ : InMux
    port map (
            O => \N__10358\,
            I => \N__10355\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__10355\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_9\
        );

    \I__1413\ : InMux
    port map (
            O => \N__10352\,
            I => \N__10349\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__10349\,
            I => \N__10345\
        );

    \I__1411\ : InMux
    port map (
            O => \N__10348\,
            I => \N__10342\
        );

    \I__1410\ : Odrv4
    port map (
            O => \N__10345\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__10342\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__1408\ : CascadeMux
    port map (
            O => \N__10337\,
            I => \N__10334\
        );

    \I__1407\ : InMux
    port map (
            O => \N__10334\,
            I => \N__10331\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__10331\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_10\
        );

    \I__1405\ : InMux
    port map (
            O => \N__10328\,
            I => \N__10325\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__10325\,
            I => \N__10321\
        );

    \I__1403\ : InMux
    port map (
            O => \N__10324\,
            I => \N__10318\
        );

    \I__1402\ : Odrv4
    port map (
            O => \N__10321\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__10318\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__1400\ : CascadeMux
    port map (
            O => \N__10313\,
            I => \N__10310\
        );

    \I__1399\ : InMux
    port map (
            O => \N__10310\,
            I => \N__10307\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__10307\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_11\
        );

    \I__1397\ : InMux
    port map (
            O => \N__10304\,
            I => \N__10300\
        );

    \I__1396\ : InMux
    port map (
            O => \N__10303\,
            I => \N__10297\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__10300\,
            I => \N__10294\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__10297\,
            I => \N__10291\
        );

    \I__1393\ : Odrv4
    port map (
            O => \N__10294\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__1392\ : Odrv4
    port map (
            O => \N__10291\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__1391\ : CascadeMux
    port map (
            O => \N__10286\,
            I => \N__10283\
        );

    \I__1390\ : InMux
    port map (
            O => \N__10283\,
            I => \N__10280\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__10280\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_12\
        );

    \I__1388\ : InMux
    port map (
            O => \N__10277\,
            I => \N__10274\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__10274\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13\
        );

    \I__1386\ : CascadeMux
    port map (
            O => \N__10271\,
            I => \N__10268\
        );

    \I__1385\ : InMux
    port map (
            O => \N__10268\,
            I => \N__10265\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__10265\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8\
        );

    \I__1383\ : InMux
    port map (
            O => \N__10262\,
            I => \N__10259\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__10259\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5\
        );

    \I__1381\ : CascadeMux
    port map (
            O => \N__10256\,
            I => \N__10253\
        );

    \I__1380\ : InMux
    port map (
            O => \N__10253\,
            I => \N__10250\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__10250\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4\
        );

    \I__1378\ : InMux
    port map (
            O => \N__10247\,
            I => \N__10244\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__10244\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2\
        );

    \I__1376\ : InMux
    port map (
            O => \N__10241\,
            I => \N__10237\
        );

    \I__1375\ : InMux
    port map (
            O => \N__10240\,
            I => \N__10233\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__10237\,
            I => \N__10230\
        );

    \I__1373\ : InMux
    port map (
            O => \N__10236\,
            I => \N__10227\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__10233\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__1371\ : Odrv4
    port map (
            O => \N__10230\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__10227\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__1369\ : CascadeMux
    port map (
            O => \N__10220\,
            I => \N__10217\
        );

    \I__1368\ : InMux
    port map (
            O => \N__10217\,
            I => \N__10214\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__10214\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_1\
        );

    \I__1366\ : InMux
    port map (
            O => \N__10211\,
            I => \N__10207\
        );

    \I__1365\ : InMux
    port map (
            O => \N__10210\,
            I => \N__10204\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__10207\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__10204\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__1362\ : InMux
    port map (
            O => \N__10199\,
            I => \N__10196\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__10196\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_2\
        );

    \I__1360\ : InMux
    port map (
            O => \N__10193\,
            I => \N__10189\
        );

    \I__1359\ : InMux
    port map (
            O => \N__10192\,
            I => \N__10186\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__10189\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__10186\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__1356\ : CascadeMux
    port map (
            O => \N__10181\,
            I => \N__10178\
        );

    \I__1355\ : InMux
    port map (
            O => \N__10178\,
            I => \N__10175\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__10175\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_3\
        );

    \I__1353\ : InMux
    port map (
            O => \N__10172\,
            I => \N__10168\
        );

    \I__1352\ : InMux
    port map (
            O => \N__10171\,
            I => \N__10165\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__10168\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__10165\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__1349\ : CascadeMux
    port map (
            O => \N__10160\,
            I => \N__10157\
        );

    \I__1348\ : InMux
    port map (
            O => \N__10157\,
            I => \N__10154\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__10154\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_4\
        );

    \I__1346\ : InMux
    port map (
            O => \N__10151\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__1345\ : CascadeMux
    port map (
            O => \N__10148\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO_cascade_\
        );

    \I__1344\ : CascadeMux
    port map (
            O => \N__10145\,
            I => \N__10142\
        );

    \I__1343\ : InMux
    port map (
            O => \N__10142\,
            I => \N__10139\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__10139\,
            I => \N__10136\
        );

    \I__1341\ : Span4Mux_s3_h
    port map (
            O => \N__10136\,
            I => \N__10133\
        );

    \I__1340\ : Odrv4
    port map (
            O => \N__10133\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\
        );

    \I__1339\ : InMux
    port map (
            O => \N__10130\,
            I => \N__10126\
        );

    \I__1338\ : InMux
    port map (
            O => \N__10129\,
            I => \N__10122\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__10126\,
            I => \N__10119\
        );

    \I__1336\ : InMux
    port map (
            O => \N__10125\,
            I => \N__10116\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__10122\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__1334\ : Odrv4
    port map (
            O => \N__10119\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__10116\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__1332\ : InMux
    port map (
            O => \N__10109\,
            I => \N__10106\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__10106\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0\
        );

    \I__1330\ : InMux
    port map (
            O => \N__10103\,
            I => \N__10100\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__10100\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16\
        );

    \I__1328\ : CascadeMux
    port map (
            O => \N__10097\,
            I => \N__10094\
        );

    \I__1327\ : InMux
    port map (
            O => \N__10094\,
            I => \N__10091\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__10091\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15\
        );

    \I__1325\ : InMux
    port map (
            O => \N__10088\,
            I => \N__10085\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__10085\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14\
        );

    \I__1323\ : CascadeMux
    port map (
            O => \N__10082\,
            I => \N__10079\
        );

    \I__1322\ : InMux
    port map (
            O => \N__10079\,
            I => \N__10076\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__10076\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6\
        );

    \I__1320\ : InMux
    port map (
            O => \N__10073\,
            I => \N__10070\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__10070\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7\
        );

    \I__1318\ : CascadeMux
    port map (
            O => \N__10067\,
            I => \N__10064\
        );

    \I__1317\ : InMux
    port map (
            O => \N__10064\,
            I => \N__10061\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__10061\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3\
        );

    \I__1315\ : InMux
    port map (
            O => \N__10058\,
            I => \N__10054\
        );

    \I__1314\ : InMux
    port map (
            O => \N__10057\,
            I => \N__10051\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__10054\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__10051\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__1311\ : CascadeMux
    port map (
            O => \N__10046\,
            I => \N__10043\
        );

    \I__1310\ : InMux
    port map (
            O => \N__10043\,
            I => \N__10040\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__10040\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\
        );

    \I__1308\ : InMux
    port map (
            O => \N__10037\,
            I => \N__10033\
        );

    \I__1307\ : InMux
    port map (
            O => \N__10036\,
            I => \N__10030\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__10033\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__10030\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__1304\ : CascadeMux
    port map (
            O => \N__10025\,
            I => \N__10022\
        );

    \I__1303\ : InMux
    port map (
            O => \N__10022\,
            I => \N__10019\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__10019\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\
        );

    \I__1301\ : InMux
    port map (
            O => \N__10016\,
            I => \N__10012\
        );

    \I__1300\ : InMux
    port map (
            O => \N__10015\,
            I => \N__10009\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__10012\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__10009\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__1297\ : CascadeMux
    port map (
            O => \N__10004\,
            I => \N__10001\
        );

    \I__1296\ : InMux
    port map (
            O => \N__10001\,
            I => \N__9998\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__9998\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\
        );

    \I__1294\ : InMux
    port map (
            O => \N__9995\,
            I => \N__9991\
        );

    \I__1293\ : InMux
    port map (
            O => \N__9994\,
            I => \N__9988\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__9991\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__9988\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__1290\ : CascadeMux
    port map (
            O => \N__9983\,
            I => \N__9980\
        );

    \I__1289\ : InMux
    port map (
            O => \N__9980\,
            I => \N__9977\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__9977\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_16\
        );

    \I__1287\ : InMux
    port map (
            O => \N__9974\,
            I => \N__9971\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__9971\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\
        );

    \I__1285\ : InMux
    port map (
            O => \N__9968\,
            I => \N__9964\
        );

    \I__1284\ : InMux
    port map (
            O => \N__9967\,
            I => \N__9961\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__9964\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__9961\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__1281\ : CascadeMux
    port map (
            O => \N__9956\,
            I => \N__9953\
        );

    \I__1280\ : InMux
    port map (
            O => \N__9953\,
            I => \N__9950\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__9950\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_17\
        );

    \I__1278\ : InMux
    port map (
            O => \N__9947\,
            I => \N__9944\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__9944\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\
        );

    \I__1276\ : InMux
    port map (
            O => \N__9941\,
            I => \N__9937\
        );

    \I__1275\ : InMux
    port map (
            O => \N__9940\,
            I => \N__9934\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__9937\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__9934\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__1272\ : CascadeMux
    port map (
            O => \N__9929\,
            I => \N__9926\
        );

    \I__1271\ : InMux
    port map (
            O => \N__9926\,
            I => \N__9923\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__9923\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_18\
        );

    \I__1269\ : InMux
    port map (
            O => \N__9920\,
            I => \N__9917\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__9917\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\
        );

    \I__1267\ : InMux
    port map (
            O => \N__9914\,
            I => \N__9910\
        );

    \I__1266\ : InMux
    port map (
            O => \N__9913\,
            I => \N__9907\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__9910\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__9907\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__1263\ : CascadeMux
    port map (
            O => \N__9902\,
            I => \N__9899\
        );

    \I__1262\ : InMux
    port map (
            O => \N__9899\,
            I => \N__9896\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__9896\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_19\
        );

    \I__1260\ : InMux
    port map (
            O => \N__9893\,
            I => \N__9889\
        );

    \I__1259\ : InMux
    port map (
            O => \N__9892\,
            I => \N__9886\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__9889\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__9886\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__1256\ : CascadeMux
    port map (
            O => \N__9881\,
            I => \N__9878\
        );

    \I__1255\ : InMux
    port map (
            O => \N__9878\,
            I => \N__9875\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__9875\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\
        );

    \I__1253\ : InMux
    port map (
            O => \N__9872\,
            I => \N__9868\
        );

    \I__1252\ : InMux
    port map (
            O => \N__9871\,
            I => \N__9865\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__9868\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__9865\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__1249\ : CascadeMux
    port map (
            O => \N__9860\,
            I => \N__9857\
        );

    \I__1248\ : InMux
    port map (
            O => \N__9857\,
            I => \N__9854\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__9854\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\
        );

    \I__1246\ : InMux
    port map (
            O => \N__9851\,
            I => \N__9847\
        );

    \I__1245\ : InMux
    port map (
            O => \N__9850\,
            I => \N__9844\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__9847\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__9844\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__1242\ : CascadeMux
    port map (
            O => \N__9839\,
            I => \N__9836\
        );

    \I__1241\ : InMux
    port map (
            O => \N__9836\,
            I => \N__9833\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__9833\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\
        );

    \I__1239\ : InMux
    port map (
            O => \N__9830\,
            I => \N__9826\
        );

    \I__1238\ : InMux
    port map (
            O => \N__9829\,
            I => \N__9823\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__9826\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__9823\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__1235\ : CascadeMux
    port map (
            O => \N__9818\,
            I => \N__9815\
        );

    \I__1234\ : InMux
    port map (
            O => \N__9815\,
            I => \N__9812\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__9812\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\
        );

    \I__1232\ : InMux
    port map (
            O => \N__9809\,
            I => \N__9805\
        );

    \I__1231\ : InMux
    port map (
            O => \N__9808\,
            I => \N__9802\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__9805\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__9802\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__1228\ : CascadeMux
    port map (
            O => \N__9797\,
            I => \N__9794\
        );

    \I__1227\ : InMux
    port map (
            O => \N__9794\,
            I => \N__9791\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__9791\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\
        );

    \I__1225\ : InMux
    port map (
            O => \N__9788\,
            I => \N__9784\
        );

    \I__1224\ : InMux
    port map (
            O => \N__9787\,
            I => \N__9781\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__9784\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__9781\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__1221\ : CascadeMux
    port map (
            O => \N__9776\,
            I => \N__9773\
        );

    \I__1220\ : InMux
    port map (
            O => \N__9773\,
            I => \N__9770\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__9770\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\
        );

    \I__1218\ : InMux
    port map (
            O => \N__9767\,
            I => \N__9763\
        );

    \I__1217\ : InMux
    port map (
            O => \N__9766\,
            I => \N__9760\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__9763\,
            I => \N__9757\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__9760\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__1214\ : Odrv4
    port map (
            O => \N__9757\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__1213\ : CascadeMux
    port map (
            O => \N__9752\,
            I => \N__9749\
        );

    \I__1212\ : InMux
    port map (
            O => \N__9749\,
            I => \N__9746\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__9746\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\
        );

    \I__1210\ : InMux
    port map (
            O => \N__9743\,
            I => \N__9739\
        );

    \I__1209\ : InMux
    port map (
            O => \N__9742\,
            I => \N__9736\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__9739\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__9736\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__1206\ : CascadeMux
    port map (
            O => \N__9731\,
            I => \N__9728\
        );

    \I__1205\ : InMux
    port map (
            O => \N__9728\,
            I => \N__9725\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__9725\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\
        );

    \I__1203\ : CascadeMux
    port map (
            O => \N__9722\,
            I => \N__9717\
        );

    \I__1202\ : CascadeMux
    port map (
            O => \N__9721\,
            I => \N__9714\
        );

    \I__1201\ : CascadeMux
    port map (
            O => \N__9720\,
            I => \N__9711\
        );

    \I__1200\ : InMux
    port map (
            O => \N__9717\,
            I => \N__9688\
        );

    \I__1199\ : InMux
    port map (
            O => \N__9714\,
            I => \N__9688\
        );

    \I__1198\ : InMux
    port map (
            O => \N__9711\,
            I => \N__9688\
        );

    \I__1197\ : InMux
    port map (
            O => \N__9710\,
            I => \N__9679\
        );

    \I__1196\ : InMux
    port map (
            O => \N__9709\,
            I => \N__9679\
        );

    \I__1195\ : InMux
    port map (
            O => \N__9708\,
            I => \N__9679\
        );

    \I__1194\ : InMux
    port map (
            O => \N__9707\,
            I => \N__9679\
        );

    \I__1193\ : InMux
    port map (
            O => \N__9706\,
            I => \N__9668\
        );

    \I__1192\ : InMux
    port map (
            O => \N__9705\,
            I => \N__9668\
        );

    \I__1191\ : InMux
    port map (
            O => \N__9704\,
            I => \N__9668\
        );

    \I__1190\ : InMux
    port map (
            O => \N__9703\,
            I => \N__9668\
        );

    \I__1189\ : InMux
    port map (
            O => \N__9702\,
            I => \N__9651\
        );

    \I__1188\ : InMux
    port map (
            O => \N__9701\,
            I => \N__9651\
        );

    \I__1187\ : InMux
    port map (
            O => \N__9700\,
            I => \N__9651\
        );

    \I__1186\ : InMux
    port map (
            O => \N__9699\,
            I => \N__9651\
        );

    \I__1185\ : InMux
    port map (
            O => \N__9698\,
            I => \N__9651\
        );

    \I__1184\ : InMux
    port map (
            O => \N__9697\,
            I => \N__9651\
        );

    \I__1183\ : InMux
    port map (
            O => \N__9696\,
            I => \N__9651\
        );

    \I__1182\ : InMux
    port map (
            O => \N__9695\,
            I => \N__9651\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__9688\,
            I => \N__9646\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__9679\,
            I => \N__9646\
        );

    \I__1179\ : InMux
    port map (
            O => \N__9678\,
            I => \N__9638\
        );

    \I__1178\ : InMux
    port map (
            O => \N__9677\,
            I => \N__9638\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__9668\,
            I => \N__9631\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__9651\,
            I => \N__9631\
        );

    \I__1175\ : Span4Mux_s3_h
    port map (
            O => \N__9646\,
            I => \N__9631\
        );

    \I__1174\ : InMux
    port map (
            O => \N__9645\,
            I => \N__9626\
        );

    \I__1173\ : InMux
    port map (
            O => \N__9644\,
            I => \N__9626\
        );

    \I__1172\ : InMux
    port map (
            O => \N__9643\,
            I => \N__9623\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__9638\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__1170\ : Odrv4
    port map (
            O => \N__9631\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__9626\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__9623\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__1167\ : CascadeMux
    port map (
            O => \N__9614\,
            I => \N__9595\
        );

    \I__1166\ : InMux
    port map (
            O => \N__9613\,
            I => \N__9575\
        );

    \I__1165\ : InMux
    port map (
            O => \N__9612\,
            I => \N__9575\
        );

    \I__1164\ : InMux
    port map (
            O => \N__9611\,
            I => \N__9575\
        );

    \I__1163\ : InMux
    port map (
            O => \N__9610\,
            I => \N__9575\
        );

    \I__1162\ : InMux
    port map (
            O => \N__9609\,
            I => \N__9575\
        );

    \I__1161\ : InMux
    port map (
            O => \N__9608\,
            I => \N__9575\
        );

    \I__1160\ : InMux
    port map (
            O => \N__9607\,
            I => \N__9575\
        );

    \I__1159\ : InMux
    port map (
            O => \N__9606\,
            I => \N__9575\
        );

    \I__1158\ : InMux
    port map (
            O => \N__9605\,
            I => \N__9560\
        );

    \I__1157\ : InMux
    port map (
            O => \N__9604\,
            I => \N__9560\
        );

    \I__1156\ : InMux
    port map (
            O => \N__9603\,
            I => \N__9560\
        );

    \I__1155\ : InMux
    port map (
            O => \N__9602\,
            I => \N__9560\
        );

    \I__1154\ : InMux
    port map (
            O => \N__9601\,
            I => \N__9560\
        );

    \I__1153\ : InMux
    port map (
            O => \N__9600\,
            I => \N__9560\
        );

    \I__1152\ : InMux
    port map (
            O => \N__9599\,
            I => \N__9560\
        );

    \I__1151\ : CascadeMux
    port map (
            O => \N__9598\,
            I => \N__9557\
        );

    \I__1150\ : InMux
    port map (
            O => \N__9595\,
            I => \N__9547\
        );

    \I__1149\ : InMux
    port map (
            O => \N__9594\,
            I => \N__9547\
        );

    \I__1148\ : InMux
    port map (
            O => \N__9593\,
            I => \N__9547\
        );

    \I__1147\ : InMux
    port map (
            O => \N__9592\,
            I => \N__9547\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__9575\,
            I => \N__9542\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__9560\,
            I => \N__9542\
        );

    \I__1144\ : InMux
    port map (
            O => \N__9557\,
            I => \N__9534\
        );

    \I__1143\ : InMux
    port map (
            O => \N__9556\,
            I => \N__9534\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__9547\,
            I => \N__9531\
        );

    \I__1141\ : Span4Mux_v
    port map (
            O => \N__9542\,
            I => \N__9528\
        );

    \I__1140\ : InMux
    port map (
            O => \N__9541\,
            I => \N__9523\
        );

    \I__1139\ : InMux
    port map (
            O => \N__9540\,
            I => \N__9523\
        );

    \I__1138\ : InMux
    port map (
            O => \N__9539\,
            I => \N__9520\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__9534\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__1136\ : Odrv4
    port map (
            O => \N__9531\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__1135\ : Odrv4
    port map (
            O => \N__9528\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__9523\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__9520\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__1132\ : InMux
    port map (
            O => \N__9509\,
            I => \N__9494\
        );

    \I__1131\ : InMux
    port map (
            O => \N__9508\,
            I => \N__9494\
        );

    \I__1130\ : InMux
    port map (
            O => \N__9507\,
            I => \N__9494\
        );

    \I__1129\ : InMux
    port map (
            O => \N__9506\,
            I => \N__9494\
        );

    \I__1128\ : InMux
    port map (
            O => \N__9505\,
            I => \N__9476\
        );

    \I__1127\ : InMux
    port map (
            O => \N__9504\,
            I => \N__9469\
        );

    \I__1126\ : InMux
    port map (
            O => \N__9503\,
            I => \N__9469\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__9494\,
            I => \N__9466\
        );

    \I__1124\ : InMux
    port map (
            O => \N__9493\,
            I => \N__9449\
        );

    \I__1123\ : InMux
    port map (
            O => \N__9492\,
            I => \N__9449\
        );

    \I__1122\ : InMux
    port map (
            O => \N__9491\,
            I => \N__9449\
        );

    \I__1121\ : InMux
    port map (
            O => \N__9490\,
            I => \N__9449\
        );

    \I__1120\ : InMux
    port map (
            O => \N__9489\,
            I => \N__9449\
        );

    \I__1119\ : InMux
    port map (
            O => \N__9488\,
            I => \N__9449\
        );

    \I__1118\ : InMux
    port map (
            O => \N__9487\,
            I => \N__9449\
        );

    \I__1117\ : InMux
    port map (
            O => \N__9486\,
            I => \N__9449\
        );

    \I__1116\ : InMux
    port map (
            O => \N__9485\,
            I => \N__9434\
        );

    \I__1115\ : InMux
    port map (
            O => \N__9484\,
            I => \N__9434\
        );

    \I__1114\ : InMux
    port map (
            O => \N__9483\,
            I => \N__9434\
        );

    \I__1113\ : InMux
    port map (
            O => \N__9482\,
            I => \N__9434\
        );

    \I__1112\ : InMux
    port map (
            O => \N__9481\,
            I => \N__9434\
        );

    \I__1111\ : InMux
    port map (
            O => \N__9480\,
            I => \N__9434\
        );

    \I__1110\ : InMux
    port map (
            O => \N__9479\,
            I => \N__9434\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__9476\,
            I => \N__9431\
        );

    \I__1108\ : InMux
    port map (
            O => \N__9475\,
            I => \N__9426\
        );

    \I__1107\ : InMux
    port map (
            O => \N__9474\,
            I => \N__9426\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__9469\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__1105\ : Odrv4
    port map (
            O => \N__9466\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__9449\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__9434\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__1102\ : Odrv4
    port map (
            O => \N__9431\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__9426\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__1100\ : CascadeMux
    port map (
            O => \N__9413\,
            I => \N__9403\
        );

    \I__1099\ : CascadeMux
    port map (
            O => \N__9412\,
            I => \N__9400\
        );

    \I__1098\ : CascadeMux
    port map (
            O => \N__9411\,
            I => \N__9397\
        );

    \I__1097\ : CascadeMux
    port map (
            O => \N__9410\,
            I => \N__9394\
        );

    \I__1096\ : CascadeMux
    port map (
            O => \N__9409\,
            I => \N__9387\
        );

    \I__1095\ : CascadeMux
    port map (
            O => \N__9408\,
            I => \N__9384\
        );

    \I__1094\ : CascadeMux
    port map (
            O => \N__9407\,
            I => \N__9381\
        );

    \I__1093\ : CascadeMux
    port map (
            O => \N__9406\,
            I => \N__9378\
        );

    \I__1092\ : InMux
    port map (
            O => \N__9403\,
            I => \N__9360\
        );

    \I__1091\ : InMux
    port map (
            O => \N__9400\,
            I => \N__9360\
        );

    \I__1090\ : InMux
    port map (
            O => \N__9397\,
            I => \N__9360\
        );

    \I__1089\ : InMux
    port map (
            O => \N__9394\,
            I => \N__9360\
        );

    \I__1088\ : InMux
    port map (
            O => \N__9393\,
            I => \N__9351\
        );

    \I__1087\ : InMux
    port map (
            O => \N__9392\,
            I => \N__9351\
        );

    \I__1086\ : InMux
    port map (
            O => \N__9391\,
            I => \N__9351\
        );

    \I__1085\ : InMux
    port map (
            O => \N__9390\,
            I => \N__9351\
        );

    \I__1084\ : InMux
    port map (
            O => \N__9387\,
            I => \N__9339\
        );

    \I__1083\ : InMux
    port map (
            O => \N__9384\,
            I => \N__9339\
        );

    \I__1082\ : InMux
    port map (
            O => \N__9381\,
            I => \N__9339\
        );

    \I__1081\ : InMux
    port map (
            O => \N__9378\,
            I => \N__9339\
        );

    \I__1080\ : InMux
    port map (
            O => \N__9377\,
            I => \N__9334\
        );

    \I__1079\ : InMux
    port map (
            O => \N__9376\,
            I => \N__9334\
        );

    \I__1078\ : InMux
    port map (
            O => \N__9375\,
            I => \N__9325\
        );

    \I__1077\ : InMux
    port map (
            O => \N__9374\,
            I => \N__9325\
        );

    \I__1076\ : InMux
    port map (
            O => \N__9373\,
            I => \N__9325\
        );

    \I__1075\ : InMux
    port map (
            O => \N__9372\,
            I => \N__9325\
        );

    \I__1074\ : InMux
    port map (
            O => \N__9371\,
            I => \N__9318\
        );

    \I__1073\ : InMux
    port map (
            O => \N__9370\,
            I => \N__9318\
        );

    \I__1072\ : InMux
    port map (
            O => \N__9369\,
            I => \N__9318\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__9360\,
            I => \N__9313\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__9351\,
            I => \N__9313\
        );

    \I__1069\ : InMux
    port map (
            O => \N__9350\,
            I => \N__9310\
        );

    \I__1068\ : InMux
    port map (
            O => \N__9349\,
            I => \N__9305\
        );

    \I__1067\ : InMux
    port map (
            O => \N__9348\,
            I => \N__9305\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__9339\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__9334\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__9325\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__9318\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__1062\ : Odrv4
    port map (
            O => \N__9313\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__9310\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__9305\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__1059\ : CascadeMux
    port map (
            O => \N__9290\,
            I => \N__9287\
        );

    \I__1058\ : InMux
    port map (
            O => \N__9287\,
            I => \N__9284\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__9284\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\
        );

    \I__1056\ : CascadeMux
    port map (
            O => \N__9281\,
            I => \N__9278\
        );

    \I__1055\ : InMux
    port map (
            O => \N__9278\,
            I => \N__9274\
        );

    \I__1054\ : InMux
    port map (
            O => \N__9277\,
            I => \N__9271\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__9274\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__9271\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__1051\ : CascadeMux
    port map (
            O => \N__9266\,
            I => \N__9263\
        );

    \I__1050\ : InMux
    port map (
            O => \N__9263\,
            I => \N__9260\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__9260\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\
        );

    \I__1048\ : InMux
    port map (
            O => \N__9257\,
            I => \N__9254\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__9254\,
            I => \N__9250\
        );

    \I__1046\ : InMux
    port map (
            O => \N__9253\,
            I => \N__9247\
        );

    \I__1045\ : Odrv4
    port map (
            O => \N__9250\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__9247\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__1043\ : CascadeMux
    port map (
            O => \N__9242\,
            I => \N__9239\
        );

    \I__1042\ : InMux
    port map (
            O => \N__9239\,
            I => \N__9236\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__9236\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\
        );

    \I__1040\ : InMux
    port map (
            O => \N__9233\,
            I => \N__9229\
        );

    \I__1039\ : InMux
    port map (
            O => \N__9232\,
            I => \N__9226\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__9229\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__9226\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__1036\ : CascadeMux
    port map (
            O => \N__9221\,
            I => \N__9218\
        );

    \I__1035\ : InMux
    port map (
            O => \N__9218\,
            I => \N__9215\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__9215\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\
        );

    \I__1033\ : InMux
    port map (
            O => \N__9212\,
            I => \N__9208\
        );

    \I__1032\ : InMux
    port map (
            O => \N__9211\,
            I => \N__9205\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__9208\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__9205\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__1029\ : CascadeMux
    port map (
            O => \N__9200\,
            I => \N__9197\
        );

    \I__1028\ : InMux
    port map (
            O => \N__9197\,
            I => \N__9194\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__9194\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_16\
        );

    \I__1026\ : InMux
    port map (
            O => \N__9191\,
            I => \N__9187\
        );

    \I__1025\ : InMux
    port map (
            O => \N__9190\,
            I => \N__9184\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__9187\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__9184\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__1022\ : CascadeMux
    port map (
            O => \N__9179\,
            I => \N__9176\
        );

    \I__1021\ : InMux
    port map (
            O => \N__9176\,
            I => \N__9173\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__9173\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_17\
        );

    \I__1019\ : InMux
    port map (
            O => \N__9170\,
            I => \N__9167\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__9167\,
            I => \N__9164\
        );

    \I__1017\ : Span4Mux_v
    port map (
            O => \N__9164\,
            I => \N__9161\
        );

    \I__1016\ : Odrv4
    port map (
            O => \N__9161\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\
        );

    \I__1015\ : InMux
    port map (
            O => \N__9158\,
            I => \N__9154\
        );

    \I__1014\ : InMux
    port map (
            O => \N__9157\,
            I => \N__9151\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__9154\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__9151\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__1011\ : CascadeMux
    port map (
            O => \N__9146\,
            I => \N__9143\
        );

    \I__1010\ : InMux
    port map (
            O => \N__9143\,
            I => \N__9140\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__9140\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_18\
        );

    \I__1008\ : InMux
    port map (
            O => \N__9137\,
            I => \N__9133\
        );

    \I__1007\ : InMux
    port map (
            O => \N__9136\,
            I => \N__9130\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__9133\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__9130\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__1004\ : CascadeMux
    port map (
            O => \N__9125\,
            I => \N__9122\
        );

    \I__1003\ : InMux
    port map (
            O => \N__9122\,
            I => \N__9119\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__9119\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_19\
        );

    \I__1001\ : InMux
    port map (
            O => \N__9116\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__1000\ : CascadeMux
    port map (
            O => \N__9113\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_\
        );

    \I__999\ : CascadeMux
    port map (
            O => \N__9110\,
            I => \N__9107\
        );

    \I__998\ : InMux
    port map (
            O => \N__9107\,
            I => \N__9104\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__9104\,
            I => \N__9101\
        );

    \I__996\ : Span4Mux_v
    port map (
            O => \N__9101\,
            I => \N__9098\
        );

    \I__995\ : Odrv4
    port map (
            O => \N__9098\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\
        );

    \I__994\ : InMux
    port map (
            O => \N__9095\,
            I => \N__9092\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__9092\,
            I => \N__9089\
        );

    \I__992\ : Odrv4
    port map (
            O => \N__9089\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\
        );

    \I__991\ : CascadeMux
    port map (
            O => \N__9086\,
            I => \N__9083\
        );

    \I__990\ : InMux
    port map (
            O => \N__9083\,
            I => \N__9079\
        );

    \I__989\ : InMux
    port map (
            O => \N__9082\,
            I => \N__9076\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__9079\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__9076\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__986\ : CascadeMux
    port map (
            O => \N__9071\,
            I => \N__9068\
        );

    \I__985\ : InMux
    port map (
            O => \N__9068\,
            I => \N__9065\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__9065\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\
        );

    \I__983\ : InMux
    port map (
            O => \N__9062\,
            I => \N__9058\
        );

    \I__982\ : InMux
    port map (
            O => \N__9061\,
            I => \N__9055\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__9058\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__9055\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__979\ : CascadeMux
    port map (
            O => \N__9050\,
            I => \N__9047\
        );

    \I__978\ : InMux
    port map (
            O => \N__9047\,
            I => \N__9044\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__9044\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\
        );

    \I__976\ : InMux
    port map (
            O => \N__9041\,
            I => \N__9037\
        );

    \I__975\ : InMux
    port map (
            O => \N__9040\,
            I => \N__9034\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__9037\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__9034\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__972\ : CascadeMux
    port map (
            O => \N__9029\,
            I => \N__9026\
        );

    \I__971\ : InMux
    port map (
            O => \N__9026\,
            I => \N__9023\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__9023\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\
        );

    \I__969\ : InMux
    port map (
            O => \N__9020\,
            I => \N__9016\
        );

    \I__968\ : InMux
    port map (
            O => \N__9019\,
            I => \N__9013\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__9016\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__9013\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__965\ : CascadeMux
    port map (
            O => \N__9008\,
            I => \N__9005\
        );

    \I__964\ : InMux
    port map (
            O => \N__9005\,
            I => \N__9002\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__9002\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\
        );

    \I__962\ : InMux
    port map (
            O => \N__8999\,
            I => \N__8995\
        );

    \I__961\ : InMux
    port map (
            O => \N__8998\,
            I => \N__8992\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__8995\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__8992\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__958\ : CascadeMux
    port map (
            O => \N__8987\,
            I => \N__8984\
        );

    \I__957\ : InMux
    port map (
            O => \N__8984\,
            I => \N__8981\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__8981\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\
        );

    \I__955\ : InMux
    port map (
            O => \N__8978\,
            I => \N__8974\
        );

    \I__954\ : InMux
    port map (
            O => \N__8977\,
            I => \N__8971\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__8974\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__8971\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__951\ : CascadeMux
    port map (
            O => \N__8966\,
            I => \N__8963\
        );

    \I__950\ : InMux
    port map (
            O => \N__8963\,
            I => \N__8960\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__8960\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\
        );

    \I__948\ : InMux
    port map (
            O => \N__8957\,
            I => \N__8953\
        );

    \I__947\ : InMux
    port map (
            O => \N__8956\,
            I => \N__8950\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__8953\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__8950\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__944\ : CascadeMux
    port map (
            O => \N__8945\,
            I => \N__8942\
        );

    \I__943\ : InMux
    port map (
            O => \N__8942\,
            I => \N__8939\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__8939\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\
        );

    \I__941\ : InMux
    port map (
            O => \N__8936\,
            I => \N__8932\
        );

    \I__940\ : InMux
    port map (
            O => \N__8935\,
            I => \N__8929\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__8932\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__8929\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__937\ : CascadeMux
    port map (
            O => \N__8924\,
            I => \N__8921\
        );

    \I__936\ : InMux
    port map (
            O => \N__8921\,
            I => \N__8918\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__8918\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\
        );

    \I__934\ : InMux
    port map (
            O => \N__8915\,
            I => \N__8911\
        );

    \I__933\ : InMux
    port map (
            O => \N__8914\,
            I => \N__8907\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__8911\,
            I => \N__8904\
        );

    \I__931\ : InMux
    port map (
            O => \N__8910\,
            I => \N__8901\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__8907\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__929\ : Odrv4
    port map (
            O => \N__8904\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__8901\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__927\ : CascadeMux
    port map (
            O => \N__8894\,
            I => \N__8891\
        );

    \I__926\ : InMux
    port map (
            O => \N__8891\,
            I => \N__8888\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__8888\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\
        );

    \I__924\ : InMux
    port map (
            O => \N__8885\,
            I => \N__8881\
        );

    \I__923\ : InMux
    port map (
            O => \N__8884\,
            I => \N__8878\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__8881\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__8878\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__920\ : CascadeMux
    port map (
            O => \N__8873\,
            I => \N__8870\
        );

    \I__919\ : InMux
    port map (
            O => \N__8870\,
            I => \N__8867\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__8867\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\
        );

    \I__917\ : InMux
    port map (
            O => \N__8864\,
            I => \N__8860\
        );

    \I__916\ : InMux
    port map (
            O => \N__8863\,
            I => \N__8857\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__8860\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__8857\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__913\ : CascadeMux
    port map (
            O => \N__8852\,
            I => \N__8849\
        );

    \I__912\ : InMux
    port map (
            O => \N__8849\,
            I => \N__8846\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__8846\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\
        );

    \I__910\ : InMux
    port map (
            O => \N__8843\,
            I => \N__8839\
        );

    \I__909\ : InMux
    port map (
            O => \N__8842\,
            I => \N__8836\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__8839\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__8836\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__906\ : CascadeMux
    port map (
            O => \N__8831\,
            I => \N__8828\
        );

    \I__905\ : InMux
    port map (
            O => \N__8828\,
            I => \N__8825\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__8825\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\
        );

    \I__903\ : InMux
    port map (
            O => \N__8822\,
            I => \N__8818\
        );

    \I__902\ : InMux
    port map (
            O => \N__8821\,
            I => \N__8815\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__8818\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__8815\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__899\ : CascadeMux
    port map (
            O => \N__8810\,
            I => \N__8807\
        );

    \I__898\ : InMux
    port map (
            O => \N__8807\,
            I => \N__8804\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__8804\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\
        );

    \I__896\ : InMux
    port map (
            O => \N__8801\,
            I => \N__8797\
        );

    \I__895\ : InMux
    port map (
            O => \N__8800\,
            I => \N__8794\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__8797\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__8794\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__892\ : CascadeMux
    port map (
            O => \N__8789\,
            I => \N__8786\
        );

    \I__891\ : InMux
    port map (
            O => \N__8786\,
            I => \N__8783\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__8783\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\
        );

    \I__889\ : InMux
    port map (
            O => \N__8780\,
            I => \N__8776\
        );

    \I__888\ : InMux
    port map (
            O => \N__8779\,
            I => \N__8773\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__8776\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__8773\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__885\ : InMux
    port map (
            O => \N__8768\,
            I => \N__8765\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__8765\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\
        );

    \I__883\ : CascadeMux
    port map (
            O => \N__8762\,
            I => \N__8759\
        );

    \I__882\ : InMux
    port map (
            O => \N__8759\,
            I => \N__8756\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__8756\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\
        );

    \I__880\ : CascadeMux
    port map (
            O => \N__8753\,
            I => \N__8750\
        );

    \I__879\ : InMux
    port map (
            O => \N__8750\,
            I => \N__8747\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__8747\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18\
        );

    \I__877\ : InMux
    port map (
            O => \N__8744\,
            I => \N__8741\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__8741\,
            I => \N__8738\
        );

    \I__875\ : Odrv4
    port map (
            O => \N__8738\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11\
        );

    \I__874\ : CascadeMux
    port map (
            O => \N__8735\,
            I => \phase_controller_slave.stoper_hc.time_passed11_cascade_\
        );

    \I__873\ : CascadeMux
    port map (
            O => \N__8732\,
            I => \N__8729\
        );

    \I__872\ : InMux
    port map (
            O => \N__8729\,
            I => \N__8726\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__8726\,
            I => \N__8723\
        );

    \I__870\ : Span4Mux_h
    port map (
            O => \N__8723\,
            I => \N__8720\
        );

    \I__869\ : Odrv4
    port map (
            O => \N__8720\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0\
        );

    \I__868\ : InMux
    port map (
            O => \N__8717\,
            I => \N__8714\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__8714\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0\
        );

    \I__866\ : InMux
    port map (
            O => \N__8711\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14\
        );

    \I__865\ : InMux
    port map (
            O => \N__8708\,
            I => \bfn_2_25_0_\
        );

    \I__864\ : InMux
    port map (
            O => \N__8705\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16\
        );

    \I__863\ : InMux
    port map (
            O => \N__8702\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17\
        );

    \I__862\ : InMux
    port map (
            O => \N__8699\,
            I => \N__8696\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__8696\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17\
        );

    \I__860\ : InMux
    port map (
            O => \N__8693\,
            I => \N__8690\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__8690\,
            I => \N__8687\
        );

    \I__858\ : Odrv4
    port map (
            O => \N__8687\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12\
        );

    \I__857\ : InMux
    port map (
            O => \N__8684\,
            I => \N__8681\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__8681\,
            I => \N__8678\
        );

    \I__855\ : Odrv4
    port map (
            O => \N__8678\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9\
        );

    \I__854\ : InMux
    port map (
            O => \N__8675\,
            I => \N__8672\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__8672\,
            I => \N__8669\
        );

    \I__852\ : Odrv4
    port map (
            O => \N__8669\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10\
        );

    \I__851\ : InMux
    port map (
            O => \N__8666\,
            I => \N__8663\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__8663\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19\
        );

    \I__849\ : InMux
    port map (
            O => \N__8660\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5\
        );

    \I__848\ : InMux
    port map (
            O => \N__8657\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6\
        );

    \I__847\ : InMux
    port map (
            O => \N__8654\,
            I => \bfn_2_24_0_\
        );

    \I__846\ : InMux
    port map (
            O => \N__8651\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8\
        );

    \I__845\ : InMux
    port map (
            O => \N__8648\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9\
        );

    \I__844\ : InMux
    port map (
            O => \N__8645\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10\
        );

    \I__843\ : InMux
    port map (
            O => \N__8642\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11\
        );

    \I__842\ : InMux
    port map (
            O => \N__8639\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12\
        );

    \I__841\ : InMux
    port map (
            O => \N__8636\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13\
        );

    \I__840\ : InMux
    port map (
            O => \N__8633\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0\
        );

    \I__839\ : InMux
    port map (
            O => \N__8630\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1\
        );

    \I__838\ : InMux
    port map (
            O => \N__8627\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2\
        );

    \I__837\ : InMux
    port map (
            O => \N__8624\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3\
        );

    \I__836\ : InMux
    port map (
            O => \N__8621\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4\
        );

    \I__835\ : InMux
    port map (
            O => \N__8618\,
            I => \N__8615\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__8615\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\
        );

    \I__833\ : InMux
    port map (
            O => \N__8612\,
            I => \N__8609\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__8609\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\
        );

    \I__831\ : InMux
    port map (
            O => \N__8606\,
            I => \N__8603\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__8603\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\
        );

    \I__829\ : InMux
    port map (
            O => \N__8600\,
            I => \N__8597\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__8597\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\
        );

    \I__827\ : InMux
    port map (
            O => \N__8594\,
            I => \N__8591\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__8591\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\
        );

    \I__825\ : InMux
    port map (
            O => \N__8588\,
            I => \N__8585\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__8585\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\
        );

    \I__823\ : InMux
    port map (
            O => \N__8582\,
            I => \N__8579\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__8579\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\
        );

    \I__821\ : InMux
    port map (
            O => \N__8576\,
            I => \N__8573\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__8573\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\
        );

    \I__819\ : InMux
    port map (
            O => \N__8570\,
            I => \N__8567\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__8567\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\
        );

    \I__817\ : InMux
    port map (
            O => \N__8564\,
            I => \N__8561\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__8561\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\
        );

    \I__815\ : InMux
    port map (
            O => \N__8558\,
            I => \N__8555\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__8555\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\
        );

    \I__813\ : InMux
    port map (
            O => \N__8552\,
            I => \N__8549\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__8549\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\
        );

    \I__811\ : InMux
    port map (
            O => \N__8546\,
            I => \N__8543\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__8543\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\
        );

    \I__809\ : InMux
    port map (
            O => \N__8540\,
            I => \N__8537\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__8537\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\
        );

    \I__807\ : InMux
    port map (
            O => \N__8534\,
            I => \N__8531\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__8531\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\
        );

    \I__805\ : InMux
    port map (
            O => \N__8528\,
            I => \N__8525\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__8525\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\
        );

    \I__803\ : InMux
    port map (
            O => \N__8522\,
            I => \N__8519\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__8519\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\
        );

    \I__801\ : InMux
    port map (
            O => \N__8516\,
            I => \N__8513\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__8513\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\
        );

    \I__799\ : InMux
    port map (
            O => \N__8510\,
            I => \N__8507\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__8507\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\
        );

    \I__797\ : InMux
    port map (
            O => \N__8504\,
            I => \N__8501\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__8501\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\
        );

    \I__795\ : CascadeMux
    port map (
            O => \N__8498\,
            I => \N__8495\
        );

    \I__794\ : InMux
    port map (
            O => \N__8495\,
            I => \N__8492\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__8492\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\
        );

    \I__792\ : InMux
    port map (
            O => \N__8489\,
            I => \N__8486\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__8486\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0\
        );

    \I__790\ : CascadeMux
    port map (
            O => \N__8483\,
            I => \phase_controller_inst1.stoper_tr.time_passed11_cascade_\
        );

    \I__789\ : CascadeMux
    port map (
            O => \N__8480\,
            I => \N__8477\
        );

    \I__788\ : InMux
    port map (
            O => \N__8477\,
            I => \N__8474\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__8474\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0\
        );

    \I__786\ : CascadeMux
    port map (
            O => \N__8471\,
            I => \phase_controller_inst1.stoper_hc.time_passed11_cascade_\
        );

    \I__785\ : CascadeMux
    port map (
            O => \N__8468\,
            I => \N__8465\
        );

    \I__784\ : InMux
    port map (
            O => \N__8465\,
            I => \N__8462\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__8462\,
            I => \N__8459\
        );

    \I__782\ : Span4Mux_s2_h
    port map (
            O => \N__8459\,
            I => \N__8456\
        );

    \I__781\ : Odrv4
    port map (
            O => \N__8456\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0\
        );

    \I__780\ : InMux
    port map (
            O => \N__8453\,
            I => \N__8450\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__8450\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\
        );

    \I__778\ : CascadeMux
    port map (
            O => \N__8447\,
            I => \N__8444\
        );

    \I__777\ : InMux
    port map (
            O => \N__8444\,
            I => \N__8441\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__8441\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\
        );

    \I__775\ : InMux
    port map (
            O => \N__8438\,
            I => \N__8435\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__8435\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\
        );

    \I__773\ : CascadeMux
    port map (
            O => \N__8432\,
            I => \N__8429\
        );

    \I__772\ : InMux
    port map (
            O => \N__8429\,
            I => \N__8426\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__8426\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\
        );

    \I__770\ : InMux
    port map (
            O => \N__8423\,
            I => \N__8420\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__8420\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\
        );

    \I__768\ : CascadeMux
    port map (
            O => \N__8417\,
            I => \N__8414\
        );

    \I__767\ : InMux
    port map (
            O => \N__8414\,
            I => \N__8411\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__8411\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\
        );

    \I__765\ : InMux
    port map (
            O => \N__8408\,
            I => \N__8405\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__8405\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\
        );

    \I__763\ : CascadeMux
    port map (
            O => \N__8402\,
            I => \N__8399\
        );

    \I__762\ : InMux
    port map (
            O => \N__8399\,
            I => \N__8396\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__8396\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\
        );

    \I__760\ : InMux
    port map (
            O => \N__8393\,
            I => \N__8390\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__8390\,
            I => \rgb_drv_RNOZ0\
        );

    \I__758\ : InMux
    port map (
            O => \N__8387\,
            I => \N__8384\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__8384\,
            I => \N_39_i_i\
        );

    \I__756\ : InMux
    port map (
            O => \N__8381\,
            I => \N__8378\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__8378\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\
        );

    \I__754\ : InMux
    port map (
            O => \N__8375\,
            I => \N__8372\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__8372\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\
        );

    \I__752\ : InMux
    port map (
            O => \N__8369\,
            I => \N__8366\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__8366\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\
        );

    \I__750\ : InMux
    port map (
            O => \N__8363\,
            I => \N__8360\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__8360\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\
        );

    \I__748\ : InMux
    port map (
            O => \N__8357\,
            I => \N__8354\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__8354\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\
        );

    \I__746\ : InMux
    port map (
            O => \N__8351\,
            I => \N__8348\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__8348\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\
        );

    \I__744\ : InMux
    port map (
            O => \N__8345\,
            I => \N__8342\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__8342\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\
        );

    \I__742\ : InMux
    port map (
            O => \N__8339\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\
        );

    \I__741\ : InMux
    port map (
            O => \N__8336\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\
        );

    \I__740\ : InMux
    port map (
            O => \N__8333\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\
        );

    \I__739\ : InMux
    port map (
            O => \N__8330\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\
        );

    \I__738\ : InMux
    port map (
            O => \N__8327\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\
        );

    \I__737\ : InMux
    port map (
            O => \N__8324\,
            I => \bfn_1_19_0_\
        );

    \I__736\ : InMux
    port map (
            O => \N__8321\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\
        );

    \I__735\ : InMux
    port map (
            O => \N__8318\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\
        );

    \I__734\ : InMux
    port map (
            O => \N__8315\,
            I => \N__8312\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__8312\,
            I => \N__8309\
        );

    \I__732\ : Span12Mux_s3_v
    port map (
            O => \N__8309\,
            I => \N__8306\
        );

    \I__731\ : Span12Mux_h
    port map (
            O => \N__8306\,
            I => \N__8303\
        );

    \I__730\ : Span12Mux_h
    port map (
            O => \N__8303\,
            I => \N__8297\
        );

    \I__729\ : InMux
    port map (
            O => \N__8302\,
            I => \N__8294\
        );

    \I__728\ : InMux
    port map (
            O => \N__8301\,
            I => \N__8291\
        );

    \I__727\ : InMux
    port map (
            O => \N__8300\,
            I => \N__8288\
        );

    \I__726\ : Odrv12
    port map (
            O => \N__8297\,
            I => \CONSTANT_ONE_NET\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__8294\,
            I => \CONSTANT_ONE_NET\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__8291\,
            I => \CONSTANT_ONE_NET\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__8288\,
            I => \CONSTANT_ONE_NET\
        );

    \I__722\ : InMux
    port map (
            O => \N__8279\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\
        );

    \I__721\ : InMux
    port map (
            O => \N__8276\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\
        );

    \I__720\ : InMux
    port map (
            O => \N__8273\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\
        );

    \I__719\ : InMux
    port map (
            O => \N__8270\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\
        );

    \I__718\ : InMux
    port map (
            O => \N__8267\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\
        );

    \I__717\ : InMux
    port map (
            O => \N__8264\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\
        );

    \I__716\ : InMux
    port map (
            O => \N__8261\,
            I => \bfn_1_18_0_\
        );

    \I__715\ : InMux
    port map (
            O => \N__8258\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\
        );

    \I__714\ : InMux
    port map (
            O => \N__8255\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\
        );

    \I__713\ : InMux
    port map (
            O => \N__8252\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\
        );

    \I__712\ : InMux
    port map (
            O => \N__8249\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\
        );

    \I__711\ : InMux
    port map (
            O => \N__8246\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\
        );

    \I__710\ : InMux
    port map (
            O => \N__8243\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\
        );

    \I__709\ : InMux
    port map (
            O => \N__8240\,
            I => \bfn_1_16_0_\
        );

    \I__708\ : InMux
    port map (
            O => \N__8237\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\
        );

    \I__707\ : InMux
    port map (
            O => \N__8234\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\
        );

    \I__706\ : InMux
    port map (
            O => \N__8231\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\
        );

    \I__705\ : InMux
    port map (
            O => \N__8228\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\
        );

    \I__704\ : InMux
    port map (
            O => \N__8225\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\
        );

    \I__703\ : InMux
    port map (
            O => \N__8222\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\
        );

    \I__702\ : InMux
    port map (
            O => \N__8219\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\
        );

    \I__701\ : InMux
    port map (
            O => \N__8216\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\
        );

    \I__700\ : InMux
    port map (
            O => \N__8213\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\
        );

    \I__699\ : InMux
    port map (
            O => \N__8210\,
            I => \bfn_1_15_0_\
        );

    \I__698\ : InMux
    port map (
            O => \N__8207\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\
        );

    \I__697\ : InMux
    port map (
            O => \N__8204\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\
        );

    \I__696\ : InMux
    port map (
            O => \N__8201\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\
        );

    \I__695\ : InMux
    port map (
            O => \N__8198\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\
        );

    \IN_MUX_bfv_8_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_17_0_\
        );

    \IN_MUX_bfv_8_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_8_18_0_\
        );

    \IN_MUX_bfv_8_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_8_19_0_\
        );

    \IN_MUX_bfv_2_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_23_0_\
        );

    \IN_MUX_bfv_2_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_2_24_0_\
        );

    \IN_MUX_bfv_2_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_2_25_0_\
        );

    \IN_MUX_bfv_1_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_17_0_\
        );

    \IN_MUX_bfv_1_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_1_18_0_\
        );

    \IN_MUX_bfv_1_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_1_19_0_\
        );

    \IN_MUX_bfv_1_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_14_0_\
        );

    \IN_MUX_bfv_1_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_1_15_0_\
        );

    \IN_MUX_bfv_1_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_1_16_0_\
        );

    \IN_MUX_bfv_5_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_17_0_\
        );

    \IN_MUX_bfv_5_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8\,
            carryinitout => \bfn_5_18_0_\
        );

    \IN_MUX_bfv_5_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16\,
            carryinitout => \bfn_5_19_0_\
        );

    \IN_MUX_bfv_3_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_25_0_\
        );

    \IN_MUX_bfv_3_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8\,
            carryinitout => \bfn_3_26_0_\
        );

    \IN_MUX_bfv_3_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16\,
            carryinitout => \bfn_3_27_0_\
        );

    \IN_MUX_bfv_3_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_19_0_\
        );

    \IN_MUX_bfv_3_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            carryinitout => \bfn_3_20_0_\
        );

    \IN_MUX_bfv_3_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            carryinitout => \bfn_3_21_0_\
        );

    \IN_MUX_bfv_3_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_15_0_\
        );

    \IN_MUX_bfv_3_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            carryinitout => \bfn_3_16_0_\
        );

    \IN_MUX_bfv_3_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            carryinitout => \bfn_3_17_0_\
        );

    \IN_MUX_bfv_9_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_13_0_\
        );

    \IN_MUX_bfv_9_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_9_14_0_\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_9_15_0_\
        );

    \IN_MUX_bfv_9_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_9_16_0_\
        );

    \IN_MUX_bfv_8_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_13_0_\
        );

    \IN_MUX_bfv_8_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            carryinitout => \bfn_8_14_0_\
        );

    \IN_MUX_bfv_8_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            carryinitout => \bfn_8_15_0_\
        );

    \IN_MUX_bfv_8_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            carryinitout => \bfn_8_16_0_\
        );

    \IN_MUX_bfv_10_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_21_0_\
        );

    \IN_MUX_bfv_10_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_10_22_0_\
        );

    \IN_MUX_bfv_10_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_10_23_0_\
        );

    \IN_MUX_bfv_10_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_10_24_0_\
        );

    \IN_MUX_bfv_9_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_21_0_\
        );

    \IN_MUX_bfv_9_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            carryinitout => \bfn_9_22_0_\
        );

    \IN_MUX_bfv_9_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            carryinitout => \bfn_9_23_0_\
        );

    \IN_MUX_bfv_9_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            carryinitout => \bfn_9_24_0_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__19934\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.delay_tr_timer.N_255_i_g\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__20702\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.delay_hc_timer.N_253_i_g\
        );

    \osc\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b10"
        )
    port map (
            CLKHFPU => \N__8300\,
            CLKHFEN => \N__8302\,
            CLKHF => clk_12mhz
        );

    \rgb_drv\ : SB_RGBA_DRV
    generic map (
            RGB2_CURRENT => "0b111111",
            CURRENT_MODE => "0b0",
            RGB0_CURRENT => "0b111111",
            RGB1_CURRENT => "0b111111"
        )
    port map (
            RGBLEDEN => \N__8301\,
            RGB2PWM => \N__8387\,
            RGB1 => rgb_g_wire,
            CURREN => \N__8315\,
            RGB2 => rgb_b_wire,
            RGB1PWM => \N__8393\,
            RGB0PWM => \N__20466\,
            RGB0 => rgb_r_wire
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__20048\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.delay_tr_timer.N_256_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8915\,
            in2 => \N__9110\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_14_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8885\,
            in2 => \_gnd_net_\,
            in3 => \N__8198\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8864\,
            in2 => \N__8468\,
            in3 => \N__8228\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8843\,
            in2 => \_gnd_net_\,
            in3 => \N__8225\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8822\,
            in2 => \_gnd_net_\,
            in3 => \N__8222\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8801\,
            in2 => \_gnd_net_\,
            in3 => \N__8219\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8780\,
            in2 => \_gnd_net_\,
            in3 => \N__8216\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9086\,
            in3 => \N__8213\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9062\,
            in2 => \_gnd_net_\,
            in3 => \N__8210\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_1_15_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9041\,
            in2 => \_gnd_net_\,
            in3 => \N__8207\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9020\,
            in2 => \_gnd_net_\,
            in3 => \N__8204\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8999\,
            in2 => \_gnd_net_\,
            in3 => \N__8201\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8978\,
            in2 => \_gnd_net_\,
            in3 => \N__8252\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8957\,
            in2 => \_gnd_net_\,
            in3 => \N__8249\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8936\,
            in2 => \_gnd_net_\,
            in3 => \N__8246\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9212\,
            in2 => \_gnd_net_\,
            in3 => \N__8243\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9191\,
            in2 => \_gnd_net_\,
            in3 => \N__8240\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_1_16_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9158\,
            in2 => \_gnd_net_\,
            in3 => \N__8237\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9137\,
            in2 => \_gnd_net_\,
            in3 => \N__8234\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10130\,
            in2 => \N__10145\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_17_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9281\,
            in3 => \N__8231\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9257\,
            in2 => \N__8480\,
            in3 => \N__8279\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9233\,
            in2 => \_gnd_net_\,
            in3 => \N__8276\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9893\,
            in2 => \_gnd_net_\,
            in3 => \N__8273\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_1_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9872\,
            in2 => \_gnd_net_\,
            in3 => \N__8270\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9851\,
            in2 => \_gnd_net_\,
            in3 => \N__8267\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_1_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9830\,
            in2 => \_gnd_net_\,
            in3 => \N__8264\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_1_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9809\,
            in2 => \_gnd_net_\,
            in3 => \N__8261\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\,
            ltout => OPEN,
            carryin => \bfn_1_18_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_1_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9788\,
            in2 => \_gnd_net_\,
            in3 => \N__8258\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_1_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9766\,
            in2 => \_gnd_net_\,
            in3 => \N__8255\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_1_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9743\,
            in2 => \_gnd_net_\,
            in3 => \N__8339\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_1_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10058\,
            in2 => \_gnd_net_\,
            in3 => \N__8336\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_1_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10037\,
            in2 => \_gnd_net_\,
            in3 => \N__8333\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_1_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10016\,
            in2 => \_gnd_net_\,
            in3 => \N__8330\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_1_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9995\,
            in2 => \_gnd_net_\,
            in3 => \N__8327\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_1_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9968\,
            in2 => \_gnd_net_\,
            in3 => \N__8324\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\,
            ltout => OPEN,
            carryin => \bfn_1_19_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_1_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9941\,
            in2 => \_gnd_net_\,
            in3 => \N__8321\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_1_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9914\,
            in2 => \_gnd_net_\,
            in3 => \N__8318\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_1_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_drv_RNO_LC_1_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__20465\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13085\,
            lcout => \rgb_drv_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_drv_RNO_0_LC_1_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__20464\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13084\,
            lcout => \N_39_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__9601\,
            in1 => \N__11915\,
            in2 => \N__9722\,
            in3 => \N__8381\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20942\,
            ce => 'H',
            sr => \N__20382\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__9710\,
            in1 => \N__9605\,
            in2 => \N__11941\,
            in3 => \N__8375\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20942\,
            ce => 'H',
            sr => \N__20382\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__9708\,
            in1 => \N__9603\,
            in2 => \N__11939\,
            in3 => \N__8369\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20942\,
            ce => 'H',
            sr => \N__20382\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__9599\,
            in1 => \N__11913\,
            in2 => \N__9720\,
            in3 => \N__8363\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20942\,
            ce => 'H',
            sr => \N__20382\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__9707\,
            in1 => \N__9602\,
            in2 => \N__11938\,
            in3 => \N__8357\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20942\,
            ce => 'H',
            sr => \N__20382\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__9600\,
            in1 => \N__11914\,
            in2 => \N__9721\,
            in3 => \N__8351\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20942\,
            ce => 'H',
            sr => \N__20382\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__9709\,
            in1 => \N__9604\,
            in2 => \N__11940\,
            in3 => \N__8345\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20942\,
            ce => 'H',
            sr => \N__20382\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__9607\,
            in1 => \N__9700\,
            in2 => \N__11933\,
            in3 => \N__8453\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20940\,
            ce => 'H',
            sr => \N__20390\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__9695\,
            in1 => \N__11902\,
            in2 => \N__8447\,
            in3 => \N__9610\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20940\,
            ce => 'H',
            sr => \N__20390\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__9606\,
            in1 => \N__9699\,
            in2 => \N__11932\,
            in3 => \N__8438\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20940\,
            ce => 'H',
            sr => \N__20390\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__9696\,
            in1 => \N__11903\,
            in2 => \N__8432\,
            in3 => \N__9611\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20940\,
            ce => 'H',
            sr => \N__20390\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__9609\,
            in1 => \N__9702\,
            in2 => \N__11935\,
            in3 => \N__8423\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20940\,
            ce => 'H',
            sr => \N__20390\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__9697\,
            in1 => \N__11904\,
            in2 => \N__8417\,
            in3 => \N__9612\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20940\,
            ce => 'H',
            sr => \N__20390\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__9608\,
            in1 => \N__9701\,
            in2 => \N__11934\,
            in3 => \N__8408\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20940\,
            ce => 'H',
            sr => \N__20390\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__9698\,
            in1 => \N__11901\,
            in2 => \N__8402\,
            in3 => \N__9613\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20940\,
            ce => 'H',
            sr => \N__20390\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010100010"
        )
    port map (
            in0 => \N__8489\,
            in1 => \N__9706\,
            in2 => \N__9614\,
            in3 => \N__11912\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20938\,
            ce => 'H',
            sr => \N__20395\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__9594\,
            in1 => \N__9705\,
            in2 => \N__11937\,
            in3 => \N__8510\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20938\,
            ce => 'H',
            sr => \N__20395\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__9593\,
            in1 => \N__9704\,
            in2 => \N__11936\,
            in3 => \N__8504\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20938\,
            ce => 'H',
            sr => \N__20395\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__9592\,
            in1 => \N__9703\,
            in2 => \N__8498\,
            in3 => \N__11911\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20938\,
            ce => 'H',
            sr => \N__20395\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__12169\,
            in1 => \N__9349\,
            in2 => \_gnd_net_\,
            in3 => \N__9475\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_2_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__11042\,
            in1 => \N__8914\,
            in2 => \_gnd_net_\,
            in3 => \N__11005\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9348\,
            in2 => \_gnd_net_\,
            in3 => \N__9474\,
            lcout => \phase_controller_inst1.stoper_tr.time_passed11\,
            ltout => \phase_controller_inst1.stoper_tr.time_passed11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_2_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8483\,
            in3 => \N__11080\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9643\,
            in2 => \_gnd_net_\,
            in3 => \N__9539\,
            lcout => \phase_controller_inst1.stoper_hc.time_passed11\,
            ltout => \phase_controller_inst1.stoper_hc.time_passed11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_2_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8471\,
            in3 => \N__11041\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__9485\,
            in1 => \N__12231\,
            in2 => \N__9413\,
            in3 => \N__8570\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20933\,
            ce => 'H',
            sr => \N__20405\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_2_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__9371\,
            in1 => \N__9484\,
            in2 => \N__12245\,
            in3 => \N__8564\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20933\,
            ce => 'H',
            sr => \N__20405\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__9482\,
            in1 => \N__12230\,
            in2 => \N__9412\,
            in3 => \N__8558\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20933\,
            ce => 'H',
            sr => \N__20405\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__9369\,
            in1 => \N__9479\,
            in2 => \N__12243\,
            in3 => \N__8552\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20933\,
            ce => 'H',
            sr => \N__20405\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__9480\,
            in1 => \N__12228\,
            in2 => \N__9410\,
            in3 => \N__8546\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20933\,
            ce => 'H',
            sr => \N__20405\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_2_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__9370\,
            in1 => \N__9483\,
            in2 => \N__12244\,
            in3 => \N__8540\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20933\,
            ce => 'H',
            sr => \N__20405\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_2_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__9481\,
            in1 => \N__12229\,
            in2 => \N__9411\,
            in3 => \N__8534\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20933\,
            ce => 'H',
            sr => \N__20405\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__9373\,
            in1 => \N__9488\,
            in2 => \N__12225\,
            in3 => \N__8528\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20927\,
            ce => 'H',
            sr => \N__20410\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_2_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__9487\,
            in1 => \N__12183\,
            in2 => \N__9406\,
            in3 => \N__8522\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20927\,
            ce => 'H',
            sr => \N__20410\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_2_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__9375\,
            in1 => \N__9492\,
            in2 => \N__12227\,
            in3 => \N__8516\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20927\,
            ce => 'H',
            sr => \N__20410\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_2_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__9491\,
            in1 => \N__12185\,
            in2 => \N__9408\,
            in3 => \N__8618\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20927\,
            ce => 'H',
            sr => \N__20410\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_2_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__9372\,
            in1 => \N__9486\,
            in2 => \N__12224\,
            in3 => \N__8612\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20927\,
            ce => 'H',
            sr => \N__20410\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_2_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__9493\,
            in1 => \N__12186\,
            in2 => \N__9409\,
            in3 => \N__8606\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20927\,
            ce => 'H',
            sr => \N__20410\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_2_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__9374\,
            in1 => \N__9490\,
            in2 => \N__12226\,
            in3 => \N__8600\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20927\,
            ce => 'H',
            sr => \N__20410\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_2_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__9489\,
            in1 => \N__12184\,
            in2 => \N__9407\,
            in3 => \N__8594\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20927\,
            ce => 'H',
            sr => \N__20410\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_2_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__9509\,
            in1 => \N__9393\,
            in2 => \N__12220\,
            in3 => \N__10109\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20923\,
            ce => 'H',
            sr => \N__20413\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_2_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__9392\,
            in1 => \N__9508\,
            in2 => \N__12223\,
            in3 => \N__8588\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20923\,
            ce => 'H',
            sr => \N__20413\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_2_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__9391\,
            in1 => \N__9507\,
            in2 => \N__12222\,
            in3 => \N__8582\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20923\,
            ce => 'H',
            sr => \N__20413\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_2_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__9390\,
            in1 => \N__9506\,
            in2 => \N__12221\,
            in3 => \N__8576\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20923\,
            ce => 'H',
            sr => \N__20413\
        );

    \phase_controller_inst1.stoper_tr.target_time_18_LC_2_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16793\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20919\,
            ce => \N__11262\,
            sr => \N__20415\
        );

    \phase_controller_inst1.stoper_tr.target_time_17_LC_2_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16754\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20919\,
            ce => \N__11262\,
            sr => \N__20415\
        );

    \phase_controller_inst1.stoper_tr.target_time_19_LC_2_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18551\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20919\,
            ce => \N__11262\,
            sr => \N__20415\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_2_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10241\,
            in2 => \N__10907\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_23_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_2_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10211\,
            in2 => \_gnd_net_\,
            in3 => \N__8633\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_2_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10193\,
            in2 => \N__8732\,
            in3 => \N__8630\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_2_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10172\,
            in2 => \_gnd_net_\,
            in3 => \N__8627\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_2_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10460\,
            in2 => \_gnd_net_\,
            in3 => \N__8624\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_2_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10439\,
            in2 => \_gnd_net_\,
            in3 => \N__8621\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_2_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10418\,
            in2 => \_gnd_net_\,
            in3 => \N__8660\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_2_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10397\,
            in2 => \_gnd_net_\,
            in3 => \N__8657\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_2_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10376\,
            in2 => \_gnd_net_\,
            in3 => \N__8654\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9\,
            ltout => OPEN,
            carryin => \bfn_2_24_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_2_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10352\,
            in2 => \_gnd_net_\,
            in3 => \N__8651\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_2_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10328\,
            in2 => \_gnd_net_\,
            in3 => \N__8648\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_2_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10304\,
            in2 => \_gnd_net_\,
            in3 => \N__8645\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_2_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10618\,
            in2 => \_gnd_net_\,
            in3 => \N__8642\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_2_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10594\,
            in2 => \_gnd_net_\,
            in3 => \N__8639\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_2_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10570\,
            in2 => \_gnd_net_\,
            in3 => \N__8636\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_2_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10546\,
            in2 => \_gnd_net_\,
            in3 => \N__8711\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_2_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10523\,
            in2 => \_gnd_net_\,
            in3 => \N__8708\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17\,
            ltout => OPEN,
            carryin => \bfn_2_25_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_2_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10502\,
            in2 => \_gnd_net_\,
            in3 => \N__8705\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_2_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10481\,
            in2 => \_gnd_net_\,
            in3 => \N__8702\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_17_LC_2_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__10775\,
            in1 => \N__10874\,
            in2 => \N__12913\,
            in3 => \N__8699\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20894\,
            ce => 'H',
            sr => \N__20424\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_12_LC_2_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__10871\,
            in1 => \N__10779\,
            in2 => \N__12910\,
            in3 => \N__8693\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20894\,
            ce => 'H',
            sr => \N__20424\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_9_LC_2_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__10777\,
            in1 => \N__10875\,
            in2 => \N__12914\,
            in3 => \N__8684\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20894\,
            ce => 'H',
            sr => \N__20424\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_1_LC_2_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010100010"
        )
    port map (
            in0 => \N__8717\,
            in1 => \N__12892\,
            in2 => \N__10892\,
            in3 => \N__10781\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20894\,
            ce => 'H',
            sr => \N__20424\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_10_LC_2_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__10774\,
            in1 => \N__10873\,
            in2 => \N__12912\,
            in3 => \N__8675\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20894\,
            ce => 'H',
            sr => \N__20424\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_19_LC_2_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__10872\,
            in1 => \N__10780\,
            in2 => \N__12911\,
            in3 => \N__8666\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20894\,
            ce => 'H',
            sr => \N__20424\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_18_LC_2_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__10776\,
            in1 => \N__12888\,
            in2 => \N__8753\,
            in3 => \N__10879\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20894\,
            ce => 'H',
            sr => \N__20424\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_11_LC_2_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__10870\,
            in1 => \N__10778\,
            in2 => \N__12909\,
            in3 => \N__8744\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20894\,
            ce => 'H',
            sr => \N__20424\
        );

    \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_2_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10816\,
            in2 => \_gnd_net_\,
            in3 => \N__10709\,
            lcout => \phase_controller_slave.stoper_hc.time_passed11\,
            ltout => \phase_controller_slave.stoper_hc.time_passed11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_2_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8735\,
            in3 => \N__11962\,
            lcout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_2_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__11963\,
            in1 => \N__11992\,
            in2 => \_gnd_net_\,
            in3 => \N__10240\,
            lcout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.stoper_state_0_LC_2_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__10720\,
            in1 => \N__10842\,
            in2 => \N__12904\,
            in3 => \N__11964\,
            lcout => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20880\,
            ce => \N__20191\,
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.stoper_state_1_LC_2_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001010000"
        )
    port map (
            in0 => \N__11965\,
            in1 => \N__12862\,
            in2 => \N__10880\,
            in3 => \N__10721\,
            lcout => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20880\,
            ce => \N__20191\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_LC_3_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11442\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13883\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20941\,
            ce => \N__11146\,
            sr => \N__20376\
        );

    \phase_controller_inst1.stoper_hc.target_time_18_LC_3_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13934\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20941\,
            ce => \N__11146\,
            sr => \N__20376\
        );

    \phase_controller_inst1.stoper_hc.target_time_8_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11443\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13847\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20941\,
            ce => \N__11146\,
            sr => \N__20376\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_3_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10643\,
            in2 => \N__8894\,
            in3 => \N__8910\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_3_15_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_3_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10652\,
            in2 => \N__8873\,
            in3 => \N__8884\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10988\,
            in2 => \N__8852\,
            in3 => \N__8863\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_3_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10634\,
            in2 => \N__8831\,
            in3 => \N__8842\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10964\,
            in2 => \N__8810\,
            in3 => \N__8821\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10628\,
            in2 => \N__8789\,
            in3 => \N__8800\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_3_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__8779\,
            in1 => \N__8768\,
            in2 => \N__8762\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_3_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9095\,
            in2 => \N__9071\,
            in3 => \N__9082\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_3_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11156\,
            in2 => \N__9050\,
            in3 => \N__9061\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_3_16_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_3_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10922\,
            in2 => \N__9029\,
            in3 => \N__9040\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10934\,
            in2 => \N__9008\,
            in3 => \N__9019\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_3_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__8998\,
            in1 => \N__10979\,
            in2 => \N__8987\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_3_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__8977\,
            in1 => \N__10949\,
            in2 => \N__8966\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_3_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10955\,
            in2 => \N__8945\,
            in3 => \N__8956\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_3_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11165\,
            in2 => \N__8924\,
            in3 => \N__8935\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_3_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10973\,
            in2 => \N__9200\,
            in3 => \N__9211\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10940\,
            in2 => \N__9179\,
            in3 => \N__9190\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_3_17_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_3_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9170\,
            in2 => \N__9146\,
            in3 => \N__9157\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_3_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10928\,
            in2 => \N__9125\,
            in3 => \N__9136\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_3_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9116\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_3_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9113\,
            in3 => \N__11004\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_3_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__9645\,
            in1 => \N__11882\,
            in2 => \_gnd_net_\,
            in3 => \N__9540\,
            lcout => \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__9350\,
            in1 => \N__12170\,
            in2 => \_gnd_net_\,
            in3 => \N__9505\,
            lcout => \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_3_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__9644\,
            in1 => \N__11881\,
            in2 => \_gnd_net_\,
            in3 => \N__9541\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_1_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001010000"
        )
    port map (
            in0 => \N__11044\,
            in1 => \N__11928\,
            in2 => \N__9598\,
            in3 => \N__9678\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20928\,
            ce => \N__20195\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_0_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__9677\,
            in1 => \N__9556\,
            in2 => \N__11942\,
            in3 => \N__11043\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20928\,
            ce => \N__20195\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_0_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__9376\,
            in1 => \N__9503\,
            in2 => \N__12241\,
            in3 => \N__11075\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20928\,
            ce => \N__20195\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_1_LC_3_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000001100100"
        )
    port map (
            in0 => \N__9377\,
            in1 => \N__9504\,
            in2 => \N__12242\,
            in3 => \N__11076\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20928\,
            ce => \N__20195\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11216\,
            in2 => \N__9290\,
            in3 => \N__10125\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_3_19_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_3_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11210\,
            in2 => \N__9266\,
            in3 => \N__9277\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11237\,
            in2 => \N__9242\,
            in3 => \N__9253\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11228\,
            in2 => \N__9221\,
            in3 => \N__9232\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_3_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11204\,
            in2 => \N__9881\,
            in3 => \N__9892\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_3_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11222\,
            in2 => \N__9860\,
            in3 => \N__9871\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11174\,
            in2 => \N__9839\,
            in3 => \N__9850\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_3_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11198\,
            in2 => \N__9818\,
            in3 => \N__9829\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_3_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11297\,
            in2 => \N__9797\,
            in3 => \N__9808\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_3_20_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_3_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11279\,
            in2 => \N__9776\,
            in3 => \N__9787\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_3_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11303\,
            in2 => \N__9752\,
            in3 => \N__9767\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_3_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11309\,
            in2 => \N__9731\,
            in3 => \N__9742\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_3_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11183\,
            in2 => \N__10046\,
            in3 => \N__10057\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_3_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11288\,
            in2 => \N__10025\,
            in3 => \N__10036\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_3_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11189\,
            in2 => \N__10004\,
            in3 => \N__10015\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_3_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11318\,
            in2 => \N__9983\,
            in3 => \N__9994\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_3_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9974\,
            in2 => \N__9956\,
            in3 => \N__9967\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_3_21_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_3_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9947\,
            in2 => \N__9929\,
            in3 => \N__9940\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_3_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9920\,
            in2 => \N__9902\,
            in3 => \N__9913\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_3_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10151\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_3_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10148\,
            in3 => \N__11116\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_3_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__11117\,
            in1 => \N__11071\,
            in2 => \_gnd_net_\,
            in3 => \N__10129\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_16_LC_3_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__10764\,
            in1 => \N__10883\,
            in2 => \N__12903\,
            in3 => \N__10103\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20902\,
            ce => 'H',
            sr => \N__20416\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_15_LC_3_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__10881\,
            in1 => \N__12854\,
            in2 => \N__10097\,
            in3 => \N__10765\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20902\,
            ce => 'H',
            sr => \N__20416\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_14_LC_3_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__10763\,
            in1 => \N__10882\,
            in2 => \N__12902\,
            in3 => \N__10088\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20902\,
            ce => 'H',
            sr => \N__20416\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_6_LC_3_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__10886\,
            in1 => \N__12880\,
            in2 => \N__10082\,
            in3 => \N__10772\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20898\,
            ce => 'H',
            sr => \N__20419\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_7_LC_3_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__10769\,
            in1 => \N__10891\,
            in2 => \N__12908\,
            in3 => \N__10073\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20898\,
            ce => 'H',
            sr => \N__20419\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_3_LC_3_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__10884\,
            in1 => \N__12878\,
            in2 => \N__10067\,
            in3 => \N__10770\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20898\,
            ce => 'H',
            sr => \N__20419\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_13_LC_3_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__10766\,
            in1 => \N__10888\,
            in2 => \N__12905\,
            in3 => \N__10277\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20898\,
            ce => 'H',
            sr => \N__20419\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_8_LC_3_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__10887\,
            in1 => \N__12881\,
            in2 => \N__10271\,
            in3 => \N__10773\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20898\,
            ce => 'H',
            sr => \N__20419\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_5_LC_3_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__10768\,
            in1 => \N__10890\,
            in2 => \N__12907\,
            in3 => \N__10262\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20898\,
            ce => 'H',
            sr => \N__20419\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_4_LC_3_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__10885\,
            in1 => \N__12879\,
            in2 => \N__10256\,
            in3 => \N__10771\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20898\,
            ce => 'H',
            sr => \N__20419\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_2_LC_3_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__10767\,
            in1 => \N__10889\,
            in2 => \N__12906\,
            in3 => \N__10247\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20898\,
            ce => 'H',
            sr => \N__20419\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_3_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11582\,
            in2 => \N__10220\,
            in3 => \N__10236\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_3_25_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_3_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10199\,
            in2 => \N__11534\,
            in3 => \N__10210\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_3_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11450\,
            in2 => \N__10181\,
            in3 => \N__10192\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_3_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11525\,
            in2 => \N__10160\,
            in3 => \N__10171\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_3_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11594\,
            in2 => \N__10448\,
            in3 => \N__10459\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_3_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10438\,
            in1 => \N__11564\,
            in2 => \N__10427\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_3_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10417\,
            in1 => \N__11576\,
            in2 => \N__10406\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_3_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11369\,
            in2 => \N__10385\,
            in3 => \N__10396\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_3_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11726\,
            in2 => \N__10361\,
            in3 => \N__10372\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_3_26_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_3_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11765\,
            in2 => \N__10337\,
            in3 => \N__10348\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_3_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11663\,
            in2 => \N__10313\,
            in3 => \N__10324\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_3_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11759\,
            in2 => \N__10286\,
            in3 => \N__10303\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_3_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11771\,
            in2 => \N__10604\,
            in3 => \N__10619\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_3_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11618\,
            in2 => \N__10580\,
            in3 => \N__10595\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_3_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11360\,
            in2 => \N__10556\,
            in3 => \N__10571\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_3_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11612\,
            in2 => \N__10532\,
            in3 => \N__10547\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_3_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11600\,
            in2 => \N__10511\,
            in3 => \N__10522\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_3_27_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_3_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12050\,
            in2 => \N__10490\,
            in3 => \N__10501\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_3_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11606\,
            in2 => \N__10469\,
            in3 => \N__10480\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_3_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10913\,
            lcout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_3_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10910\,
            in3 => \N__11991\,
            lcout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_3_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__10817\,
            in1 => \N__12853\,
            in2 => \_gnd_net_\,
            in3 => \N__10710\,
            lcout => \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_3_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__12861\,
            in1 => \N__10818\,
            in2 => \_gnd_net_\,
            in3 => \N__10711\,
            lcout => \phase_controller_slave.stoper_hc.time_passed_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_3_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__10679\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_clk_12mhz_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_2_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__11558\,
            in1 => \N__13343\,
            in2 => \N__11444\,
            in3 => \N__11515\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20936\,
            ce => \N__11147\,
            sr => \N__20377\
        );

    \phase_controller_inst1.stoper_hc.target_time_1_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__11514\,
            in1 => \N__11434\,
            in2 => \N__13652\,
            in3 => \N__11557\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20936\,
            ce => \N__11147\,
            sr => \N__20377\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__11439\,
            in1 => \N__11517\,
            in2 => \_gnd_net_\,
            in3 => \N__13703\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20936\,
            ce => \N__11147\,
            sr => \N__20377\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__11519\,
            in1 => \N__11441\,
            in2 => \_gnd_net_\,
            in3 => \N__14099\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20936\,
            ce => \N__11147\,
            sr => \N__20377\
        );

    \phase_controller_inst1.stoper_hc.target_time_3_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__11438\,
            in1 => \N__11516\,
            in2 => \N__13742\,
            in3 => \N__11468\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20936\,
            ce => \N__11147\,
            sr => \N__20377\
        );

    \phase_controller_inst1.stoper_hc.target_time_12_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11712\,
            in2 => \_gnd_net_\,
            in3 => \N__13772\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20936\,
            ce => \N__11147\,
            sr => \N__20377\
        );

    \phase_controller_inst1.stoper_hc.target_time_16_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14024\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20936\,
            ce => \N__11147\,
            sr => \N__20377\
        );

    \phase_controller_inst1.stoper_hc.target_time_5_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__11518\,
            in1 => \N__13382\,
            in2 => \_gnd_net_\,
            in3 => \N__11440\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20936\,
            ce => \N__11147\,
            sr => \N__20377\
        );

    \phase_controller_inst1.stoper_hc.target_time_14_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__13555\,
            in1 => \N__11650\,
            in2 => \_gnd_net_\,
            in3 => \N__13979\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20934\,
            ce => \N__11145\,
            sr => \N__20383\
        );

    \phase_controller_inst1.stoper_hc.target_time_13_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11708\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15776\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20934\,
            ce => \N__11145\,
            sr => \N__20383\
        );

    \phase_controller_inst1.stoper_hc.target_time_17_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14066\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20934\,
            ce => \N__11145\,
            sr => \N__20383\
        );

    \phase_controller_inst1.stoper_hc.target_time_11_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11707\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13802\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20934\,
            ce => \N__11145\,
            sr => \N__20383\
        );

    \phase_controller_inst1.stoper_hc.target_time_19_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13498\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20934\,
            ce => \N__11145\,
            sr => \N__20383\
        );

    \phase_controller_inst1.stoper_hc.target_time_10_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11706\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13619\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20934\,
            ce => \N__11145\,
            sr => \N__20383\
        );

    \phase_controller_inst1.stoper_hc.target_time_15_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13554\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11651\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20934\,
            ce => \N__11145\,
            sr => \N__20383\
        );

    \phase_controller_inst1.stoper_hc.target_time_9_LC_4_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111110101011"
        )
    port map (
            in0 => \N__13589\,
            in1 => \N__11750\,
            in2 => \N__11714\,
            in3 => \N__13556\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20934\,
            ce => \N__11145\,
            sr => \N__20383\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_4_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__15468\,
            in1 => \N__15146\,
            in2 => \N__15342\,
            in3 => \N__14309\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20929\,
            ce => 'H',
            sr => \N__20391\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_1_LC_4_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__15141\,
            in1 => \N__15316\,
            in2 => \N__15479\,
            in3 => \N__12617\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20929\,
            ce => 'H',
            sr => \N__20391\
        );

    \phase_controller_inst1.stoper_tr.time_passed_LC_4_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__12378\,
            in1 => \N__11115\,
            in2 => \N__11093\,
            in3 => \N__11081\,
            lcout => \phase_controller_inst1.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20929\,
            ce => 'H',
            sr => \N__20391\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_6_LC_4_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__15144\,
            in1 => \N__15319\,
            in2 => \N__14243\,
            in3 => \N__15471\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20929\,
            ce => 'H',
            sr => \N__20391\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_2_LC_4_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__15467\,
            in1 => \N__15145\,
            in2 => \N__15341\,
            in3 => \N__14387\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20929\,
            ce => 'H',
            sr => \N__20391\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_5_LC_4_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__15143\,
            in1 => \N__15318\,
            in2 => \N__14276\,
            in3 => \N__15470\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20929\,
            ce => 'H',
            sr => \N__20391\
        );

    \phase_controller_inst1.stoper_hc.time_passed_LC_4_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110111000000"
        )
    port map (
            in0 => \N__11045\,
            in1 => \N__12314\,
            in2 => \N__11021\,
            in3 => \N__11009\,
            lcout => \phase_controller_inst1.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20929\,
            ce => 'H',
            sr => \N__20391\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_3_LC_4_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__15142\,
            in1 => \N__15317\,
            in2 => \N__14342\,
            in3 => \N__15469\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20929\,
            ce => 'H',
            sr => \N__20391\
        );

    \phase_controller_slave.stoper_tr.target_time_3_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__14827\,
            in1 => \N__14717\,
            in2 => \N__16420\,
            in3 => \N__17099\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20924\,
            ce => \N__12666\,
            sr => \N__20396\
        );

    \phase_controller_slave.stoper_tr.target_time_9_LC_4_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011111101"
        )
    port map (
            in0 => \N__16564\,
            in1 => \N__16997\,
            in2 => \N__16532\,
            in3 => \N__12737\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20924\,
            ce => \N__12666\,
            sr => \N__20396\
        );

    \phase_controller_slave.stoper_tr.target_time_8_LC_4_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14720\,
            in2 => \_gnd_net_\,
            in3 => \N__18717\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20924\,
            ce => \N__12666\,
            sr => \N__20396\
        );

    \phase_controller_slave.stoper_tr.target_time_11_LC_4_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12735\,
            in2 => \_gnd_net_\,
            in3 => \N__16645\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20924\,
            ce => \N__12666\,
            sr => \N__20396\
        );

    \phase_controller_slave.stoper_tr.target_time_2_LC_4_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__14826\,
            in1 => \N__14887\,
            in2 => \N__16460\,
            in3 => \N__14716\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20924\,
            ce => \N__12666\,
            sr => \N__20396\
        );

    \phase_controller_slave.stoper_tr.target_time_12_LC_4_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12736\,
            in2 => \_gnd_net_\,
            in3 => \N__16672\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20924\,
            ce => \N__12666\,
            sr => \N__20396\
        );

    \phase_controller_slave.stoper_tr.target_time_6_LC_4_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__14828\,
            in1 => \N__14718\,
            in2 => \_gnd_net_\,
            in3 => \N__16819\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20924\,
            ce => \N__12666\,
            sr => \N__20396\
        );

    \phase_controller_slave.stoper_tr.target_time_7_LC_4_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__14719\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17851\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20924\,
            ce => \N__12666\,
            sr => \N__20396\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_LC_4_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__14696\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17855\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20920\,
            ce => \N__11269\,
            sr => \N__20398\
        );

    \phase_controller_inst1.stoper_tr.target_time_3_LC_4_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__14798\,
            in1 => \N__14692\,
            in2 => \N__16421\,
            in3 => \N__17092\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20920\,
            ce => \N__11269\,
            sr => \N__20398\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_LC_4_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__14693\,
            in1 => \N__14799\,
            in2 => \_gnd_net_\,
            in3 => \N__17069\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20920\,
            ce => \N__11269\,
            sr => \N__20398\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_LC_4_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000001111"
        )
    port map (
            in0 => \N__16820\,
            in1 => \_gnd_net_\,
            in2 => \N__14815\,
            in3 => \N__14695\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20920\,
            ce => \N__11269\,
            sr => \N__20398\
        );

    \phase_controller_inst1.stoper_tr.target_time_1_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__14690\,
            in1 => \N__14794\,
            in2 => \N__16487\,
            in3 => \N__14879\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20920\,
            ce => \N__11269\,
            sr => \N__20398\
        );

    \phase_controller_inst1.stoper_tr.target_time_2_LC_4_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__14880\,
            in1 => \N__16456\,
            in2 => \N__14814\,
            in3 => \N__14691\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20920\,
            ce => \N__11269\,
            sr => \N__20398\
        );

    \phase_controller_inst1.stoper_tr.target_time_5_LC_4_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__14694\,
            in1 => \N__14800\,
            in2 => \_gnd_net_\,
            in3 => \N__16931\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20920\,
            ce => \N__11269\,
            sr => \N__20398\
        );

    \phase_controller_inst1.stoper_tr.target_time_8_LC_4_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18725\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14697\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20920\,
            ce => \N__11269\,
            sr => \N__20398\
        );

    \phase_controller_inst1.stoper_tr.target_time_15_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__14759\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17000\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20913\,
            ce => \N__11273\,
            sr => \N__20406\
        );

    \phase_controller_inst1.stoper_tr.target_time_13_LC_4_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12726\,
            in2 => \_gnd_net_\,
            in3 => \N__16622\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20913\,
            ce => \N__11273\,
            sr => \N__20406\
        );

    \phase_controller_inst1.stoper_tr.target_time_16_LC_4_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16715\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20913\,
            ce => \N__11273\,
            sr => \N__20406\
        );

    \phase_controller_inst1.stoper_tr.target_time_12_LC_4_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12725\,
            in2 => \_gnd_net_\,
            in3 => \N__16676\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20913\,
            ce => \N__11273\,
            sr => \N__20406\
        );

    \phase_controller_inst1.stoper_tr.target_time_11_LC_4_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__12724\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16652\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20913\,
            ce => \N__11273\,
            sr => \N__20406\
        );

    \phase_controller_inst1.stoper_tr.target_time_9_LC_4_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100100011"
        )
    port map (
            in0 => \N__16998\,
            in1 => \N__12727\,
            in2 => \N__16565\,
            in3 => \N__16531\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20913\,
            ce => \N__11273\,
            sr => \N__20406\
        );

    \phase_controller_inst1.stoper_tr.target_time_14_LC_4_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__14758\,
            in1 => \N__16999\,
            in2 => \_gnd_net_\,
            in3 => \N__17039\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20913\,
            ce => \N__11273\,
            sr => \N__20406\
        );

    \phase_controller_inst1.stoper_tr.target_time_10_LC_4_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12723\,
            in2 => \_gnd_net_\,
            in3 => \N__16592\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20913\,
            ce => \N__11273\,
            sr => \N__20406\
        );

    \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_4_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__15221\,
            in1 => \N__15466\,
            in2 => \_gnd_net_\,
            in3 => \N__15140\,
            lcout => \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_f0_0_a2_4_3_LC_4_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13973\,
            in1 => \N__13377\,
            in2 => \N__13553\,
            in3 => \N__13692\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_6_f0_0_a2_4Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_f0_0_a2_3_3_LC_4_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13922\,
            in1 => \N__14061\,
            in2 => \N__13499\,
            in3 => \N__14019\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.target_time_6_f0_0_a2_3Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_f0_0_a2_3_LC_4_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11354\,
            in1 => \N__11327\,
            in2 => \N__11348\,
            in3 => \N__11339\,
            lcout => \phase_controller_inst1.stoper_hc.N_144\,
            ltout => \phase_controller_inst1.stoper_hc.N_144_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_f0_0_a3_1_LC_4_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011110000"
        )
    port map (
            in0 => \N__13725\,
            in1 => \_gnd_net_\,
            in2 => \N__11345\,
            in3 => \N__13332\,
            lcout => \phase_controller_inst1.stoper_hc.N_122\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_0_6_LC_4_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13761\,
            in1 => \N__13791\,
            in2 => \N__15771\,
            in3 => \N__13611\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_0Z0Z_6\,
            ltout => \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_9_LC_4_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__13584\,
            in1 => \_gnd_net_\,
            in2 => \N__11342\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2Z0Z_9\,
            ltout => \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_o2_6_LC_4_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010111011"
        )
    port map (
            in0 => \N__11634\,
            in1 => \N__13540\,
            in2 => \N__11333\,
            in3 => \N__13974\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_o2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_i_o2_15_LC_4_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__13926\,
            in1 => \N__14054\,
            in2 => \N__13490\,
            in3 => \N__14015\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_6_i_o2Z0Z_15\,
            ltout => \phase_controller_inst1.stoper_hc.target_time_6_i_o2Z0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_o2_9_LC_4_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110001"
        )
    port map (
            in0 => \N__13541\,
            in1 => \N__13966\,
            in2 => \N__11330\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_o2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_1_6_LC_4_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__13881\,
            in1 => \N__13846\,
            in2 => \_gnd_net_\,
            in3 => \N__14088\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_1Z0Z_6\,
            ltout => \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_1Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a3_0_6_LC_4_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__11742\,
            in1 => \_gnd_net_\,
            in2 => \N__11321\,
            in3 => \N__13542\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a3_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.target_time_5_LC_4_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__11403\,
            in1 => \N__11493\,
            in2 => \_gnd_net_\,
            in3 => \N__13378\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20895\,
            ce => \N__12044\,
            sr => \N__20417\
        );

    \phase_controller_slave.stoper_hc.target_time_1_LC_4_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__11489\,
            in1 => \N__11397\,
            in2 => \N__13648\,
            in3 => \N__11555\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20895\,
            ce => \N__12044\,
            sr => \N__20417\
        );

    \phase_controller_slave.stoper_hc.target_time_7_LC_4_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__13882\,
            in1 => \_gnd_net_\,
            in2 => \N__11415\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20895\,
            ce => \N__12044\,
            sr => \N__20417\
        );

    \phase_controller_slave.stoper_hc.target_time_6_LC_4_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__11494\,
            in1 => \N__11404\,
            in2 => \_gnd_net_\,
            in3 => \N__14095\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20895\,
            ce => \N__12044\,
            sr => \N__20417\
        );

    \phase_controller_slave.stoper_hc.target_time_2_LC_4_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__11556\,
            in1 => \N__13339\,
            in2 => \N__11414\,
            in3 => \N__11490\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20895\,
            ce => \N__12044\,
            sr => \N__20417\
        );

    \phase_controller_slave.stoper_hc.target_time_4_LC_4_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__11492\,
            in1 => \N__13699\,
            in2 => \_gnd_net_\,
            in3 => \N__11402\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20895\,
            ce => \N__12044\,
            sr => \N__20417\
        );

    \phase_controller_slave.stoper_hc.target_time_3_LC_4_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__11401\,
            in1 => \N__11491\,
            in2 => \N__13741\,
            in3 => \N__11467\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20895\,
            ce => \N__12044\,
            sr => \N__20417\
        );

    \phase_controller_slave.stoper_hc.target_time_8_LC_4_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11408\,
            in2 => \_gnd_net_\,
            in3 => \N__13842\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20895\,
            ce => \N__12044\,
            sr => \N__20417\
        );

    \phase_controller_slave.stoper_hc.target_time_15_LC_4_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__11644\,
            in1 => \N__13550\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20887\,
            ce => \N__12042\,
            sr => \N__20420\
        );

    \phase_controller_slave.stoper_hc.target_time_13_LC_4_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11702\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15772\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20887\,
            ce => \N__12042\,
            sr => \N__20420\
        );

    \phase_controller_slave.stoper_hc.target_time_10_LC_4_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11699\,
            in2 => \_gnd_net_\,
            in3 => \N__13618\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20887\,
            ce => \N__12042\,
            sr => \N__20420\
        );

    \phase_controller_slave.stoper_hc.target_time_12_LC_4_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11701\,
            in2 => \_gnd_net_\,
            in3 => \N__13768\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20887\,
            ce => \N__12042\,
            sr => \N__20420\
        );

    \phase_controller_slave.stoper_hc.target_time_9_LC_4_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100001011"
        )
    port map (
            in0 => \N__13552\,
            in1 => \N__11749\,
            in2 => \N__11713\,
            in3 => \N__13585\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20887\,
            ce => \N__12042\,
            sr => \N__20420\
        );

    \phase_controller_slave.stoper_hc.target_time_11_LC_4_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11700\,
            in2 => \_gnd_net_\,
            in3 => \N__13798\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20887\,
            ce => \N__12042\,
            sr => \N__20420\
        );

    \phase_controller_slave.stoper_hc.target_time_14_LC_4_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__13551\,
            in1 => \N__11643\,
            in2 => \_gnd_net_\,
            in3 => \N__13975\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20887\,
            ce => \N__12042\,
            sr => \N__20420\
        );

    \phase_controller_slave.stoper_hc.target_time_16_LC_4_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14020\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20881\,
            ce => \N__12043\,
            sr => \N__20422\
        );

    \phase_controller_slave.stoper_hc.target_time_19_LC_4_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13491\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20875\,
            ce => \N__12035\,
            sr => \N__20423\
        );

    \phase_controller_slave.stoper_hc.target_time_17_LC_4_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14062\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20875\,
            ce => \N__12035\,
            sr => \N__20423\
        );

    \phase_controller_slave.stoper_hc.target_time_18_LC_4_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13933\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20875\,
            ce => \N__12035\,
            sr => \N__20423\
        );

    \phase_controller_slave.stoper_hc.time_passed_LC_4_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__13281\,
            in1 => \N__11999\,
            in2 => \N__11975\,
            in3 => \N__11966\,
            lcout => \phase_controller_slave.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20870\,
            ce => 'H',
            sr => \N__20425\
        );

    \phase_controller_inst1.state_2_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__13217\,
            in1 => \N__12340\,
            in2 => \N__16890\,
            in3 => \N__12323\,
            lcout => \phase_controller_inst1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20939\,
            ce => 'H',
            sr => \N__20368\
        );

    \phase_controller_inst1.state_3_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111011111110"
        )
    port map (
            in0 => \N__11786\,
            in1 => \N__12257\,
            in2 => \N__16891\,
            in3 => \N__13216\,
            lcout => \phase_controller_inst1.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20939\,
            ce => 'H',
            sr => \N__20368\
        );

    \phase_controller_inst1.state_4_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__13057\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12285\,
            lcout => \phase_controller_inst1.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20939\,
            ce => 'H',
            sr => \N__20368\
        );

    \phase_controller_inst1.start_timer_hc_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010111010"
        )
    port map (
            in0 => \N__13193\,
            in1 => \N__12284\,
            in2 => \N__11888\,
            in3 => \N__11777\,
            lcout => \phase_controller_inst1.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20939\,
            ce => 'H',
            sr => \N__20368\
        );

    \phase_controller_inst1.state_RNI7NN7_0_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12379\,
            in2 => \_gnd_net_\,
            in3 => \N__12358\,
            lcout => \phase_controller_inst1.N_107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_RNO_0_3_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13058\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12277\,
            lcout => \phase_controller_inst1.N_110\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_RNO_0_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12339\,
            in2 => \_gnd_net_\,
            in3 => \N__12322\,
            lcout => \phase_controller_inst1.N_112\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_0_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010001000100"
        )
    port map (
            in0 => \N__12380\,
            in1 => \N__12359\,
            in2 => \N__19915\,
            in3 => \N__13160\,
            lcout => \phase_controller_inst1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20935\,
            ce => 'H',
            sr => \N__20373\
        );

    \phase_controller_inst1.T01_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010111010"
        )
    port map (
            in0 => \N__12346\,
            in1 => \N__13138\,
            in2 => \N__13016\,
            in3 => \N__12286\,
            lcout => shift_flag_start,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20935\,
            ce => 'H',
            sr => \N__20373\
        );

    \phase_controller_inst1.state_1_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__12347\,
            in1 => \N__12321\,
            in2 => \N__19914\,
            in3 => \N__13159\,
            lcout => \phase_controller_inst1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20935\,
            ce => 'H',
            sr => \N__20373\
        );

    \phase_controller_inst1.start_timer_tr_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001110"
        )
    port map (
            in0 => \N__12127\,
            in1 => \N__13139\,
            in2 => \N__12290\,
            in3 => \N__12256\,
            lcout => \phase_controller_inst1.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20935\,
            ce => 'H',
            sr => \N__20373\
        );

    \phase_controller_slave.stoper_tr.target_time_4_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__14824\,
            in1 => \N__17068\,
            in2 => \_gnd_net_\,
            in3 => \N__14722\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20930\,
            ce => \N__12671\,
            sr => \N__20378\
        );

    \phase_controller_slave.stoper_tr.target_time_5_LC_5_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__14723\,
            in1 => \N__14825\,
            in2 => \_gnd_net_\,
            in3 => \N__16927\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20930\,
            ce => \N__12671\,
            sr => \N__20378\
        );

    \phase_controller_slave.stoper_tr.target_time_1_LC_5_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__14823\,
            in1 => \N__14721\,
            in2 => \N__16483\,
            in3 => \N__14888\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20930\,
            ce => \N__12671\,
            sr => \N__20378\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__14433\,
            in1 => \N__12089\,
            in2 => \N__12080\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_5_17_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_5_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12071\,
            in2 => \N__12059\,
            in3 => \N__14398\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12497\,
            in2 => \N__12491\,
            in3 => \N__14368\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__14320\,
            in1 => \N__12482\,
            in2 => \N__12476\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_5_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12467\,
            in2 => \N__12461\,
            in3 => \N__14287\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12452\,
            in2 => \N__12446\,
            in3 => \N__14254\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12437\,
            in2 => \N__12428\,
            in3 => \N__14225\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_5_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12419\,
            in2 => \N__12413\,
            in3 => \N__14651\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_5_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12404\,
            in2 => \N__12398\,
            in3 => \N__14621\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_5_18_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12599\,
            in2 => \N__12389\,
            in3 => \N__14597\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12584\,
            in2 => \N__12575\,
            in3 => \N__14570\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_5_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12566\,
            in2 => \N__12560\,
            in3 => \N__14546\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12695\,
            in2 => \N__12551\,
            in3 => \N__14516\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__14492\,
            in1 => \N__12755\,
            in2 => \N__12542\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_5_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__14465\,
            in1 => \N__12746\,
            in2 => \N__12533\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_5_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12608\,
            in2 => \N__12524\,
            in3 => \N__14987\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12677\,
            in2 => \N__12515\,
            in3 => \N__14960\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_5_19_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12686\,
            in2 => \N__12506\,
            in3 => \N__14936\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12590\,
            in2 => \N__12632\,
            in3 => \N__14912\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_5_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12623\,
            lcout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_5_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12620\,
            in3 => \N__14846\,
            lcout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__14848\,
            in1 => \N__15168\,
            in2 => \_gnd_net_\,
            in3 => \N__14441\,
            lcout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_9_LC_5_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__14745\,
            in1 => \N__16994\,
            in2 => \_gnd_net_\,
            in3 => \N__17031\,
            lcout => \phase_controller_inst1.stoper_tr.N_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_5_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__14847\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15167\,
            lcout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.target_time_16_LC_5_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16711\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20907\,
            ce => \N__12667\,
            sr => \N__20399\
        );

    \phase_controller_slave.stoper_tr.target_time_10_LC_5_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__12721\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16588\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20907\,
            ce => \N__12667\,
            sr => \N__20399\
        );

    \phase_controller_slave.stoper_tr.target_time_19_LC_5_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18547\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20907\,
            ce => \N__12667\,
            sr => \N__20399\
        );

    \phase_controller_slave.stoper_tr.target_time_14_LC_5_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__14756\,
            in1 => \N__16996\,
            in2 => \_gnd_net_\,
            in3 => \N__17038\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20907\,
            ce => \N__12667\,
            sr => \N__20399\
        );

    \phase_controller_slave.stoper_tr.target_time_15_LC_5_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__16995\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14757\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20907\,
            ce => \N__12667\,
            sr => \N__20399\
        );

    \phase_controller_slave.stoper_tr.target_time_13_LC_5_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__12722\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16618\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20907\,
            ce => \N__12667\,
            sr => \N__20399\
        );

    \phase_controller_slave.stoper_tr.target_time_18_LC_5_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16792\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20907\,
            ce => \N__12667\,
            sr => \N__20399\
        );

    \phase_controller_slave.stoper_tr.target_time_17_LC_5_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16750\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20907\,
            ce => \N__12667\,
            sr => \N__20399\
        );

    \phase_controller_slave.stoper_tr.time_passed_LC_5_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__13126\,
            in1 => \N__14852\,
            in2 => \N__13445\,
            in3 => \N__15177\,
            lcout => \phase_controller_slave.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20903\,
            ce => 'H',
            sr => \N__20407\
        );

    \phase_controller_slave.state_4_LC_5_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010111011101110"
        )
    port map (
            in0 => \N__13094\,
            in1 => \N__12927\,
            in2 => \N__13083\,
            in3 => \N__13015\,
            lcout => \phase_controller_slave.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20899\,
            ce => 'H',
            sr => \N__20411\
        );

    \phase_controller_slave.start_timer_tr_LC_5_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101110"
        )
    port map (
            in0 => \N__12638\,
            in1 => \N__15235\,
            in2 => \N__12936\,
            in3 => \N__13093\,
            lcout => \phase_controller_slave.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20899\,
            ce => 'H',
            sr => \N__20411\
        );

    \phase_controller_slave.state_0_LC_5_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__13417\,
            in1 => \N__13125\,
            in2 => \N__15707\,
            in3 => \N__13106\,
            lcout => \phase_controller_slave.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20899\,
            ce => 'H',
            sr => \N__20411\
        );

    \phase_controller_slave.start_timer_tr_RNO_0_LC_5_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15699\,
            in2 => \_gnd_net_\,
            in3 => \N__13416\,
            lcout => \phase_controller_slave.start_timer_tr_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.state_RNIVDE2_0_LC_5_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13127\,
            in2 => \_gnd_net_\,
            in3 => \N__13105\,
            lcout => \phase_controller_slave.state_RNIVDE2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.state_RNO_0_3_LC_5_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13071\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13014\,
            lcout => \phase_controller_slave.state_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MAX_D2_LC_5_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12977\,
            lcout => \il_max_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20888\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.start_timer_hc_RNO_1_LC_5_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17264\,
            in2 => \_gnd_net_\,
            in3 => \N__12960\,
            lcout => \phase_controller_slave.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MAX_D1_LC_5_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12992\,
            lcout => \il_max_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20888\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.state_1_LC_5_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001100"
        )
    port map (
            in0 => \N__13288\,
            in1 => \N__15695\,
            in2 => \N__13421\,
            in3 => \N__13306\,
            lcout => \phase_controller_slave.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20882\,
            ce => 'H',
            sr => \N__20418\
        );

    \phase_controller_slave.state_3_LC_5_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000010101100"
        )
    port map (
            in0 => \N__12971\,
            in1 => \N__17265\,
            in2 => \N__12941\,
            in3 => \N__12961\,
            lcout => \phase_controller_slave.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20882\,
            ce => 'H',
            sr => \N__20418\
        );

    \phase_controller_slave.state_2_LC_5_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__17266\,
            in1 => \N__13289\,
            in2 => \N__13307\,
            in3 => \N__12962\,
            lcout => \phase_controller_slave.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20882\,
            ce => 'H',
            sr => \N__20418\
        );

    \phase_controller_slave.start_timer_hc_LC_5_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001110"
        )
    port map (
            in0 => \N__12799\,
            in1 => \N__12947\,
            in2 => \N__13262\,
            in3 => \N__12940\,
            lcout => \phase_controller_slave.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20882\,
            ce => 'H',
            sr => \N__20418\
        );

    \phase_controller_slave.start_timer_hc_RNO_0_LC_5_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13302\,
            in2 => \_gnd_net_\,
            in3 => \N__13282\,
            lcout => \phase_controller_slave.start_timer_hc_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D1_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13250\,
            lcout => \il_max_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20937\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MIN_D1_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13235\,
            lcout => \il_min_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20937\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D2_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13223\,
            lcout => \il_max_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20937\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_RNO_1_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16889\,
            in2 => \_gnd_net_\,
            in3 => \N__13204\,
            lcout => \phase_controller_inst1.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D2_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13166\,
            lcout => \il_min_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20931\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D1_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13184\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_min_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20931\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_RNIR0JF_1_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19910\,
            in2 => \_gnd_net_\,
            in3 => \N__13150\,
            lcout => \phase_controller_inst1.T01_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_8_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__15147\,
            in1 => \N__15330\,
            in2 => \N__14633\,
            in3 => \N__15459\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20914\,
            ce => 'H',
            sr => \N__20374\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_7_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__15458\,
            in1 => \N__15148\,
            in2 => \N__15346\,
            in3 => \N__14210\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20914\,
            ce => 'H',
            sr => \N__20374\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_16_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__15453\,
            in1 => \N__15135\,
            in2 => \N__15336\,
            in3 => \N__14969\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20908\,
            ce => 'H',
            sr => \N__20379\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_12_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__15130\,
            in1 => \N__15304\,
            in2 => \N__14528\,
            in3 => \N__15456\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20908\,
            ce => 'H',
            sr => \N__20379\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_15_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__15452\,
            in1 => \N__15134\,
            in2 => \N__15335\,
            in3 => \N__14450\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20908\,
            ce => 'H',
            sr => \N__20379\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_14_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__15132\,
            in1 => \N__15306\,
            in2 => \N__14477\,
            in3 => \N__15457\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20908\,
            ce => 'H',
            sr => \N__20379\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_11_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__15451\,
            in1 => \N__15133\,
            in2 => \N__15334\,
            in3 => \N__14555\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20908\,
            ce => 'H',
            sr => \N__20379\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_13_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__15131\,
            in1 => \N__15305\,
            in2 => \N__15478\,
            in3 => \N__14501\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20908\,
            ce => 'H',
            sr => \N__20379\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_9_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__15454\,
            in1 => \N__15136\,
            in2 => \N__15337\,
            in3 => \N__14606\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20908\,
            ce => 'H',
            sr => \N__20379\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_10_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__15129\,
            in1 => \N__15303\,
            in2 => \N__14582\,
            in3 => \N__15455\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20908\,
            ce => 'H',
            sr => \N__20379\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_19_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__15105\,
            in1 => \N__15434\,
            in2 => \N__15344\,
            in3 => \N__14894\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20904\,
            ce => 'H',
            sr => \N__20384\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_17_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__15104\,
            in1 => \N__15433\,
            in2 => \N__15343\,
            in3 => \N__14945\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20904\,
            ce => 'H',
            sr => \N__20384\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_18_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__15432\,
            in1 => \N__15320\,
            in2 => \N__15149\,
            in3 => \N__14921\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20904\,
            ce => 'H',
            sr => \N__20384\
        );

    \phase_controller_slave.stoper_tr.stoper_state_1_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000001100100"
        )
    port map (
            in0 => \N__15435\,
            in1 => \N__15107\,
            in2 => \N__15345\,
            in3 => \N__15184\,
            lcout => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20900\,
            ce => \N__20190\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGUTL_6_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18845\,
            in2 => \_gnd_net_\,
            in3 => \N__18326\,
            lcout => \delay_measurement_inst.delay_hc_reg_3_0_a2_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__15285\,
            in1 => \N__15420\,
            in2 => \_gnd_net_\,
            in3 => \N__15103\,
            lcout => \phase_controller_slave.stoper_tr.time_passed_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_4_LC_7_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18373\,
            in2 => \_gnd_net_\,
            in3 => \N__18415\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_232_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MIN_D2_LC_7_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13430\,
            lcout => \il_min_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20896\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_esr_5_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__15831\,
            in1 => \N__13670\,
            in2 => \N__15539\,
            in3 => \N__18377\,
            lcout => measured_delay_hc_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20889\,
            ce => \N__15740\,
            sr => \N__20400\
        );

    \delay_measurement_inst.delay_hc_reg_esr_2_LC_7_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__15002\,
            in1 => \N__15532\,
            in2 => \N__13673\,
            in3 => \N__15829\,
            lcout => measured_delay_hc_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20889\,
            ce => \N__15740\,
            sr => \N__20400\
        );

    \delay_measurement_inst.delay_hc_reg_esr_11_LC_7_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__15802\,
            in1 => \N__19569\,
            in2 => \_gnd_net_\,
            in3 => \N__19046\,
            lcout => measured_delay_hc_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20889\,
            ce => \N__15740\,
            sr => \N__20400\
        );

    \delay_measurement_inst.delay_hc_reg_esr_12_LC_7_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__19568\,
            in1 => \N__15803\,
            in2 => \_gnd_net_\,
            in3 => \N__19007\,
            lcout => measured_delay_hc_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20889\,
            ce => \N__15740\,
            sr => \N__20400\
        );

    \delay_measurement_inst.delay_hc_reg_ess_3_LC_7_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__15833\,
            in1 => \N__15538\,
            in2 => \N__18467\,
            in3 => \N__13672\,
            lcout => measured_delay_hc_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20889\,
            ce => \N__15740\,
            sr => \N__20400\
        );

    \delay_measurement_inst.delay_hc_reg_esr_4_LC_7_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__13669\,
            in1 => \N__15533\,
            in2 => \N__18425\,
            in3 => \N__15830\,
            lcout => measured_delay_hc_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20889\,
            ce => \N__15740\,
            sr => \N__20400\
        );

    \delay_measurement_inst.delay_hc_reg_ess_1_LC_7_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111000010000000"
        )
    port map (
            in0 => \N__15832\,
            in1 => \N__13671\,
            in2 => \N__15035\,
            in3 => \N__15537\,
            lcout => measured_delay_hc_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20889\,
            ce => \N__15740\,
            sr => \N__20400\
        );

    \delay_measurement_inst.delay_hc_reg_esr_10_LC_7_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__19567\,
            in1 => \N__15801\,
            in2 => \_gnd_net_\,
            in3 => \N__19085\,
            lcout => measured_delay_hc_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20889\,
            ce => \N__15740\,
            sr => \N__20400\
        );

    \delay_measurement_inst.delay_hc_reg_esr_9_LC_7_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000110001"
        )
    port map (
            in0 => \N__19558\,
            in1 => \N__15548\,
            in2 => \N__19154\,
            in3 => \N__15800\,
            lcout => measured_delay_hc_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20883\,
            ce => \N__15732\,
            sr => \N__20408\
        );

    \delay_measurement_inst.delay_hc_reg_esr_15_LC_7_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011001000"
        )
    port map (
            in0 => \N__15500\,
            in1 => \N__18853\,
            in2 => \N__19571\,
            in3 => \N__19829\,
            lcout => measured_delay_hc_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20883\,
            ce => \N__15732\,
            sr => \N__20408\
        );

    \delay_measurement_inst.delay_hc_reg_esr_19_LC_7_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__19826\,
            in1 => \N__19562\,
            in2 => \_gnd_net_\,
            in3 => \N__19309\,
            lcout => measured_delay_hc_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20883\,
            ce => \N__15732\,
            sr => \N__20408\
        );

    \delay_measurement_inst.delay_hc_reg_esr_6_LC_7_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010011110101"
        )
    port map (
            in0 => \N__15529\,
            in1 => \N__18854\,
            in2 => \N__18335\,
            in3 => \N__15828\,
            lcout => measured_delay_hc_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20883\,
            ce => \N__15732\,
            sr => \N__20408\
        );

    \delay_measurement_inst.delay_hc_reg_esr_17_LC_7_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__19825\,
            in1 => \N__19561\,
            in2 => \_gnd_net_\,
            in3 => \N__19408\,
            lcout => measured_delay_hc_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20883\,
            ce => \N__15732\,
            sr => \N__20408\
        );

    \delay_measurement_inst.delay_hc_reg_esr_16_LC_7_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__19559\,
            in1 => \N__19459\,
            in2 => \_gnd_net_\,
            in3 => \N__19827\,
            lcout => measured_delay_hc_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20883\,
            ce => \N__15732\,
            sr => \N__20408\
        );

    \delay_measurement_inst.delay_hc_reg_esr_14_LC_7_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__19557\,
            in1 => \N__15799\,
            in2 => \_gnd_net_\,
            in3 => \N__18916\,
            lcout => measured_delay_hc_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20883\,
            ce => \N__15732\,
            sr => \N__20408\
        );

    \delay_measurement_inst.delay_hc_reg_esr_18_LC_7_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__19560\,
            in1 => \N__19355\,
            in2 => \_gnd_net_\,
            in3 => \N__19828\,
            lcout => measured_delay_hc_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20883\,
            ce => \N__15732\,
            sr => \N__20408\
        );

    \delay_measurement_inst.delay_hc_reg_7_LC_7_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__13871\,
            in1 => \N__15530\,
            in2 => \N__18281\,
            in3 => \N__15559\,
            lcout => measured_delay_hc_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20876\,
            ce => 'H',
            sr => \N__20412\
        );

    \delay_measurement_inst.delay_hc_reg_8_LC_7_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__13838\,
            in1 => \N__15531\,
            in2 => \N__18236\,
            in3 => \N__15560\,
            lcout => measured_delay_hc_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20876\,
            ce => 'H',
            sr => \N__20412\
        );

    \delay_measurement_inst.delay_tr_timer.counter_0_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17559\,
            in1 => \N__17232\,
            in2 => \_gnd_net_\,
            in3 => \N__13808\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_13_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            clk => \N__20932\,
            ce => \N__14171\,
            sr => \N__20353\
        );

    \delay_measurement_inst.delay_tr_timer.counter_1_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17554\,
            in1 => \N__17211\,
            in2 => \_gnd_net_\,
            in3 => \N__13805\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            clk => \N__20932\,
            ce => \N__14171\,
            sr => \N__20353\
        );

    \delay_measurement_inst.delay_tr_timer.counter_2_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17560\,
            in1 => \N__15657\,
            in2 => \_gnd_net_\,
            in3 => \N__14126\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            clk => \N__20932\,
            ce => \N__14171\,
            sr => \N__20353\
        );

    \delay_measurement_inst.delay_tr_timer.counter_3_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17555\,
            in1 => \N__15633\,
            in2 => \_gnd_net_\,
            in3 => \N__14123\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            clk => \N__20932\,
            ce => \N__14171\,
            sr => \N__20353\
        );

    \delay_measurement_inst.delay_tr_timer.counter_4_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17561\,
            in1 => \N__15611\,
            in2 => \_gnd_net_\,
            in3 => \N__14120\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            clk => \N__20932\,
            ce => \N__14171\,
            sr => \N__20353\
        );

    \delay_measurement_inst.delay_tr_timer.counter_5_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17556\,
            in1 => \N__16037\,
            in2 => \_gnd_net_\,
            in3 => \N__14117\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            clk => \N__20932\,
            ce => \N__14171\,
            sr => \N__20353\
        );

    \delay_measurement_inst.delay_tr_timer.counter_6_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17558\,
            in1 => \N__16017\,
            in2 => \_gnd_net_\,
            in3 => \N__14114\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            clk => \N__20932\,
            ce => \N__14171\,
            sr => \N__20353\
        );

    \delay_measurement_inst.delay_tr_timer.counter_7_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17557\,
            in1 => \N__15993\,
            in2 => \_gnd_net_\,
            in3 => \N__14111\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            clk => \N__20932\,
            ce => \N__14171\,
            sr => \N__20353\
        );

    \delay_measurement_inst.delay_tr_timer.counter_8_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17532\,
            in1 => \N__15970\,
            in2 => \_gnd_net_\,
            in3 => \N__14108\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_14_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            clk => \N__20925\,
            ce => \N__14172\,
            sr => \N__20355\
        );

    \delay_measurement_inst.delay_tr_timer.counter_9_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17567\,
            in1 => \N__15949\,
            in2 => \_gnd_net_\,
            in3 => \N__14105\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            clk => \N__20925\,
            ce => \N__14172\,
            sr => \N__20355\
        );

    \delay_measurement_inst.delay_tr_timer.counter_10_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17529\,
            in1 => \N__15927\,
            in2 => \_gnd_net_\,
            in3 => \N__14102\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            clk => \N__20925\,
            ce => \N__14172\,
            sr => \N__20355\
        );

    \delay_measurement_inst.delay_tr_timer.counter_11_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17564\,
            in1 => \N__15903\,
            in2 => \_gnd_net_\,
            in3 => \N__14156\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            clk => \N__20925\,
            ce => \N__14172\,
            sr => \N__20355\
        );

    \delay_measurement_inst.delay_tr_timer.counter_12_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17530\,
            in1 => \N__15881\,
            in2 => \_gnd_net_\,
            in3 => \N__14153\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            clk => \N__20925\,
            ce => \N__14172\,
            sr => \N__20355\
        );

    \delay_measurement_inst.delay_tr_timer.counter_13_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17565\,
            in1 => \N__15863\,
            in2 => \_gnd_net_\,
            in3 => \N__14150\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            clk => \N__20925\,
            ce => \N__14172\,
            sr => \N__20355\
        );

    \delay_measurement_inst.delay_tr_timer.counter_14_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17531\,
            in1 => \N__16209\,
            in2 => \_gnd_net_\,
            in3 => \N__14147\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            clk => \N__20925\,
            ce => \N__14172\,
            sr => \N__20355\
        );

    \delay_measurement_inst.delay_tr_timer.counter_15_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17566\,
            in1 => \N__16185\,
            in2 => \_gnd_net_\,
            in3 => \N__14144\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            clk => \N__20925\,
            ce => \N__14172\,
            sr => \N__20355\
        );

    \delay_measurement_inst.delay_tr_timer.counter_16_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17542\,
            in1 => \N__16162\,
            in2 => \_gnd_net_\,
            in3 => \N__14141\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_8_15_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            clk => \N__20921\,
            ce => \N__14173\,
            sr => \N__20361\
        );

    \delay_measurement_inst.delay_tr_timer.counter_17_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17546\,
            in1 => \N__16141\,
            in2 => \_gnd_net_\,
            in3 => \N__14138\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            clk => \N__20921\,
            ce => \N__14173\,
            sr => \N__20361\
        );

    \delay_measurement_inst.delay_tr_timer.counter_18_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17543\,
            in1 => \N__16119\,
            in2 => \_gnd_net_\,
            in3 => \N__14135\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            clk => \N__20921\,
            ce => \N__14173\,
            sr => \N__20361\
        );

    \delay_measurement_inst.delay_tr_timer.counter_19_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17547\,
            in1 => \N__16095\,
            in2 => \_gnd_net_\,
            in3 => \N__14132\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            clk => \N__20921\,
            ce => \N__14173\,
            sr => \N__20361\
        );

    \delay_measurement_inst.delay_tr_timer.counter_20_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17544\,
            in1 => \N__16073\,
            in2 => \_gnd_net_\,
            in3 => \N__14129\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            clk => \N__20921\,
            ce => \N__14173\,
            sr => \N__20361\
        );

    \delay_measurement_inst.delay_tr_timer.counter_21_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17548\,
            in1 => \N__16055\,
            in2 => \_gnd_net_\,
            in3 => \N__14201\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            clk => \N__20921\,
            ce => \N__14173\,
            sr => \N__20361\
        );

    \delay_measurement_inst.delay_tr_timer.counter_22_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17545\,
            in1 => \N__16374\,
            in2 => \_gnd_net_\,
            in3 => \N__14198\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            clk => \N__20921\,
            ce => \N__14173\,
            sr => \N__20361\
        );

    \delay_measurement_inst.delay_tr_timer.counter_23_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17549\,
            in1 => \N__16350\,
            in2 => \_gnd_net_\,
            in3 => \N__14195\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            clk => \N__20921\,
            ce => \N__14173\,
            sr => \N__20361\
        );

    \delay_measurement_inst.delay_tr_timer.counter_24_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17550\,
            in1 => \N__16327\,
            in2 => \_gnd_net_\,
            in3 => \N__14192\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_8_16_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            clk => \N__20915\,
            ce => \N__14174\,
            sr => \N__20369\
        );

    \delay_measurement_inst.delay_tr_timer.counter_25_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17562\,
            in1 => \N__16306\,
            in2 => \_gnd_net_\,
            in3 => \N__14189\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            clk => \N__20915\,
            ce => \N__14174\,
            sr => \N__20369\
        );

    \delay_measurement_inst.delay_tr_timer.counter_26_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17551\,
            in1 => \N__16272\,
            in2 => \_gnd_net_\,
            in3 => \N__14186\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            clk => \N__20915\,
            ce => \N__14174\,
            sr => \N__20369\
        );

    \delay_measurement_inst.delay_tr_timer.counter_27_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17563\,
            in1 => \N__16236\,
            in2 => \_gnd_net_\,
            in3 => \N__14183\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            clk => \N__20915\,
            ce => \N__14174\,
            sr => \N__20369\
        );

    \delay_measurement_inst.delay_tr_timer.counter_28_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17552\,
            in1 => \N__16286\,
            in2 => \_gnd_net_\,
            in3 => \N__14180\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_28\,
            clk => \N__20915\,
            ce => \N__14174\,
            sr => \N__20369\
        );

    \delay_measurement_inst.delay_tr_timer.counter_29_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__16250\,
            in1 => \N__17553\,
            in2 => \_gnd_net_\,
            in3 => \N__14177\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20915\,
            ce => \N__14174\,
            sr => \N__20369\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14440\,
            in2 => \N__14417\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_17_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_8_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14402\,
            in2 => \_gnd_net_\,
            in3 => \N__14375\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14372\,
            in2 => \N__14357\,
            in3 => \N__14330\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14327\,
            in3 => \N__14297\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14294\,
            in3 => \N__14261\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14258\,
            in2 => \_gnd_net_\,
            in3 => \N__14228\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14224\,
            in2 => \_gnd_net_\,
            in3 => \N__14204\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14650\,
            in2 => \_gnd_net_\,
            in3 => \N__14624\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14620\,
            in2 => \_gnd_net_\,
            in3 => \N__14600\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9\,
            ltout => OPEN,
            carryin => \bfn_8_18_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14596\,
            in2 => \_gnd_net_\,
            in3 => \N__14573\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14569\,
            in2 => \_gnd_net_\,
            in3 => \N__14549\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_8_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14542\,
            in2 => \_gnd_net_\,
            in3 => \N__14519\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14515\,
            in2 => \_gnd_net_\,
            in3 => \N__14495\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14491\,
            in2 => \_gnd_net_\,
            in3 => \N__14468\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_8_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14464\,
            in2 => \_gnd_net_\,
            in3 => \N__14444\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_8_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14983\,
            in2 => \_gnd_net_\,
            in3 => \N__14963\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14959\,
            in2 => \_gnd_net_\,
            in3 => \N__14939\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17\,
            ltout => OPEN,
            carryin => \bfn_8_19_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14935\,
            in2 => \_gnd_net_\,
            in3 => \N__14915\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14911\,
            in2 => \_gnd_net_\,
            in3 => \N__14897\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a3_1_LC_8_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__16401\,
            in1 => \N__16449\,
            in2 => \_gnd_net_\,
            in3 => \N__17085\,
            lcout => \phase_controller_inst1.stoper_tr.N_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15398\,
            in2 => \_gnd_net_\,
            in3 => \N__15074\,
            lcout => \phase_controller_slave.stoper_tr.time_passed11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0_6_LC_8_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__16548\,
            in1 => \N__16964\,
            in2 => \_gnd_net_\,
            in3 => \N__17111\,
            lcout => \phase_controller_inst1.stoper_tr.N_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_i_o2_15_LC_8_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__16698\,
            in1 => \N__16778\,
            in2 => \N__18546\,
            in3 => \N__16737\,
            lcout => \phase_controller_inst1.stoper_tr.N_32\,
            ltout => \phase_controller_inst1.stoper_tr.N_32_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_6_LC_8_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110001"
        )
    port map (
            in0 => \N__17022\,
            in1 => \N__16965\,
            in2 => \N__14726\,
            in3 => \N__16493\,
            lcout => \phase_controller_inst1.stoper_tr.N_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.stoper_state_0_LC_8_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__15436\,
            in1 => \N__15106\,
            in2 => \N__15347\,
            in3 => \N__15185\,
            lcout => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20897\,
            ce => \N__20189\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_8_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18443\,
            lcout => \delay_measurement_inst.elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20890\,
            ce => \N__19496\,
            sr => \N__20392\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_8_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18485\,
            lcout => \delay_measurement_inst.elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20890\,
            ce => \N__19496\,
            sr => \N__20392\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNID3EH4_1_LC_8_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__15008\,
            in1 => \N__15498\,
            in2 => \N__15017\,
            in3 => \N__15590\,
            lcout => \delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_8_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19003\,
            in1 => \N__19045\,
            in2 => \N__18964\,
            in3 => \N__19084\,
            lcout => \delay_measurement_inst.N_243\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_6_LC_8_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19145\,
            in2 => \_gnd_net_\,
            in3 => \N__18331\,
            lcout => \delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3GIH1_1_LC_8_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__18910\,
            in1 => \N__18462\,
            in2 => \N__15034\,
            in3 => \N__15001\,
            lcout => \delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3HO31_6_LC_8_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__18837\,
            in1 => \N__19144\,
            in2 => \_gnd_net_\,
            in3 => \N__18330\,
            lcout => \delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0TRB1_18_LC_8_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__19347\,
            in1 => \N__18463\,
            in2 => \N__19310\,
            in3 => \N__15000\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0QNN2_16_LC_8_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__19404\,
            in1 => \N__19460\,
            in2 => \N__15593\,
            in3 => \N__15589\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2PJ34_14_LC_8_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__15581\,
            in1 => \N__18911\,
            in2 => \N__15575\,
            in3 => \N__18838\,
            lcout => \delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4ESID_31_LC_8_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001111"
        )
    port map (
            in0 => \N__15572\,
            in1 => \N__15566\,
            in2 => \N__19570\,
            in3 => \N__15827\,
            lcout => \delay_measurement_inst.un3_elapsed_time_hc_0_i\,
            ltout => \delay_measurement_inst.un3_elapsed_time_hc_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBNQQD_31_LC_8_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15551\,
            in3 => \N__20463\,
            lcout => \delay_measurement_inst.un3_elapsed_time_hc_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_esr_RNO_0_9_LC_8_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__19824\,
            in1 => \N__15845\,
            in2 => \N__19153\,
            in3 => \N__18851\,
            lcout => \delay_measurement_inst.N_219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4TEU1_14_LC_8_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100100011"
        )
    port map (
            in0 => \N__15844\,
            in1 => \N__18839\,
            in2 => \N__18917\,
            in3 => \N__19146\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.N_237_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE5L06_31_LC_8_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111011100"
        )
    port map (
            in0 => \N__19823\,
            in1 => \N__19566\,
            in2 => \N__15542\,
            in3 => \N__15499\,
            lcout => \delay_measurement_inst.N_209\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_8_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__19458\,
            in1 => \N__19308\,
            in2 => \N__19409\,
            in3 => \N__19354\,
            lcout => \delay_measurement_inst.N_207\,
            ltout => \delay_measurement_inst.N_207_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBM7A4_14_LC_8_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010001"
        )
    port map (
            in0 => \N__19822\,
            in1 => \N__18852\,
            in2 => \N__15482\,
            in3 => \N__18915\,
            lcout => \delay_measurement_inst.N_216_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN2LL4_7_LC_8_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__15843\,
            in1 => \N__18277\,
            in2 => \N__18235\,
            in3 => \N__19821\,
            lcout => \delay_measurement_inst.N_247\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_esr_13_LC_8_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__19553\,
            in1 => \N__15798\,
            in2 => \_gnd_net_\,
            in3 => \N__18965\,
            lcout => measured_delay_hc_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20871\,
            ce => \N__15739\,
            sr => \N__20409\
        );

    \phase_controller_slave.S2_LC_8_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15706\,
            lcout => s4_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20866\,
            ce => 'H',
            sr => \N__20414\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17233\,
            in2 => \N__15658\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.elapsed_time_tr_3\,
            ltout => OPEN,
            carryin => \bfn_9_13_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__20926\,
            ce => \N__17194\,
            sr => \N__20352\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17212\,
            in2 => \N__15634\,
            in3 => \N__15662\,
            lcout => \delay_measurement_inst.elapsed_time_tr_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__20926\,
            ce => \N__17194\,
            sr => \N__20352\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15609\,
            in2 => \N__15659\,
            in3 => \N__15638\,
            lcout => \delay_measurement_inst.elapsed_time_tr_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__20926\,
            ce => \N__17194\,
            sr => \N__20352\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16035\,
            in2 => \N__15635\,
            in3 => \N__15614\,
            lcout => \delay_measurement_inst.delay_tr_reg3lto6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__20926\,
            ce => \N__17194\,
            sr => \N__20352\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15610\,
            in2 => \N__16018\,
            in3 => \N__15596\,
            lcout => \delay_measurement_inst.elapsed_time_tr_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__20926\,
            ce => \N__17194\,
            sr => \N__20352\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16036\,
            in2 => \N__15994\,
            in3 => \N__16022\,
            lcout => \delay_measurement_inst.elapsed_time_tr_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__20926\,
            ce => \N__17194\,
            sr => \N__20352\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15969\,
            in2 => \N__16019\,
            in3 => \N__15998\,
            lcout => \delay_measurement_inst.delay_tr_reg3lto9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__20926\,
            ce => \N__17194\,
            sr => \N__20352\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15948\,
            in2 => \N__15995\,
            in3 => \N__15974\,
            lcout => \delay_measurement_inst.elapsed_time_tr_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__20926\,
            ce => \N__17194\,
            sr => \N__20352\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15971\,
            in2 => \N__15928\,
            in3 => \N__15953\,
            lcout => \delay_measurement_inst.elapsed_time_tr_11\,
            ltout => OPEN,
            carryin => \bfn_9_14_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__20922\,
            ce => \N__17193\,
            sr => \N__20354\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15950\,
            in2 => \N__15904\,
            in3 => \N__15932\,
            lcout => \delay_measurement_inst.elapsed_time_tr_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__20922\,
            ce => \N__17193\,
            sr => \N__20354\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15879\,
            in2 => \N__15929\,
            in3 => \N__15908\,
            lcout => \delay_measurement_inst.elapsed_time_tr_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__20922\,
            ce => \N__17193\,
            sr => \N__20354\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15861\,
            in2 => \N__15905\,
            in3 => \N__15884\,
            lcout => \delay_measurement_inst.delay_tr_reg3lto14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__20922\,
            ce => \N__17193\,
            sr => \N__20354\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15880\,
            in2 => \N__16210\,
            in3 => \N__15866\,
            lcout => \delay_measurement_inst.delay_tr_reg3lto15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__20922\,
            ce => \N__17193\,
            sr => \N__20354\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15862\,
            in2 => \N__16186\,
            in3 => \N__15848\,
            lcout => \delay_measurement_inst.elapsed_time_tr_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__20922\,
            ce => \N__17193\,
            sr => \N__20354\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16161\,
            in2 => \N__16211\,
            in3 => \N__16190\,
            lcout => \delay_measurement_inst.elapsed_time_tr_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__20922\,
            ce => \N__17193\,
            sr => \N__20354\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16140\,
            in2 => \N__16187\,
            in3 => \N__16166\,
            lcout => \delay_measurement_inst.elapsed_time_tr_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__20922\,
            ce => \N__17193\,
            sr => \N__20354\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16163\,
            in2 => \N__16120\,
            in3 => \N__16145\,
            lcout => \delay_measurement_inst.elapsed_time_tr_19\,
            ltout => OPEN,
            carryin => \bfn_9_15_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__20916\,
            ce => \N__17192\,
            sr => \N__20356\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16142\,
            in2 => \N__16096\,
            in3 => \N__16124\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__20916\,
            ce => \N__17192\,
            sr => \N__20356\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16071\,
            in2 => \N__16121\,
            in3 => \N__16100\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__20916\,
            ce => \N__17192\,
            sr => \N__20356\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16053\,
            in2 => \N__16097\,
            in3 => \N__16076\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__20916\,
            ce => \N__17192\,
            sr => \N__20356\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16072\,
            in2 => \N__16375\,
            in3 => \N__16058\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__20916\,
            ce => \N__17192\,
            sr => \N__20356\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16054\,
            in2 => \N__16351\,
            in3 => \N__16040\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__20916\,
            ce => \N__17192\,
            sr => \N__20356\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16326\,
            in2 => \N__16376\,
            in3 => \N__16355\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__20916\,
            ce => \N__17192\,
            sr => \N__20356\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16305\,
            in2 => \N__16352\,
            in3 => \N__16331\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__20916\,
            ce => \N__17192\,
            sr => \N__20356\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16328\,
            in2 => \N__16273\,
            in3 => \N__16310\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\,
            ltout => OPEN,
            carryin => \bfn_9_16_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__20909\,
            ce => \N__17191\,
            sr => \N__20362\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16307\,
            in2 => \N__16237\,
            in3 => \N__16289\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__20909\,
            ce => \N__17191\,
            sr => \N__20362\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16285\,
            in2 => \N__16274\,
            in3 => \N__16253\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__20909\,
            ce => \N__17191\,
            sr => \N__20362\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16249\,
            in2 => \N__16238\,
            in3 => \N__16217\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__20909\,
            ce => \N__17191\,
            sr => \N__20362\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16214\,
            lcout => \delay_measurement_inst.elapsed_time_tr_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20909\,
            ce => \N__17191\,
            sr => \N__20362\
        );

    \delay_measurement_inst.delay_tr_reg_esr_15_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011001000"
        )
    port map (
            in0 => \N__18023\,
            in1 => \N__17941\,
            in2 => \N__18688\,
            in3 => \N__18579\,
            lcout => measured_delay_tr_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20905\,
            ce => \N__18501\,
            sr => \N__20370\
        );

    \delay_measurement_inst.delay_tr_reg_esr_9_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000100011"
        )
    port map (
            in0 => \N__18105\,
            in1 => \N__18203\,
            in2 => \N__18689\,
            in3 => \N__18147\,
            lcout => measured_delay_tr_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20905\,
            ce => \N__18501\,
            sr => \N__20370\
        );

    \delay_measurement_inst.delay_tr_reg_esr_4_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__18193\,
            in1 => \N__18775\,
            in2 => \N__17903\,
            in3 => \N__17417\,
            lcout => measured_delay_tr_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20905\,
            ce => \N__18501\,
            sr => \N__20370\
        );

    \delay_measurement_inst.delay_tr_reg_esr_5_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000010100000"
        )
    port map (
            in0 => \N__18776\,
            in1 => \N__18194\,
            in2 => \N__17438\,
            in3 => \N__17899\,
            lcout => measured_delay_tr_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20905\,
            ce => \N__18501\,
            sr => \N__20370\
        );

    \delay_measurement_inst.delay_tr_reg_esr_6_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011111101"
        )
    port map (
            in0 => \N__18195\,
            in1 => \N__17942\,
            in2 => \N__17981\,
            in3 => \N__18777\,
            lcout => measured_delay_tr_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20905\,
            ce => \N__18501\,
            sr => \N__20370\
        );

    \delay_measurement_inst.delay_tr_reg_ess_1_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110000010100000"
        )
    port map (
            in0 => \N__18778\,
            in1 => \N__18196\,
            in2 => \N__17375\,
            in3 => \N__17900\,
            lcout => measured_delay_tr_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20905\,
            ce => \N__18501\,
            sr => \N__20370\
        );

    \delay_measurement_inst.delay_tr_reg_esr_2_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__18192\,
            in1 => \N__18774\,
            in2 => \N__17902\,
            in3 => \N__17348\,
            lcout => measured_delay_tr_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20905\,
            ce => \N__18501\,
            sr => \N__20370\
        );

    \delay_measurement_inst.delay_tr_reg_ess_3_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110000010100000"
        )
    port map (
            in0 => \N__18779\,
            in1 => \N__18197\,
            in2 => \N__17402\,
            in3 => \N__17901\,
            lcout => measured_delay_tr_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20905\,
            ce => \N__18501\,
            sr => \N__20370\
        );

    \delay_measurement_inst.delay_tr_reg_esr_10_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__18676\,
            in1 => \N__18148\,
            in2 => \_gnd_net_\,
            in3 => \N__17654\,
            lcout => measured_delay_tr_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20901\,
            ce => \N__18505\,
            sr => \N__20372\
        );

    \delay_measurement_inst.delay_tr_reg_esr_12_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__18150\,
            in1 => \N__18678\,
            in2 => \_gnd_net_\,
            in3 => \N__17716\,
            lcout => measured_delay_tr_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20901\,
            ce => \N__18505\,
            sr => \N__20372\
        );

    \delay_measurement_inst.delay_tr_reg_esr_16_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__18681\,
            in1 => \N__17792\,
            in2 => \_gnd_net_\,
            in3 => \N__18591\,
            lcout => measured_delay_tr_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20901\,
            ce => \N__18505\,
            sr => \N__20372\
        );

    \delay_measurement_inst.delay_tr_reg_esr_14_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101011"
        )
    port map (
            in0 => \N__18059\,
            in1 => \N__18680\,
            in2 => \N__18155\,
            in3 => \_gnd_net_\,
            lcout => measured_delay_tr_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20901\,
            ce => \N__18505\,
            sr => \N__20372\
        );

    \delay_measurement_inst.delay_tr_reg_esr_17_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__17774\,
            in1 => \N__18683\,
            in2 => \_gnd_net_\,
            in3 => \N__18592\,
            lcout => measured_delay_tr_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20901\,
            ce => \N__18505\,
            sr => \N__20372\
        );

    \delay_measurement_inst.delay_tr_reg_esr_18_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__18593\,
            in1 => \N__18682\,
            in2 => \_gnd_net_\,
            in3 => \N__17750\,
            lcout => measured_delay_tr_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20901\,
            ce => \N__18505\,
            sr => \N__20372\
        );

    \delay_measurement_inst.delay_tr_reg_esr_11_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__18677\,
            in1 => \N__18149\,
            in2 => \_gnd_net_\,
            in3 => \N__17695\,
            lcout => measured_delay_tr_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20901\,
            ce => \N__18505\,
            sr => \N__20372\
        );

    \delay_measurement_inst.delay_tr_reg_esr_13_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__18151\,
            in1 => \N__18679\,
            in2 => \_gnd_net_\,
            in3 => \N__17675\,
            lcout => measured_delay_tr_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20901\,
            ce => \N__18505\,
            sr => \N__20372\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_6_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__16807\,
            in1 => \_gnd_net_\,
            in2 => \N__17850\,
            in3 => \N__18707\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_3_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16782\,
            in1 => \N__16736\,
            in2 => \N__18527\,
            in3 => \N__16697\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_6_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16665\,
            in1 => \N__16638\,
            in2 => \N__16611\,
            in3 => \N__16576\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_0_6\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_9_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__16515\,
            in1 => \_gnd_net_\,
            in2 => \N__16496\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_9\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16904\,
            in1 => \N__17120\,
            in2 => \N__17114\,
            in3 => \N__17110\,
            lcout => \phase_controller_inst1.stoper_tr.N_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4_3_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17061\,
            in1 => \N__17016\,
            in2 => \N__16963\,
            in3 => \N__16920\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.S1_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16898\,
            lcout => s1_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20891\,
            ce => 'H',
            sr => \N__20380\
        );

    \delay_measurement_inst.delay_hc_timer.counter_0_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20523\,
            in1 => \N__18483\,
            in2 => \_gnd_net_\,
            in3 => \N__16838\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_9_21_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            clk => \N__20884\,
            ce => \N__20651\,
            sr => \N__20385\
        );

    \delay_measurement_inst.delay_hc_timer.counter_1_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20582\,
            in1 => \N__18441\,
            in2 => \_gnd_net_\,
            in3 => \N__16835\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            clk => \N__20884\,
            ce => \N__20651\,
            sr => \N__20385\
        );

    \delay_measurement_inst.delay_hc_timer.counter_2_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20524\,
            in1 => \N__18396\,
            in2 => \_gnd_net_\,
            in3 => \N__16832\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            clk => \N__20884\,
            ce => \N__20651\,
            sr => \N__20385\
        );

    \delay_measurement_inst.delay_hc_timer.counter_3_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20583\,
            in1 => \N__18354\,
            in2 => \_gnd_net_\,
            in3 => \N__16829\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            clk => \N__20884\,
            ce => \N__20651\,
            sr => \N__20385\
        );

    \delay_measurement_inst.delay_hc_timer.counter_4_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20525\,
            in1 => \N__18296\,
            in2 => \_gnd_net_\,
            in3 => \N__16826\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            clk => \N__20884\,
            ce => \N__20651\,
            sr => \N__20385\
        );

    \delay_measurement_inst.delay_hc_timer.counter_5_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20584\,
            in1 => \N__18251\,
            in2 => \_gnd_net_\,
            in3 => \N__16823\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            clk => \N__20884\,
            ce => \N__20651\,
            sr => \N__20385\
        );

    \delay_measurement_inst.delay_hc_timer.counter_6_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20526\,
            in1 => \N__19173\,
            in2 => \_gnd_net_\,
            in3 => \N__17147\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            clk => \N__20884\,
            ce => \N__20651\,
            sr => \N__20385\
        );

    \delay_measurement_inst.delay_hc_timer.counter_7_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20585\,
            in1 => \N__19104\,
            in2 => \_gnd_net_\,
            in3 => \N__17144\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            clk => \N__20884\,
            ce => \N__20651\,
            sr => \N__20385\
        );

    \delay_measurement_inst.delay_hc_timer.counter_8_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20581\,
            in1 => \N__19063\,
            in2 => \_gnd_net_\,
            in3 => \N__17141\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_9_22_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            clk => \N__20877\,
            ce => \N__20659\,
            sr => \N__20393\
        );

    \delay_measurement_inst.delay_hc_timer.counter_9_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20593\,
            in1 => \N__19024\,
            in2 => \_gnd_net_\,
            in3 => \N__17138\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            clk => \N__20877\,
            ce => \N__20659\,
            sr => \N__20393\
        );

    \delay_measurement_inst.delay_hc_timer.counter_10_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20578\,
            in1 => \N__18984\,
            in2 => \_gnd_net_\,
            in3 => \N__17135\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            clk => \N__20877\,
            ce => \N__20659\,
            sr => \N__20393\
        );

    \delay_measurement_inst.delay_hc_timer.counter_11_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20590\,
            in1 => \N__18936\,
            in2 => \_gnd_net_\,
            in3 => \N__17132\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            clk => \N__20877\,
            ce => \N__20659\,
            sr => \N__20393\
        );

    \delay_measurement_inst.delay_hc_timer.counter_12_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20579\,
            in1 => \N__18869\,
            in2 => \_gnd_net_\,
            in3 => \N__17129\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            clk => \N__20877\,
            ce => \N__20659\,
            sr => \N__20393\
        );

    \delay_measurement_inst.delay_hc_timer.counter_13_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20591\,
            in1 => \N__19475\,
            in2 => \_gnd_net_\,
            in3 => \N__17126\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            clk => \N__20877\,
            ce => \N__20659\,
            sr => \N__20393\
        );

    \delay_measurement_inst.delay_hc_timer.counter_14_LC_9_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20580\,
            in1 => \N__19428\,
            in2 => \_gnd_net_\,
            in3 => \N__17123\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            clk => \N__20877\,
            ce => \N__20659\,
            sr => \N__20393\
        );

    \delay_measurement_inst.delay_hc_timer.counter_15_LC_9_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20592\,
            in1 => \N__19374\,
            in2 => \_gnd_net_\,
            in3 => \N__17174\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            clk => \N__20877\,
            ce => \N__20659\,
            sr => \N__20393\
        );

    \delay_measurement_inst.delay_hc_timer.counter_16_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20594\,
            in1 => \N__19327\,
            in2 => \_gnd_net_\,
            in3 => \N__17171\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_9_23_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            clk => \N__20872\,
            ce => \N__20658\,
            sr => \N__20397\
        );

    \delay_measurement_inst.delay_hc_timer.counter_17_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20586\,
            in1 => \N__19276\,
            in2 => \_gnd_net_\,
            in3 => \N__17168\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            clk => \N__20872\,
            ce => \N__20658\,
            sr => \N__20397\
        );

    \delay_measurement_inst.delay_hc_timer.counter_18_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20595\,
            in1 => \N__19254\,
            in2 => \_gnd_net_\,
            in3 => \N__17165\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            clk => \N__20872\,
            ce => \N__20658\,
            sr => \N__20397\
        );

    \delay_measurement_inst.delay_hc_timer.counter_19_LC_9_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20587\,
            in1 => \N__19230\,
            in2 => \_gnd_net_\,
            in3 => \N__17162\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            clk => \N__20872\,
            ce => \N__20658\,
            sr => \N__20397\
        );

    \delay_measurement_inst.delay_hc_timer.counter_20_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20596\,
            in1 => \N__19208\,
            in2 => \_gnd_net_\,
            in3 => \N__17159\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            clk => \N__20872\,
            ce => \N__20658\,
            sr => \N__20397\
        );

    \delay_measurement_inst.delay_hc_timer.counter_21_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20588\,
            in1 => \N__19190\,
            in2 => \_gnd_net_\,
            in3 => \N__17156\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            clk => \N__20872\,
            ce => \N__20658\,
            sr => \N__20397\
        );

    \delay_measurement_inst.delay_hc_timer.counter_22_LC_9_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20597\,
            in1 => \N__19734\,
            in2 => \_gnd_net_\,
            in3 => \N__17153\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            clk => \N__20872\,
            ce => \N__20658\,
            sr => \N__20397\
        );

    \delay_measurement_inst.delay_hc_timer.counter_23_LC_9_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20589\,
            in1 => \N__19710\,
            in2 => \_gnd_net_\,
            in3 => \N__17150\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            clk => \N__20872\,
            ce => \N__20658\,
            sr => \N__20397\
        );

    \delay_measurement_inst.delay_hc_timer.counter_24_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20527\,
            in1 => \N__19687\,
            in2 => \_gnd_net_\,
            in3 => \N__17294\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_9_24_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            clk => \N__20868\,
            ce => \N__20663\,
            sr => \N__20401\
        );

    \delay_measurement_inst.delay_hc_timer.counter_25_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20531\,
            in1 => \N__19666\,
            in2 => \_gnd_net_\,
            in3 => \N__17291\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            clk => \N__20868\,
            ce => \N__20663\,
            sr => \N__20401\
        );

    \delay_measurement_inst.delay_hc_timer.counter_26_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20528\,
            in1 => \N__19632\,
            in2 => \_gnd_net_\,
            in3 => \N__17288\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            clk => \N__20868\,
            ce => \N__20663\,
            sr => \N__20401\
        );

    \delay_measurement_inst.delay_hc_timer.counter_27_LC_9_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20532\,
            in1 => \N__19596\,
            in2 => \_gnd_net_\,
            in3 => \N__17285\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            clk => \N__20868\,
            ce => \N__20663\,
            sr => \N__20401\
        );

    \delay_measurement_inst.delay_hc_timer.counter_28_LC_9_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20529\,
            in1 => \N__19646\,
            in2 => \_gnd_net_\,
            in3 => \N__17282\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_28\,
            clk => \N__20868\,
            ce => \N__20663\,
            sr => \N__20401\
        );

    \delay_measurement_inst.delay_hc_timer.counter_29_LC_9_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__19610\,
            in1 => \N__20530\,
            in2 => \_gnd_net_\,
            in3 => \N__17279\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20868\,
            ce => \N__20663\,
            sr => \N__20401\
        );

    \phase_controller_slave.S1_LC_9_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17276\,
            lcout => s3_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20864\,
            ce => 'H',
            sr => \N__20421\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17237\,
            lcout => \delay_measurement_inst.elapsed_time_tr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20917\,
            ce => \N__17195\,
            sr => \N__20351\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17216\,
            lcout => \delay_measurement_inst.elapsed_time_tr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20917\,
            ce => \N__17195\,
            sr => \N__20351\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__17745\,
            in1 => \N__17388\,
            in2 => \N__18616\,
            in3 => \N__17337\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5OTB1_6_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18077\,
            in2 => \N__17570\,
            in3 => \N__17960\,
            lcout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20071\,
            lcout => \delay_measurement_inst.delay_tr_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17428\,
            in2 => \_gnd_net_\,
            in3 => \N__17413\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_177_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIF2PP_1_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__18043\,
            in1 => \N__17395\,
            in2 => \N__17371\,
            in3 => \N__17344\,
            lcout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17324\,
            in1 => \N__17318\,
            in2 => \N__17312\,
            in3 => \N__17303\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC841_7_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17871\,
            in1 => \N__17920\,
            in2 => \N__18056\,
            in3 => \N__18741\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQMG82_16_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__17788\,
            in1 => \N__17769\,
            in2 => \N__17297\,
            in3 => \N__17809\,
            lcout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKTUL_6_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__17921\,
            in1 => \N__18089\,
            in2 => \_gnd_net_\,
            in3 => \N__17970\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICHJG3_1_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__17810\,
            in1 => \N__17801\,
            in2 => \N__17795\,
            in3 => \N__18005\,
            lcout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__17787\,
            in1 => \N__18612\,
            in2 => \N__17773\,
            in3 => \N__17746\,
            lcout => \delay_measurement_inst.N_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17729\,
            in2 => \_gnd_net_\,
            in3 => \N__17723\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17717\,
            in1 => \N__17696\,
            in2 => \N__17674\,
            in3 => \N__17653\,
            lcout => \delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17636\,
            in1 => \N__17630\,
            in2 => \N__17624\,
            in3 => \N__17615\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17609\,
            in1 => \N__17603\,
            in2 => \N__17597\,
            in3 => \N__17594\,
            lcout => \delay_measurement_inst.N_35\,
            ltout => \delay_measurement_inst.N_35_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_6_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__18122\,
            in1 => \N__17588\,
            in2 => \N__17579\,
            in3 => \N__17576\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_177\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__18578\,
            in1 => \N__18127\,
            in2 => \N__18107\,
            in3 => \N__17940\,
            lcout => \delay_measurement_inst.N_164\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__18748\,
            in1 => \N__17878\,
            in2 => \N__18128\,
            in3 => \N__18575\,
            lcout => \delay_measurement_inst.N_187\,
            ltout => \delay_measurement_inst.N_187_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__18176\,
            in1 => \N__18647\,
            in2 => \N__18167\,
            in3 => \N__18164\,
            lcout => \delay_measurement_inst.un3_elapsed_time_tr_0_i\,
            ltout => \delay_measurement_inst.un3_elapsed_time_tr_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_31_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__20461\,
            in1 => \_gnd_net_\,
            in2 => \N__18158\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010001"
        )
    port map (
            in0 => \N__18576\,
            in1 => \N__17939\,
            in2 => \N__18022\,
            in3 => \N__18058\,
            lcout => \delay_measurement_inst.N_162_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000110011"
        )
    port map (
            in0 => \N__18126\,
            in1 => \N__17937\,
            in2 => \N__18106\,
            in3 => \N__18057\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.N_180_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010100"
        )
    port map (
            in0 => \N__18577\,
            in1 => \N__18018\,
            in2 => \N__17984\,
            in3 => \N__18648\,
            lcout => \delay_measurement_inst.N_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI654I_6_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17977\,
            in2 => \_gnd_net_\,
            in3 => \N__17938\,
            lcout => \delay_measurement_inst.delay_tr_reg_5_0_a2_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_7_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__18772\,
            in1 => \N__18787\,
            in2 => \N__17849\,
            in3 => \N__17879\,
            lcout => measured_delay_tr_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20892\,
            ce => 'H',
            sr => \N__20366\
        );

    \delay_measurement_inst.delay_tr_reg_8_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__18788\,
            in1 => \N__18773\,
            in2 => \N__18721\,
            in3 => \N__18749\,
            lcout => measured_delay_tr_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20892\,
            ce => 'H',
            sr => \N__20366\
        );

    \delay_measurement_inst.delay_tr_reg_esr_19_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__18687\,
            in1 => \N__18620\,
            in2 => \_gnd_net_\,
            in3 => \N__18590\,
            lcout => measured_delay_tr_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20885\,
            ce => \N__18506\,
            sr => \N__20371\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18484\,
            in2 => \N__18397\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.elapsed_time_hc_3\,
            ltout => OPEN,
            carryin => \bfn_10_21_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__20873\,
            ce => \N__19495\,
            sr => \N__20375\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18442\,
            in2 => \N__18355\,
            in3 => \N__18401\,
            lcout => \delay_measurement_inst.elapsed_time_hc_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__20873\,
            ce => \N__19495\,
            sr => \N__20375\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18294\,
            in2 => \N__18398\,
            in3 => \N__18359\,
            lcout => \delay_measurement_inst.elapsed_time_hc_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__20873\,
            ce => \N__19495\,
            sr => \N__20375\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18249\,
            in2 => \N__18356\,
            in3 => \N__18299\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__20873\,
            ce => \N__19495\,
            sr => \N__20375\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18295\,
            in2 => \N__19174\,
            in3 => \N__18254\,
            lcout => \delay_measurement_inst.elapsed_time_hc_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__20873\,
            ce => \N__19495\,
            sr => \N__20375\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18250\,
            in2 => \N__19105\,
            in3 => \N__18206\,
            lcout => \delay_measurement_inst.elapsed_time_hc_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__20873\,
            ce => \N__19495\,
            sr => \N__20375\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19062\,
            in2 => \N__19175\,
            in3 => \N__19109\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__20873\,
            ce => \N__19495\,
            sr => \N__20375\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19023\,
            in2 => \N__19106\,
            in3 => \N__19067\,
            lcout => \delay_measurement_inst.elapsed_time_hc_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__20873\,
            ce => \N__19495\,
            sr => \N__20375\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19064\,
            in2 => \N__18985\,
            in3 => \N__19028\,
            lcout => \delay_measurement_inst.elapsed_time_hc_11\,
            ltout => OPEN,
            carryin => \bfn_10_22_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__20869\,
            ce => \N__19494\,
            sr => \N__20381\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19025\,
            in2 => \N__18937\,
            in3 => \N__18989\,
            lcout => \delay_measurement_inst.elapsed_time_hc_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__20869\,
            ce => \N__19494\,
            sr => \N__20381\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18867\,
            in2 => \N__18986\,
            in3 => \N__18941\,
            lcout => \delay_measurement_inst.elapsed_time_hc_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__20869\,
            ce => \N__19494\,
            sr => \N__20381\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19473\,
            in2 => \N__18938\,
            in3 => \N__18872\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__20869\,
            ce => \N__19494\,
            sr => \N__20381\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18868\,
            in2 => \N__19429\,
            in3 => \N__18791\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__20869\,
            ce => \N__19494\,
            sr => \N__20381\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19474\,
            in2 => \N__19375\,
            in3 => \N__19433\,
            lcout => \delay_measurement_inst.elapsed_time_hc_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__20869\,
            ce => \N__19494\,
            sr => \N__20381\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19326\,
            in2 => \N__19430\,
            in3 => \N__19379\,
            lcout => \delay_measurement_inst.elapsed_time_hc_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__20869\,
            ce => \N__19494\,
            sr => \N__20381\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19275\,
            in2 => \N__19376\,
            in3 => \N__19331\,
            lcout => \delay_measurement_inst.elapsed_time_hc_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__20869\,
            ce => \N__19494\,
            sr => \N__20381\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19328\,
            in2 => \N__19255\,
            in3 => \N__19280\,
            lcout => \delay_measurement_inst.elapsed_time_hc_19\,
            ltout => OPEN,
            carryin => \bfn_10_23_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__20867\,
            ce => \N__19493\,
            sr => \N__20389\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19277\,
            in2 => \N__19231\,
            in3 => \N__19259\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__20867\,
            ce => \N__19493\,
            sr => \N__20389\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19206\,
            in2 => \N__19256\,
            in3 => \N__19235\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__20867\,
            ce => \N__19493\,
            sr => \N__20389\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19188\,
            in2 => \N__19232\,
            in3 => \N__19211\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__20867\,
            ce => \N__19493\,
            sr => \N__20389\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19207\,
            in2 => \N__19735\,
            in3 => \N__19193\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__20867\,
            ce => \N__19493\,
            sr => \N__20389\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19189\,
            in2 => \N__19711\,
            in3 => \N__19739\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__20867\,
            ce => \N__19493\,
            sr => \N__20389\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19686\,
            in2 => \N__19736\,
            in3 => \N__19715\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__20867\,
            ce => \N__19493\,
            sr => \N__20389\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_10_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19665\,
            in2 => \N__19712\,
            in3 => \N__19691\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__20867\,
            ce => \N__19493\,
            sr => \N__20389\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_10_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19688\,
            in2 => \N__19633\,
            in3 => \N__19670\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\,
            ltout => OPEN,
            carryin => \bfn_10_24_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__20865\,
            ce => \N__19492\,
            sr => \N__20394\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19667\,
            in2 => \N__19597\,
            in3 => \N__19649\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__20865\,
            ce => \N__19492\,
            sr => \N__20394\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_10_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19645\,
            in2 => \N__19634\,
            in3 => \N__19613\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__20865\,
            ce => \N__19492\,
            sr => \N__20394\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_10_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19609\,
            in2 => \N__19598\,
            in3 => \N__19577\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__20865\,
            ce => \N__19492\,
            sr => \N__20394\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_10_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19574\,
            lcout => \delay_measurement_inst.elapsed_time_hc_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20865\,
            ce => \N__19492\,
            sr => \N__20394\
        );

    \delay_measurement_inst.delay_tr_timer.running_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__20102\,
            in1 => \N__20090\,
            in2 => \_gnd_net_\,
            in3 => \N__20072\,
            lcout => \delay_measurement_inst.delay_tr_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20911\,
            ce => 'H',
            sr => \N__20350\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20089\,
            in2 => \_gnd_net_\,
            in3 => \N__20069\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_255_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.S2_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19919\,
            lcout => s2_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20878\,
            ce => 'H',
            sr => \N__20367\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19865\,
            in1 => \N__19859\,
            in2 => \N__19853\,
            in3 => \N__19844\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_o2_7_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19838\,
            in1 => \N__19763\,
            in2 => \N__19832\,
            in3 => \N__19745\,
            lcout => \delay_measurement_inst.N_276\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAAI01_25_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19790\,
            in1 => \N__19784\,
            in2 => \N__19778\,
            in3 => \N__19769\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_o2_6_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI23AG_29_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19757\,
            in2 => \_gnd_net_\,
            in3 => \N__19751\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_o2_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.start_timer_tr_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001100110"
        )
    port map (
            in0 => \N__19973\,
            in1 => \N__20009\,
            in2 => \_gnd_net_\,
            in3 => \N__19989\,
            lcout => \delay_measurement_inst.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20910\,
            ce => 'H',
            sr => \N__20346\
        );

    \delay_measurement_inst.prev_tr_sig_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20010\,
            lcout => \delay_measurement_inst.prev_tr_sigZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20910\,
            ce => 'H',
            sr => \N__20346\
        );

    \delay_measurement_inst.stop_timer_tr_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__20012\,
            in1 => \N__19972\,
            in2 => \N__20467\,
            in3 => \N__19990\,
            lcout => \delay_measurement_inst.stop_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20906\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__20101\,
            in1 => \N__20088\,
            in2 => \_gnd_net_\,
            in3 => \N__20070\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_256_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_TR2_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20018\,
            lcout => delay_tr_d2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20918\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_TR1_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20036\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => delay_tr_d1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20918\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.tr_state_0_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001100110"
        )
    port map (
            in0 => \N__20011\,
            in1 => \N__19971\,
            in2 => \_gnd_net_\,
            in3 => \N__19991\,
            lcout => \delay_measurement_inst.tr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20912\,
            ce => \N__20188\,
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_HC2_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19940\,
            lcout => delay_hc_d2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20893\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_HC1_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19955\,
            lcout => delay_hc_d1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20893\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.hc_state_0_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__21008\,
            in1 => \N__20982\,
            in2 => \_gnd_net_\,
            in3 => \N__20955\,
            lcout => \delay_measurement_inst.hc_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20886\,
            ce => \N__20171\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_hc_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__21004\,
            in1 => \N__20983\,
            in2 => \N__20468\,
            in3 => \N__20964\,
            lcout => \delay_measurement_inst.stop_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20879\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.prev_hc_sig_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20966\,
            lcout => \delay_measurement_inst.prev_hc_sigZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20874\,
            ce => 'H',
            sr => \N__20360\
        );

    \delay_measurement_inst.start_timer_hc_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__21003\,
            in1 => \N__20987\,
            in2 => \_gnd_net_\,
            in3 => \N__20965\,
            lcout => \delay_measurement_inst.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20874\,
            ce => 'H',
            sr => \N__20360\
        );

    \delay_measurement_inst.delay_hc_timer.running_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__20679\,
            in1 => \N__20693\,
            in2 => \_gnd_net_\,
            in3 => \N__20615\,
            lcout => \delay_measurement_inst.delay_hc_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20874\,
            ce => 'H',
            sr => \N__20360\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20680\,
            in2 => \_gnd_net_\,
            in3 => \N__20612\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_253_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__20692\,
            in1 => \N__20681\,
            in2 => \_gnd_net_\,
            in3 => \N__20614\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_254_i_g\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_13_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20613\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_ibuf_gb_io_RNI79U7_LC_13_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20462\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => red_c_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
