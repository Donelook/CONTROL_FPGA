-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Oct 20 2025 00:15:25

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MAIN" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MAIN
entity MAIN is
port (
    start_stop : in std_logic;
    s2_phy : out std_logic;
    T23 : out std_logic;
    s3_phy : out std_logic;
    il_min_comp2 : in std_logic;
    il_max_comp1 : in std_logic;
    s1_phy : out std_logic;
    reset : in std_logic;
    il_min_comp1 : in std_logic;
    delay_tr_input : in std_logic;
    T12 : out std_logic;
    s4_phy : out std_logic;
    rgb_g : out std_logic;
    rgb_r : out std_logic;
    rgb_b : out std_logic;
    pwm_output : out std_logic;
    il_max_comp2 : in std_logic;
    delay_hc_input : in std_logic);
end MAIN;

-- Architecture of MAIN
-- View name is \INTERFACE\
architecture \INTERFACE\ of MAIN is

signal \N__21833\ : std_logic;
signal \N__21832\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21784\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21766\ : std_logic;
signal \N__21759\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21748\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21739\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21681\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21679\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21676\ : std_logic;
signal \N__21675\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21594\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21575\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21534\ : std_logic;
signal \N__21531\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21499\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21480\ : std_logic;
signal \N__21477\ : std_logic;
signal \N__21474\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21419\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21387\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21370\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21367\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21339\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21311\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21282\ : std_logic;
signal \N__21279\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21249\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21223\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21193\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21188\ : std_logic;
signal \N__21187\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21184\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21163\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21148\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21124\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21112\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20902\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20899\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20880\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20863\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20835\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20832\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20827\ : std_logic;
signal \N__20826\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20823\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20821\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20818\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20800\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20794\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20791\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20788\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20785\ : std_logic;
signal \N__20784\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20779\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20776\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20766\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20760\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20589\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20570\ : std_logic;
signal \N__20567\ : std_logic;
signal \N__20564\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20553\ : std_logic;
signal \N__20550\ : std_logic;
signal \N__20547\ : std_logic;
signal \N__20544\ : std_logic;
signal \N__20541\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20511\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20478\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20451\ : std_logic;
signal \N__20448\ : std_logic;
signal \N__20445\ : std_logic;
signal \N__20442\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20403\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20376\ : std_logic;
signal \N__20373\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20364\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20353\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20347\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20308\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20302\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20288\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20261\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20257\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20209\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20202\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20173\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20080\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20070\ : std_logic;
signal \N__20067\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19986\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19930\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19923\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19702\ : std_logic;
signal \N__19699\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19674\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19657\ : std_logic;
signal \N__19654\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19648\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19633\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19620\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19612\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19591\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19557\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19545\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19485\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19476\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19449\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19437\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19389\ : std_logic;
signal \N__19386\ : std_logic;
signal \N__19383\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19353\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19303\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19284\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19281\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19279\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19276\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19273\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19269\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19166\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19137\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19131\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19086\ : std_logic;
signal \N__19083\ : std_logic;
signal \N__19080\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19069\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19057\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19045\ : std_logic;
signal \N__19044\ : std_logic;
signal \N__19041\ : std_logic;
signal \N__19038\ : std_logic;
signal \N__19035\ : std_logic;
signal \N__19032\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19012\ : std_logic;
signal \N__19009\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18999\ : std_logic;
signal \N__18996\ : std_logic;
signal \N__18993\ : std_logic;
signal \N__18990\ : std_logic;
signal \N__18987\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18963\ : std_logic;
signal \N__18960\ : std_logic;
signal \N__18957\ : std_logic;
signal \N__18950\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18936\ : std_logic;
signal \N__18933\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18924\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18912\ : std_logic;
signal \N__18909\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18866\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18847\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18829\ : std_logic;
signal \N__18826\ : std_logic;
signal \N__18823\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18811\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18795\ : std_logic;
signal \N__18792\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18769\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18762\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18734\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18728\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18723\ : std_logic;
signal \N__18722\ : std_logic;
signal \N__18721\ : std_logic;
signal \N__18720\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18714\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18711\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18708\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18705\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18702\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18699\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18697\ : std_logic;
signal \N__18696\ : std_logic;
signal \N__18687\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18669\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18621\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18605\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18595\ : std_logic;
signal \N__18594\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18577\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18541\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18478\ : std_logic;
signal \N__18475\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18458\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18436\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18400\ : std_logic;
signal \N__18397\ : std_logic;
signal \N__18394\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18373\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18352\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18328\ : std_logic;
signal \N__18325\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18310\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18304\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18293\ : std_logic;
signal \N__18290\ : std_logic;
signal \N__18289\ : std_logic;
signal \N__18286\ : std_logic;
signal \N__18283\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18272\ : std_logic;
signal \N__18269\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18265\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18247\ : std_logic;
signal \N__18246\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18240\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18224\ : std_logic;
signal \N__18221\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18214\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18196\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18190\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18182\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18164\ : std_logic;
signal \N__18163\ : std_logic;
signal \N__18160\ : std_logic;
signal \N__18157\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18149\ : std_logic;
signal \N__18146\ : std_logic;
signal \N__18143\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18139\ : std_logic;
signal \N__18136\ : std_logic;
signal \N__18133\ : std_logic;
signal \N__18128\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18119\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18112\ : std_logic;
signal \N__18109\ : std_logic;
signal \N__18106\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18092\ : std_logic;
signal \N__18091\ : std_logic;
signal \N__18088\ : std_logic;
signal \N__18085\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18064\ : std_logic;
signal \N__18061\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18040\ : std_logic;
signal \N__18039\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18031\ : std_logic;
signal \N__18028\ : std_logic;
signal \N__18025\ : std_logic;
signal \N__18024\ : std_logic;
signal \N__18019\ : std_logic;
signal \N__18016\ : std_logic;
signal \N__18009\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__18001\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17995\ : std_logic;
signal \N__17992\ : std_logic;
signal \N__17989\ : std_logic;
signal \N__17986\ : std_logic;
signal \N__17983\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17975\ : std_logic;
signal \N__17974\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17972\ : std_logic;
signal \N__17969\ : std_logic;
signal \N__17966\ : std_logic;
signal \N__17965\ : std_logic;
signal \N__17964\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17962\ : std_logic;
signal \N__17961\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17955\ : std_logic;
signal \N__17950\ : std_logic;
signal \N__17945\ : std_logic;
signal \N__17936\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17917\ : std_logic;
signal \N__17916\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17914\ : std_logic;
signal \N__17913\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17902\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17884\ : std_logic;
signal \N__17881\ : std_logic;
signal \N__17880\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17878\ : std_logic;
signal \N__17875\ : std_logic;
signal \N__17872\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17854\ : std_logic;
signal \N__17851\ : std_logic;
signal \N__17848\ : std_logic;
signal \N__17845\ : std_logic;
signal \N__17842\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17833\ : std_logic;
signal \N__17832\ : std_logic;
signal \N__17827\ : std_logic;
signal \N__17826\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17821\ : std_logic;
signal \N__17820\ : std_logic;
signal \N__17819\ : std_logic;
signal \N__17818\ : std_logic;
signal \N__17815\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17799\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17797\ : std_logic;
signal \N__17796\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17794\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17783\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17775\ : std_logic;
signal \N__17772\ : std_logic;
signal \N__17769\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17759\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17745\ : std_logic;
signal \N__17738\ : std_logic;
signal \N__17735\ : std_logic;
signal \N__17734\ : std_logic;
signal \N__17731\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17725\ : std_logic;
signal \N__17722\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17711\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17702\ : std_logic;
signal \N__17697\ : std_logic;
signal \N__17690\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17686\ : std_logic;
signal \N__17683\ : std_logic;
signal \N__17682\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17678\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17669\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17659\ : std_logic;
signal \N__17658\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17656\ : std_logic;
signal \N__17645\ : std_logic;
signal \N__17642\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17638\ : std_logic;
signal \N__17637\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17627\ : std_logic;
signal \N__17626\ : std_logic;
signal \N__17625\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17623\ : std_logic;
signal \N__17622\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17620\ : std_logic;
signal \N__17619\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17614\ : std_logic;
signal \N__17609\ : std_logic;
signal \N__17600\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17590\ : std_logic;
signal \N__17589\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17587\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17577\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17575\ : std_logic;
signal \N__17574\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17572\ : std_logic;
signal \N__17571\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17539\ : std_logic;
signal \N__17538\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17536\ : std_logic;
signal \N__17533\ : std_logic;
signal \N__17526\ : std_logic;
signal \N__17517\ : std_logic;
signal \N__17512\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17506\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17500\ : std_logic;
signal \N__17499\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17489\ : std_logic;
signal \N__17486\ : std_logic;
signal \N__17481\ : std_logic;
signal \N__17478\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17472\ : std_logic;
signal \N__17469\ : std_logic;
signal \N__17466\ : std_logic;
signal \N__17463\ : std_logic;
signal \N__17460\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17452\ : std_logic;
signal \N__17451\ : std_logic;
signal \N__17448\ : std_logic;
signal \N__17445\ : std_logic;
signal \N__17442\ : std_logic;
signal \N__17439\ : std_logic;
signal \N__17438\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17421\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17407\ : std_logic;
signal \N__17404\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17400\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17384\ : std_logic;
signal \N__17381\ : std_logic;
signal \N__17378\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17370\ : std_logic;
signal \N__17363\ : std_logic;
signal \N__17362\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17355\ : std_logic;
signal \N__17352\ : std_logic;
signal \N__17349\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17342\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17324\ : std_logic;
signal \N__17321\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17317\ : std_logic;
signal \N__17314\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17297\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17275\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17265\ : std_logic;
signal \N__17264\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17258\ : std_logic;
signal \N__17255\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17243\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17239\ : std_logic;
signal \N__17238\ : std_logic;
signal \N__17235\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17229\ : std_logic;
signal \N__17224\ : std_logic;
signal \N__17221\ : std_logic;
signal \N__17218\ : std_logic;
signal \N__17217\ : std_logic;
signal \N__17214\ : std_logic;
signal \N__17211\ : std_logic;
signal \N__17208\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17189\ : std_logic;
signal \N__17186\ : std_logic;
signal \N__17185\ : std_logic;
signal \N__17184\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17172\ : std_logic;
signal \N__17169\ : std_logic;
signal \N__17166\ : std_logic;
signal \N__17163\ : std_logic;
signal \N__17160\ : std_logic;
signal \N__17157\ : std_logic;
signal \N__17154\ : std_logic;
signal \N__17151\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17145\ : std_logic;
signal \N__17142\ : std_logic;
signal \N__17137\ : std_logic;
signal \N__17132\ : std_logic;
signal \N__17129\ : std_logic;
signal \N__17120\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17114\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17108\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17103\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17090\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17084\ : std_logic;
signal \N__17081\ : std_logic;
signal \N__17078\ : std_logic;
signal \N__17075\ : std_logic;
signal \N__17072\ : std_logic;
signal \N__17069\ : std_logic;
signal \N__17066\ : std_logic;
signal \N__17063\ : std_logic;
signal \N__17060\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17054\ : std_logic;
signal \N__17051\ : std_logic;
signal \N__17048\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17040\ : std_logic;
signal \N__17039\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17033\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17009\ : std_logic;
signal \N__17006\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16999\ : std_logic;
signal \N__16996\ : std_logic;
signal \N__16993\ : std_logic;
signal \N__16990\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16984\ : std_logic;
signal \N__16983\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16981\ : std_logic;
signal \N__16980\ : std_logic;
signal \N__16977\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16975\ : std_logic;
signal \N__16974\ : std_logic;
signal \N__16971\ : std_logic;
signal \N__16968\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16952\ : std_logic;
signal \N__16949\ : std_logic;
signal \N__16934\ : std_logic;
signal \N__16933\ : std_logic;
signal \N__16930\ : std_logic;
signal \N__16927\ : std_logic;
signal \N__16926\ : std_logic;
signal \N__16925\ : std_logic;
signal \N__16920\ : std_logic;
signal \N__16917\ : std_logic;
signal \N__16914\ : std_logic;
signal \N__16911\ : std_logic;
signal \N__16908\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16900\ : std_logic;
signal \N__16897\ : std_logic;
signal \N__16892\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16888\ : std_logic;
signal \N__16887\ : std_logic;
signal \N__16886\ : std_logic;
signal \N__16883\ : std_logic;
signal \N__16880\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16871\ : std_logic;
signal \N__16866\ : std_logic;
signal \N__16863\ : std_logic;
signal \N__16860\ : std_logic;
signal \N__16855\ : std_logic;
signal \N__16850\ : std_logic;
signal \N__16847\ : std_logic;
signal \N__16846\ : std_logic;
signal \N__16843\ : std_logic;
signal \N__16840\ : std_logic;
signal \N__16837\ : std_logic;
signal \N__16836\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16832\ : std_logic;
signal \N__16829\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16814\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16808\ : std_logic;
signal \N__16805\ : std_logic;
signal \N__16802\ : std_logic;
signal \N__16801\ : std_logic;
signal \N__16798\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16792\ : std_logic;
signal \N__16791\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16789\ : std_logic;
signal \N__16786\ : std_logic;
signal \N__16783\ : std_logic;
signal \N__16776\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16766\ : std_logic;
signal \N__16763\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16756\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16750\ : std_logic;
signal \N__16747\ : std_logic;
signal \N__16744\ : std_logic;
signal \N__16743\ : std_logic;
signal \N__16740\ : std_logic;
signal \N__16737\ : std_logic;
signal \N__16734\ : std_logic;
signal \N__16727\ : std_logic;
signal \N__16724\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16719\ : std_logic;
signal \N__16718\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16716\ : std_logic;
signal \N__16715\ : std_logic;
signal \N__16714\ : std_logic;
signal \N__16713\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16711\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16686\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16684\ : std_logic;
signal \N__16683\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16681\ : std_logic;
signal \N__16680\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16678\ : std_logic;
signal \N__16677\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16675\ : std_logic;
signal \N__16672\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16656\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16642\ : std_logic;
signal \N__16639\ : std_logic;
signal \N__16632\ : std_logic;
signal \N__16629\ : std_logic;
signal \N__16622\ : std_logic;
signal \N__16621\ : std_logic;
signal \N__16620\ : std_logic;
signal \N__16617\ : std_logic;
signal \N__16614\ : std_logic;
signal \N__16611\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16609\ : std_logic;
signal \N__16608\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16606\ : std_logic;
signal \N__16605\ : std_logic;
signal \N__16604\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16602\ : std_logic;
signal \N__16601\ : std_logic;
signal \N__16590\ : std_logic;
signal \N__16587\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16581\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16579\ : std_logic;
signal \N__16576\ : std_logic;
signal \N__16567\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16565\ : std_logic;
signal \N__16564\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16562\ : std_logic;
signal \N__16559\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16545\ : std_logic;
signal \N__16542\ : std_logic;
signal \N__16531\ : std_logic;
signal \N__16528\ : std_logic;
signal \N__16521\ : std_logic;
signal \N__16514\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16510\ : std_logic;
signal \N__16507\ : std_logic;
signal \N__16506\ : std_logic;
signal \N__16503\ : std_logic;
signal \N__16500\ : std_logic;
signal \N__16497\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16487\ : std_logic;
signal \N__16484\ : std_logic;
signal \N__16481\ : std_logic;
signal \N__16480\ : std_logic;
signal \N__16477\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16468\ : std_logic;
signal \N__16467\ : std_logic;
signal \N__16464\ : std_logic;
signal \N__16461\ : std_logic;
signal \N__16458\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16448\ : std_logic;
signal \N__16445\ : std_logic;
signal \N__16442\ : std_logic;
signal \N__16441\ : std_logic;
signal \N__16440\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16438\ : std_logic;
signal \N__16437\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16435\ : std_logic;
signal \N__16434\ : std_logic;
signal \N__16431\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16429\ : std_logic;
signal \N__16428\ : std_logic;
signal \N__16425\ : std_logic;
signal \N__16422\ : std_logic;
signal \N__16419\ : std_logic;
signal \N__16416\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16413\ : std_logic;
signal \N__16412\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16400\ : std_logic;
signal \N__16399\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16393\ : std_logic;
signal \N__16380\ : std_logic;
signal \N__16377\ : std_logic;
signal \N__16374\ : std_logic;
signal \N__16373\ : std_logic;
signal \N__16372\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16370\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16366\ : std_logic;
signal \N__16363\ : std_logic;
signal \N__16360\ : std_logic;
signal \N__16357\ : std_logic;
signal \N__16356\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16352\ : std_logic;
signal \N__16347\ : std_logic;
signal \N__16330\ : std_logic;
signal \N__16329\ : std_logic;
signal \N__16326\ : std_logic;
signal \N__16315\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16307\ : std_logic;
signal \N__16298\ : std_logic;
signal \N__16295\ : std_logic;
signal \N__16292\ : std_logic;
signal \N__16289\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16284\ : std_logic;
signal \N__16283\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16277\ : std_logic;
signal \N__16272\ : std_logic;
signal \N__16265\ : std_logic;
signal \N__16262\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16260\ : std_logic;
signal \N__16259\ : std_logic;
signal \N__16256\ : std_logic;
signal \N__16253\ : std_logic;
signal \N__16248\ : std_logic;
signal \N__16245\ : std_logic;
signal \N__16242\ : std_logic;
signal \N__16239\ : std_logic;
signal \N__16232\ : std_logic;
signal \N__16229\ : std_logic;
signal \N__16228\ : std_logic;
signal \N__16227\ : std_logic;
signal \N__16226\ : std_logic;
signal \N__16223\ : std_logic;
signal \N__16220\ : std_logic;
signal \N__16215\ : std_logic;
signal \N__16212\ : std_logic;
signal \N__16209\ : std_logic;
signal \N__16206\ : std_logic;
signal \N__16199\ : std_logic;
signal \N__16196\ : std_logic;
signal \N__16195\ : std_logic;
signal \N__16194\ : std_logic;
signal \N__16193\ : std_logic;
signal \N__16190\ : std_logic;
signal \N__16187\ : std_logic;
signal \N__16184\ : std_logic;
signal \N__16181\ : std_logic;
signal \N__16176\ : std_logic;
signal \N__16171\ : std_logic;
signal \N__16166\ : std_logic;
signal \N__16165\ : std_logic;
signal \N__16162\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16160\ : std_logic;
signal \N__16157\ : std_logic;
signal \N__16154\ : std_logic;
signal \N__16149\ : std_logic;
signal \N__16146\ : std_logic;
signal \N__16141\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16133\ : std_logic;
signal \N__16132\ : std_logic;
signal \N__16127\ : std_logic;
signal \N__16124\ : std_logic;
signal \N__16123\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16119\ : std_logic;
signal \N__16114\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16106\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16102\ : std_logic;
signal \N__16101\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16097\ : std_logic;
signal \N__16094\ : std_logic;
signal \N__16091\ : std_logic;
signal \N__16088\ : std_logic;
signal \N__16085\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16076\ : std_logic;
signal \N__16071\ : std_logic;
signal \N__16064\ : std_logic;
signal \N__16063\ : std_logic;
signal \N__16062\ : std_logic;
signal \N__16059\ : std_logic;
signal \N__16056\ : std_logic;
signal \N__16053\ : std_logic;
signal \N__16052\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16048\ : std_logic;
signal \N__16043\ : std_logic;
signal \N__16038\ : std_logic;
signal \N__16031\ : std_logic;
signal \N__16028\ : std_logic;
signal \N__16025\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16019\ : std_logic;
signal \N__16016\ : std_logic;
signal \N__16015\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16011\ : std_logic;
signal \N__16006\ : std_logic;
signal \N__16005\ : std_logic;
signal \N__16002\ : std_logic;
signal \N__15999\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15991\ : std_logic;
signal \N__15988\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15973\ : std_logic;
signal \N__15972\ : std_logic;
signal \N__15969\ : std_logic;
signal \N__15966\ : std_logic;
signal \N__15963\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15953\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15949\ : std_logic;
signal \N__15946\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15937\ : std_logic;
signal \N__15936\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15930\ : std_logic;
signal \N__15927\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15922\ : std_logic;
signal \N__15919\ : std_logic;
signal \N__15916\ : std_logic;
signal \N__15913\ : std_logic;
signal \N__15908\ : std_logic;
signal \N__15899\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15897\ : std_logic;
signal \N__15894\ : std_logic;
signal \N__15891\ : std_logic;
signal \N__15890\ : std_logic;
signal \N__15889\ : std_logic;
signal \N__15888\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15886\ : std_logic;
signal \N__15885\ : std_logic;
signal \N__15884\ : std_logic;
signal \N__15883\ : std_logic;
signal \N__15882\ : std_logic;
signal \N__15879\ : std_logic;
signal \N__15874\ : std_logic;
signal \N__15871\ : std_logic;
signal \N__15868\ : std_logic;
signal \N__15855\ : std_logic;
signal \N__15854\ : std_logic;
signal \N__15853\ : std_logic;
signal \N__15852\ : std_logic;
signal \N__15851\ : std_logic;
signal \N__15850\ : std_logic;
signal \N__15849\ : std_logic;
signal \N__15846\ : std_logic;
signal \N__15843\ : std_logic;
signal \N__15840\ : std_logic;
signal \N__15835\ : std_logic;
signal \N__15834\ : std_logic;
signal \N__15833\ : std_logic;
signal \N__15832\ : std_logic;
signal \N__15831\ : std_logic;
signal \N__15830\ : std_logic;
signal \N__15829\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15824\ : std_logic;
signal \N__15817\ : std_logic;
signal \N__15810\ : std_logic;
signal \N__15807\ : std_logic;
signal \N__15800\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15778\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15764\ : std_logic;
signal \N__15763\ : std_logic;
signal \N__15762\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15756\ : std_logic;
signal \N__15753\ : std_logic;
signal \N__15750\ : std_logic;
signal \N__15743\ : std_logic;
signal \N__15742\ : std_logic;
signal \N__15741\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15739\ : std_logic;
signal \N__15738\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15735\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15732\ : std_logic;
signal \N__15731\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15729\ : std_logic;
signal \N__15728\ : std_logic;
signal \N__15725\ : std_logic;
signal \N__15722\ : std_logic;
signal \N__15719\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15715\ : std_logic;
signal \N__15714\ : std_logic;
signal \N__15713\ : std_logic;
signal \N__15712\ : std_logic;
signal \N__15709\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15703\ : std_logic;
signal \N__15700\ : std_logic;
signal \N__15697\ : std_logic;
signal \N__15694\ : std_logic;
signal \N__15691\ : std_logic;
signal \N__15688\ : std_logic;
signal \N__15687\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15669\ : std_logic;
signal \N__15666\ : std_logic;
signal \N__15657\ : std_logic;
signal \N__15648\ : std_logic;
signal \N__15639\ : std_logic;
signal \N__15636\ : std_logic;
signal \N__15633\ : std_logic;
signal \N__15630\ : std_logic;
signal \N__15627\ : std_logic;
signal \N__15626\ : std_logic;
signal \N__15621\ : std_logic;
signal \N__15618\ : std_logic;
signal \N__15615\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15607\ : std_logic;
signal \N__15604\ : std_logic;
signal \N__15593\ : std_logic;
signal \N__15592\ : std_logic;
signal \N__15591\ : std_logic;
signal \N__15590\ : std_logic;
signal \N__15589\ : std_logic;
signal \N__15588\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15586\ : std_logic;
signal \N__15569\ : std_logic;
signal \N__15568\ : std_logic;
signal \N__15567\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15561\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15559\ : std_logic;
signal \N__15558\ : std_logic;
signal \N__15557\ : std_logic;
signal \N__15556\ : std_logic;
signal \N__15555\ : std_logic;
signal \N__15554\ : std_logic;
signal \N__15553\ : std_logic;
signal \N__15552\ : std_logic;
signal \N__15551\ : std_logic;
signal \N__15550\ : std_logic;
signal \N__15547\ : std_logic;
signal \N__15544\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15514\ : std_logic;
signal \N__15511\ : std_logic;
signal \N__15508\ : std_logic;
signal \N__15505\ : std_logic;
signal \N__15488\ : std_logic;
signal \N__15485\ : std_logic;
signal \N__15482\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15478\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15471\ : std_logic;
signal \N__15468\ : std_logic;
signal \N__15461\ : std_logic;
signal \N__15460\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15454\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15437\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15433\ : std_logic;
signal \N__15432\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15421\ : std_logic;
signal \N__15420\ : std_logic;
signal \N__15419\ : std_logic;
signal \N__15416\ : std_logic;
signal \N__15409\ : std_logic;
signal \N__15404\ : std_logic;
signal \N__15401\ : std_logic;
signal \N__15400\ : std_logic;
signal \N__15397\ : std_logic;
signal \N__15394\ : std_logic;
signal \N__15389\ : std_logic;
signal \N__15388\ : std_logic;
signal \N__15385\ : std_logic;
signal \N__15382\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15375\ : std_logic;
signal \N__15372\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15364\ : std_logic;
signal \N__15363\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15361\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15349\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15343\ : std_logic;
signal \N__15340\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15329\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15325\ : std_logic;
signal \N__15322\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15315\ : std_logic;
signal \N__15312\ : std_logic;
signal \N__15305\ : std_logic;
signal \N__15302\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15297\ : std_logic;
signal \N__15294\ : std_logic;
signal \N__15289\ : std_logic;
signal \N__15284\ : std_logic;
signal \N__15283\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15281\ : std_logic;
signal \N__15280\ : std_logic;
signal \N__15279\ : std_logic;
signal \N__15276\ : std_logic;
signal \N__15273\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15269\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15259\ : std_logic;
signal \N__15252\ : std_logic;
signal \N__15245\ : std_logic;
signal \N__15244\ : std_logic;
signal \N__15243\ : std_logic;
signal \N__15240\ : std_logic;
signal \N__15237\ : std_logic;
signal \N__15234\ : std_logic;
signal \N__15231\ : std_logic;
signal \N__15226\ : std_logic;
signal \N__15223\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15211\ : std_logic;
signal \N__15210\ : std_logic;
signal \N__15207\ : std_logic;
signal \N__15204\ : std_logic;
signal \N__15201\ : std_logic;
signal \N__15196\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15190\ : std_logic;
signal \N__15189\ : std_logic;
signal \N__15186\ : std_logic;
signal \N__15181\ : std_logic;
signal \N__15176\ : std_logic;
signal \N__15173\ : std_logic;
signal \N__15170\ : std_logic;
signal \N__15167\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15160\ : std_logic;
signal \N__15157\ : std_logic;
signal \N__15154\ : std_logic;
signal \N__15149\ : std_logic;
signal \N__15146\ : std_logic;
signal \N__15143\ : std_logic;
signal \N__15142\ : std_logic;
signal \N__15141\ : std_logic;
signal \N__15138\ : std_logic;
signal \N__15135\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15129\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15123\ : std_logic;
signal \N__15116\ : std_logic;
signal \N__15113\ : std_logic;
signal \N__15112\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15108\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15104\ : std_logic;
signal \N__15101\ : std_logic;
signal \N__15098\ : std_logic;
signal \N__15095\ : std_logic;
signal \N__15092\ : std_logic;
signal \N__15089\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15079\ : std_logic;
signal \N__15076\ : std_logic;
signal \N__15071\ : std_logic;
signal \N__15068\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15066\ : std_logic;
signal \N__15063\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15057\ : std_logic;
signal \N__15056\ : std_logic;
signal \N__15051\ : std_logic;
signal \N__15048\ : std_logic;
signal \N__15045\ : std_logic;
signal \N__15042\ : std_logic;
signal \N__15037\ : std_logic;
signal \N__15032\ : std_logic;
signal \N__15029\ : std_logic;
signal \N__15028\ : std_logic;
signal \N__15025\ : std_logic;
signal \N__15022\ : std_logic;
signal \N__15021\ : std_logic;
signal \N__15020\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15014\ : std_logic;
signal \N__15009\ : std_logic;
signal \N__15004\ : std_logic;
signal \N__15001\ : std_logic;
signal \N__14996\ : std_logic;
signal \N__14995\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14991\ : std_logic;
signal \N__14990\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14988\ : std_logic;
signal \N__14987\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14983\ : std_logic;
signal \N__14980\ : std_logic;
signal \N__14977\ : std_logic;
signal \N__14970\ : std_logic;
signal \N__14963\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14949\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14946\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14928\ : std_logic;
signal \N__14925\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14915\ : std_logic;
signal \N__14914\ : std_logic;
signal \N__14911\ : std_logic;
signal \N__14908\ : std_logic;
signal \N__14907\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14903\ : std_logic;
signal \N__14900\ : std_logic;
signal \N__14895\ : std_logic;
signal \N__14892\ : std_logic;
signal \N__14887\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14881\ : std_logic;
signal \N__14878\ : std_logic;
signal \N__14875\ : std_logic;
signal \N__14872\ : std_logic;
signal \N__14869\ : std_logic;
signal \N__14866\ : std_logic;
signal \N__14863\ : std_logic;
signal \N__14862\ : std_logic;
signal \N__14857\ : std_logic;
signal \N__14854\ : std_logic;
signal \N__14849\ : std_logic;
signal \N__14846\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14842\ : std_logic;
signal \N__14841\ : std_logic;
signal \N__14838\ : std_logic;
signal \N__14837\ : std_logic;
signal \N__14834\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14819\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14807\ : std_logic;
signal \N__14806\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14797\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14788\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14784\ : std_logic;
signal \N__14781\ : std_logic;
signal \N__14778\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14768\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14759\ : std_logic;
signal \N__14756\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14750\ : std_logic;
signal \N__14747\ : std_logic;
signal \N__14744\ : std_logic;
signal \N__14741\ : std_logic;
signal \N__14738\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14720\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14711\ : std_logic;
signal \N__14708\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14702\ : std_logic;
signal \N__14699\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14678\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14663\ : std_logic;
signal \N__14660\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14645\ : std_logic;
signal \N__14642\ : std_logic;
signal \N__14639\ : std_logic;
signal \N__14636\ : std_logic;
signal \N__14633\ : std_logic;
signal \N__14630\ : std_logic;
signal \N__14627\ : std_logic;
signal \N__14624\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14615\ : std_logic;
signal \N__14612\ : std_logic;
signal \N__14609\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14600\ : std_logic;
signal \N__14597\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14588\ : std_logic;
signal \N__14585\ : std_logic;
signal \N__14582\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14576\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14567\ : std_logic;
signal \N__14564\ : std_logic;
signal \N__14561\ : std_logic;
signal \N__14558\ : std_logic;
signal \N__14555\ : std_logic;
signal \N__14552\ : std_logic;
signal \N__14549\ : std_logic;
signal \N__14546\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14540\ : std_logic;
signal \N__14537\ : std_logic;
signal \N__14534\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14528\ : std_logic;
signal \N__14525\ : std_logic;
signal \N__14522\ : std_logic;
signal \N__14519\ : std_logic;
signal \N__14516\ : std_logic;
signal \N__14513\ : std_logic;
signal \N__14510\ : std_logic;
signal \N__14507\ : std_logic;
signal \N__14504\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14498\ : std_logic;
signal \N__14495\ : std_logic;
signal \N__14492\ : std_logic;
signal \N__14489\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14483\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14474\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14468\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14444\ : std_logic;
signal \N__14441\ : std_logic;
signal \N__14438\ : std_logic;
signal \N__14435\ : std_logic;
signal \N__14432\ : std_logic;
signal \N__14429\ : std_logic;
signal \N__14426\ : std_logic;
signal \N__14423\ : std_logic;
signal \N__14420\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14411\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14407\ : std_logic;
signal \N__14404\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14397\ : std_logic;
signal \N__14394\ : std_logic;
signal \N__14391\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14380\ : std_logic;
signal \N__14377\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14369\ : std_logic;
signal \N__14366\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14364\ : std_logic;
signal \N__14361\ : std_logic;
signal \N__14356\ : std_logic;
signal \N__14353\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14342\ : std_logic;
signal \N__14341\ : std_logic;
signal \N__14338\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14330\ : std_logic;
signal \N__14327\ : std_logic;
signal \N__14326\ : std_logic;
signal \N__14323\ : std_logic;
signal \N__14320\ : std_logic;
signal \N__14317\ : std_logic;
signal \N__14314\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14308\ : std_logic;
signal \N__14303\ : std_logic;
signal \N__14302\ : std_logic;
signal \N__14301\ : std_logic;
signal \N__14300\ : std_logic;
signal \N__14299\ : std_logic;
signal \N__14296\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14283\ : std_logic;
signal \N__14280\ : std_logic;
signal \N__14279\ : std_logic;
signal \N__14276\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14258\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14256\ : std_logic;
signal \N__14255\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14253\ : std_logic;
signal \N__14252\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14232\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14223\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14216\ : std_logic;
signal \N__14215\ : std_logic;
signal \N__14212\ : std_logic;
signal \N__14211\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14201\ : std_logic;
signal \N__14196\ : std_logic;
signal \N__14193\ : std_logic;
signal \N__14186\ : std_logic;
signal \N__14183\ : std_logic;
signal \N__14182\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14171\ : std_logic;
signal \N__14168\ : std_logic;
signal \N__14167\ : std_logic;
signal \N__14166\ : std_logic;
signal \N__14163\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14153\ : std_logic;
signal \N__14152\ : std_logic;
signal \N__14151\ : std_logic;
signal \N__14148\ : std_logic;
signal \N__14143\ : std_logic;
signal \N__14138\ : std_logic;
signal \N__14137\ : std_logic;
signal \N__14134\ : std_logic;
signal \N__14131\ : std_logic;
signal \N__14130\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14120\ : std_logic;
signal \N__14117\ : std_logic;
signal \N__14116\ : std_logic;
signal \N__14115\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14111\ : std_logic;
signal \N__14108\ : std_logic;
signal \N__14103\ : std_logic;
signal \N__14100\ : std_logic;
signal \N__14095\ : std_logic;
signal \N__14090\ : std_logic;
signal \N__14087\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14082\ : std_logic;
signal \N__14079\ : std_logic;
signal \N__14076\ : std_logic;
signal \N__14073\ : std_logic;
signal \N__14070\ : std_logic;
signal \N__14063\ : std_logic;
signal \N__14060\ : std_logic;
signal \N__14057\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14050\ : std_logic;
signal \N__14045\ : std_logic;
signal \N__14042\ : std_logic;
signal \N__14041\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14027\ : std_logic;
signal \N__14026\ : std_logic;
signal \N__14025\ : std_logic;
signal \N__14018\ : std_logic;
signal \N__14015\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14009\ : std_logic;
signal \N__14006\ : std_logic;
signal \N__14005\ : std_logic;
signal \N__14002\ : std_logic;
signal \N__13999\ : std_logic;
signal \N__13994\ : std_logic;
signal \N__13991\ : std_logic;
signal \N__13988\ : std_logic;
signal \N__13985\ : std_logic;
signal \N__13982\ : std_logic;
signal \N__13979\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13966\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13958\ : std_logic;
signal \N__13955\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13951\ : std_logic;
signal \N__13948\ : std_logic;
signal \N__13945\ : std_logic;
signal \N__13942\ : std_logic;
signal \N__13937\ : std_logic;
signal \N__13934\ : std_logic;
signal \N__13931\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13924\ : std_logic;
signal \N__13923\ : std_logic;
signal \N__13920\ : std_logic;
signal \N__13917\ : std_logic;
signal \N__13916\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13910\ : std_logic;
signal \N__13907\ : std_logic;
signal \N__13904\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13889\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13883\ : std_logic;
signal \N__13882\ : std_logic;
signal \N__13881\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13869\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13856\ : std_logic;
signal \N__13853\ : std_logic;
signal \N__13852\ : std_logic;
signal \N__13851\ : std_logic;
signal \N__13850\ : std_logic;
signal \N__13845\ : std_logic;
signal \N__13842\ : std_logic;
signal \N__13839\ : std_logic;
signal \N__13834\ : std_logic;
signal \N__13831\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13805\ : std_logic;
signal \N__13802\ : std_logic;
signal \N__13799\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13794\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13786\ : std_logic;
signal \N__13783\ : std_logic;
signal \N__13780\ : std_logic;
signal \N__13777\ : std_logic;
signal \N__13774\ : std_logic;
signal \N__13769\ : std_logic;
signal \N__13760\ : std_logic;
signal \N__13757\ : std_logic;
signal \N__13754\ : std_logic;
signal \N__13753\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13748\ : std_logic;
signal \N__13743\ : std_logic;
signal \N__13740\ : std_logic;
signal \N__13737\ : std_logic;
signal \N__13734\ : std_logic;
signal \N__13727\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13719\ : std_logic;
signal \N__13718\ : std_logic;
signal \N__13715\ : std_logic;
signal \N__13714\ : std_logic;
signal \N__13713\ : std_logic;
signal \N__13712\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13704\ : std_logic;
signal \N__13701\ : std_logic;
signal \N__13698\ : std_logic;
signal \N__13695\ : std_logic;
signal \N__13692\ : std_logic;
signal \N__13691\ : std_logic;
signal \N__13688\ : std_logic;
signal \N__13687\ : std_logic;
signal \N__13684\ : std_logic;
signal \N__13677\ : std_logic;
signal \N__13674\ : std_logic;
signal \N__13671\ : std_logic;
signal \N__13668\ : std_logic;
signal \N__13665\ : std_logic;
signal \N__13656\ : std_logic;
signal \N__13649\ : std_logic;
signal \N__13648\ : std_logic;
signal \N__13645\ : std_logic;
signal \N__13642\ : std_logic;
signal \N__13641\ : std_logic;
signal \N__13640\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13634\ : std_logic;
signal \N__13629\ : std_logic;
signal \N__13626\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13620\ : std_logic;
signal \N__13613\ : std_logic;
signal \N__13612\ : std_logic;
signal \N__13611\ : std_logic;
signal \N__13608\ : std_logic;
signal \N__13605\ : std_logic;
signal \N__13602\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13598\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13590\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13580\ : std_logic;
signal \N__13579\ : std_logic;
signal \N__13576\ : std_logic;
signal \N__13575\ : std_logic;
signal \N__13572\ : std_logic;
signal \N__13569\ : std_logic;
signal \N__13566\ : std_logic;
signal \N__13563\ : std_logic;
signal \N__13558\ : std_logic;
signal \N__13557\ : std_logic;
signal \N__13552\ : std_logic;
signal \N__13549\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13538\ : std_logic;
signal \N__13537\ : std_logic;
signal \N__13534\ : std_logic;
signal \N__13531\ : std_logic;
signal \N__13530\ : std_logic;
signal \N__13527\ : std_logic;
signal \N__13524\ : std_logic;
signal \N__13521\ : std_logic;
signal \N__13518\ : std_logic;
signal \N__13513\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13504\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13500\ : std_logic;
signal \N__13497\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13490\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13468\ : std_logic;
signal \N__13467\ : std_logic;
signal \N__13464\ : std_logic;
signal \N__13461\ : std_logic;
signal \N__13458\ : std_logic;
signal \N__13457\ : std_logic;
signal \N__13456\ : std_logic;
signal \N__13453\ : std_logic;
signal \N__13450\ : std_logic;
signal \N__13447\ : std_logic;
signal \N__13444\ : std_logic;
signal \N__13441\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13426\ : std_logic;
signal \N__13423\ : std_logic;
signal \N__13420\ : std_logic;
signal \N__13419\ : std_logic;
signal \N__13418\ : std_logic;
signal \N__13413\ : std_logic;
signal \N__13408\ : std_logic;
signal \N__13405\ : std_logic;
signal \N__13402\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13396\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13390\ : std_logic;
signal \N__13385\ : std_logic;
signal \N__13382\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13376\ : std_logic;
signal \N__13375\ : std_logic;
signal \N__13372\ : std_logic;
signal \N__13369\ : std_logic;
signal \N__13364\ : std_logic;
signal \N__13361\ : std_logic;
signal \N__13358\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13354\ : std_logic;
signal \N__13351\ : std_logic;
signal \N__13348\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13337\ : std_logic;
signal \N__13334\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13330\ : std_logic;
signal \N__13327\ : std_logic;
signal \N__13322\ : std_logic;
signal \N__13319\ : std_logic;
signal \N__13316\ : std_logic;
signal \N__13313\ : std_logic;
signal \N__13312\ : std_logic;
signal \N__13309\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13295\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13288\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13285\ : std_logic;
signal \N__13284\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13282\ : std_logic;
signal \N__13281\ : std_logic;
signal \N__13278\ : std_logic;
signal \N__13275\ : std_logic;
signal \N__13274\ : std_logic;
signal \N__13273\ : std_logic;
signal \N__13272\ : std_logic;
signal \N__13271\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13255\ : std_logic;
signal \N__13254\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13252\ : std_logic;
signal \N__13251\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13249\ : std_logic;
signal \N__13248\ : std_logic;
signal \N__13245\ : std_logic;
signal \N__13242\ : std_logic;
signal \N__13239\ : std_logic;
signal \N__13236\ : std_logic;
signal \N__13233\ : std_logic;
signal \N__13230\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13228\ : std_logic;
signal \N__13227\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13222\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13196\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13178\ : std_logic;
signal \N__13163\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13158\ : std_logic;
signal \N__13155\ : std_logic;
signal \N__13152\ : std_logic;
signal \N__13145\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13141\ : std_logic;
signal \N__13140\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13138\ : std_logic;
signal \N__13137\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13122\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13112\ : std_logic;
signal \N__13109\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13103\ : std_logic;
signal \N__13100\ : std_logic;
signal \N__13097\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13085\ : std_logic;
signal \N__13082\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13075\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13067\ : std_logic;
signal \N__13064\ : std_logic;
signal \N__13061\ : std_logic;
signal \N__13060\ : std_logic;
signal \N__13057\ : std_logic;
signal \N__13054\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13039\ : std_logic;
signal \N__13036\ : std_logic;
signal \N__13033\ : std_logic;
signal \N__13028\ : std_logic;
signal \N__13025\ : std_logic;
signal \N__13022\ : std_logic;
signal \N__13019\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13015\ : std_logic;
signal \N__13012\ : std_logic;
signal \N__13007\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12997\ : std_logic;
signal \N__12994\ : std_logic;
signal \N__12991\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12983\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12974\ : std_logic;
signal \N__12971\ : std_logic;
signal \N__12970\ : std_logic;
signal \N__12967\ : std_logic;
signal \N__12964\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12956\ : std_logic;
signal \N__12953\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12949\ : std_logic;
signal \N__12946\ : std_logic;
signal \N__12943\ : std_logic;
signal \N__12938\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12932\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12917\ : std_logic;
signal \N__12914\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12905\ : std_logic;
signal \N__12902\ : std_logic;
signal \N__12901\ : std_logic;
signal \N__12898\ : std_logic;
signal \N__12895\ : std_logic;
signal \N__12892\ : std_logic;
signal \N__12889\ : std_logic;
signal \N__12884\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12869\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12863\ : std_logic;
signal \N__12862\ : std_logic;
signal \N__12859\ : std_logic;
signal \N__12856\ : std_logic;
signal \N__12851\ : std_logic;
signal \N__12848\ : std_logic;
signal \N__12845\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12836\ : std_logic;
signal \N__12833\ : std_logic;
signal \N__12832\ : std_logic;
signal \N__12829\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12803\ : std_logic;
signal \N__12802\ : std_logic;
signal \N__12799\ : std_logic;
signal \N__12796\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12782\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12772\ : std_logic;
signal \N__12769\ : std_logic;
signal \N__12766\ : std_logic;
signal \N__12761\ : std_logic;
signal \N__12758\ : std_logic;
signal \N__12755\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12751\ : std_logic;
signal \N__12748\ : std_logic;
signal \N__12745\ : std_logic;
signal \N__12740\ : std_logic;
signal \N__12737\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12731\ : std_logic;
signal \N__12728\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12710\ : std_logic;
signal \N__12707\ : std_logic;
signal \N__12704\ : std_logic;
signal \N__12701\ : std_logic;
signal \N__12698\ : std_logic;
signal \N__12697\ : std_logic;
signal \N__12696\ : std_logic;
signal \N__12693\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12687\ : std_logic;
signal \N__12684\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12676\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12668\ : std_logic;
signal \N__12667\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12660\ : std_logic;
signal \N__12657\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12651\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12643\ : std_logic;
signal \N__12640\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12630\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12612\ : std_logic;
signal \N__12611\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12597\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12578\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12557\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12551\ : std_logic;
signal \N__12548\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12542\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12527\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12518\ : std_logic;
signal \N__12515\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12494\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12488\ : std_logic;
signal \N__12487\ : std_logic;
signal \N__12484\ : std_logic;
signal \N__12481\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12472\ : std_logic;
signal \N__12469\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12452\ : std_logic;
signal \N__12451\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12445\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12428\ : std_logic;
signal \N__12425\ : std_logic;
signal \N__12422\ : std_logic;
signal \N__12419\ : std_logic;
signal \N__12416\ : std_logic;
signal \N__12413\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12404\ : std_logic;
signal \N__12401\ : std_logic;
signal \N__12398\ : std_logic;
signal \N__12397\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12391\ : std_logic;
signal \N__12386\ : std_logic;
signal \N__12383\ : std_logic;
signal \N__12380\ : std_logic;
signal \N__12377\ : std_logic;
signal \N__12374\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12370\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12361\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12350\ : std_logic;
signal \N__12347\ : std_logic;
signal \N__12344\ : std_logic;
signal \N__12343\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12334\ : std_logic;
signal \N__12329\ : std_logic;
signal \N__12326\ : std_logic;
signal \N__12323\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12319\ : std_logic;
signal \N__12316\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12307\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12296\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12290\ : std_logic;
signal \N__12289\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12280\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12272\ : std_logic;
signal \N__12269\ : std_logic;
signal \N__12266\ : std_logic;
signal \N__12265\ : std_logic;
signal \N__12262\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12238\ : std_logic;
signal \N__12235\ : std_logic;
signal \N__12232\ : std_logic;
signal \N__12227\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12205\ : std_logic;
signal \N__12202\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12193\ : std_logic;
signal \N__12188\ : std_logic;
signal \N__12185\ : std_logic;
signal \N__12182\ : std_logic;
signal \N__12179\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12173\ : std_logic;
signal \N__12170\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12155\ : std_logic;
signal \N__12152\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12145\ : std_logic;
signal \N__12142\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12128\ : std_logic;
signal \N__12127\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12103\ : std_logic;
signal \N__12100\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12076\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12058\ : std_logic;
signal \N__12055\ : std_logic;
signal \N__12052\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12038\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12031\ : std_logic;
signal \N__12030\ : std_logic;
signal \N__12029\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12020\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12016\ : std_logic;
signal \N__12011\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__12002\ : std_logic;
signal \N__11999\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11984\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11980\ : std_logic;
signal \N__11977\ : std_logic;
signal \N__11974\ : std_logic;
signal \N__11973\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11957\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11947\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11941\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11909\ : std_logic;
signal \N__11906\ : std_logic;
signal \N__11903\ : std_logic;
signal \N__11900\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11897\ : std_logic;
signal \N__11894\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11891\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11858\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11844\ : std_logic;
signal \N__11843\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11841\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11838\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11818\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11808\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11800\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11787\ : std_logic;
signal \N__11786\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11783\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11770\ : std_logic;
signal \N__11767\ : std_logic;
signal \N__11764\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11761\ : std_logic;
signal \N__11758\ : std_logic;
signal \N__11755\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11686\ : std_logic;
signal \N__11683\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11674\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11667\ : std_logic;
signal \N__11658\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11644\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11613\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11578\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11526\ : std_logic;
signal \N__11523\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11486\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11463\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11411\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11403\ : std_logic;
signal \N__11400\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11365\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11359\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11356\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11347\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11341\ : std_logic;
signal \N__11338\ : std_logic;
signal \N__11337\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11319\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11313\ : std_logic;
signal \N__11312\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11294\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11240\ : std_logic;
signal \N__11239\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11223\ : std_logic;
signal \N__11220\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11206\ : std_logic;
signal \N__11203\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11159\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11019\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10921\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10900\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10858\ : std_logic;
signal \N__10857\ : std_logic;
signal \N__10854\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10806\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10791\ : std_logic;
signal \N__10788\ : std_logic;
signal \N__10785\ : std_logic;
signal \N__10782\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10754\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10750\ : std_logic;
signal \N__10749\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10726\ : std_logic;
signal \N__10725\ : std_logic;
signal \N__10722\ : std_logic;
signal \N__10719\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10711\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10698\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10675\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10647\ : std_logic;
signal \N__10644\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10638\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10623\ : std_logic;
signal \N__10620\ : std_logic;
signal \N__10617\ : std_logic;
signal \N__10614\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10578\ : std_logic;
signal \N__10575\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10559\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10551\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10533\ : std_logic;
signal \N__10530\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10506\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10488\ : std_logic;
signal \N__10485\ : std_logic;
signal \N__10482\ : std_logic;
signal \N__10479\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10470\ : std_logic;
signal \N__10467\ : std_logic;
signal \N__10464\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10449\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10422\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10416\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10401\ : std_logic;
signal \N__10398\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10159\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9858\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9750\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9636\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9555\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9546\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9390\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9384\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9344\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9316\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9289\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9202\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9178\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9001\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8941\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8811\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8671\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8665\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8611\ : std_logic;
signal \N__8608\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8530\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8372\ : std_logic;
signal \N__8369\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8360\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8312\ : std_logic;
signal \N__8309\ : std_logic;
signal \N__8306\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8282\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \bfn_1_18_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7\ : std_logic;
signal \bfn_1_19_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15\ : std_logic;
signal \bfn_1_20_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17\ : std_logic;
signal \N_39_i_i\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \rgb_drv_RNOZ0\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIUSZ0Z53\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_slave.stoper_tr.N_60\ : std_logic;
signal \phase_controller_slave.start_timer_trZ0\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_3_18_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_3_19_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_17\ : std_logic;
signal \bfn_3_20_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_slave.tr_time_passed\ : std_logic;
signal \phase_controller_slave.stateZ0Z_0\ : std_logic;
signal \phase_controller_slave.start_timer_tr_0_sqmuxa\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ1Z_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.stoper_state_RNII60DZ0Z_1\ : std_logic;
signal il_max_comp2_c : std_logic;
signal il_min_comp2_c : std_logic;
signal \il_min_comp2_D1\ : std_logic;
signal \il_max_comp2_D1\ : std_logic;
signal \phase_controller_slave.start_timer_hc_0_sqmuxa\ : std_logic;
signal \phase_controller_slave.start_timer_hc_RNOZ0Z_0\ : std_logic;
signal \il_min_comp2_D2\ : std_logic;
signal \phase_controller_slave.stateZ0Z_2\ : std_logic;
signal \il_max_comp2_D2\ : std_logic;
signal \phase_controller_slave.stoper_hc.N_60\ : std_logic;
signal \phase_controller_slave.hc_time_passed\ : std_logic;
signal \phase_controller_slave.state_RNIVDE2Z0Z_0\ : std_logic;
signal \phase_controller_slave.stateZ0Z_4\ : std_logic;
signal \phase_controller_slave.state_RNO_0Z0Z_3\ : std_logic;
signal shift_flag_start : std_logic;
signal \phase_controller_slave.stateZ0Z_1\ : std_logic;
signal s4_phy_c : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_7\ : std_logic;
signal \bfn_7_14_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_15\ : std_logic;
signal \bfn_7_15_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_23\ : std_logic;
signal \bfn_7_16_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_28\ : std_logic;
signal \bfn_7_17_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7\ : std_logic;
signal \bfn_7_18_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15\ : std_logic;
signal \bfn_7_19_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_startlt8_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_startlto5Z0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_startlto6Z0Z_0_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_startlt19_0_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_start\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_7_23_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ1Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_7_24_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_17\ : std_logic;
signal \bfn_7_25_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal il_max_comp1_c : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_105_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\ : std_logic;
signal \bfn_8_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\ : std_logic;
signal \bfn_8_14_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\ : std_logic;
signal \bfn_8_15_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\ : std_logic;
signal \bfn_8_16_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_178_i_g\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNI89DKZ0\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19\ : std_logic;
signal \phase_controller_slave.start_timer_hcZ0\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_startlto9_cZ0_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_startlto13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_8_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_start\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_startlto19Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_startlt15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJMZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\ : std_logic;
signal \bfn_8_25_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNI62NAZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\ : std_logic;
signal \bfn_8_26_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\ : std_logic;
signal \bfn_8_27_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_180_i\ : std_logic;
signal il_min_comp1_c : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_101\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_81_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_reset_1_i_a2_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_reset_1_i_a2_6_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_reset_1_i_a2_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_105\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_reset_1_i_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_reset_1_i_a2_9_cascade_\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_2\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_19\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_16\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_3\ : std_logic;
signal measured_delay_tr_8 : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg_5_0_o2_0_7_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg_5_0_o2_0_6_9_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg_5_0_o2_0_0_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_9_17_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ1Z_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_9_18_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_17\ : std_logic;
signal \bfn_9_19_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0\ : std_logic;
signal \il_min_comp1_D1\ : std_logic;
signal measured_delay_tr_15 : std_logic;
signal measured_delay_tr_6 : std_logic;
signal measured_delay_tr_12 : std_logic;
signal measured_delay_tr_14 : std_logic;
signal measured_delay_tr_1 : std_logic;
signal measured_delay_tr_17 : std_logic;
signal measured_delay_tr_9 : std_logic;
signal measured_delay_tr_5 : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_reset_i_a2_5_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_reset_i_a2_9_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_160_cascade_\ : std_logic;
signal \delay_measurement_inst.tr_state_RNIVV8GZ0Z_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_reset_i_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_2\ : std_logic;
signal measured_delay_tr_7 : std_logic;
signal measured_delay_tr_16 : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_slave.stateZ0Z_3\ : std_logic;
signal s3_phy_c : std_logic;
signal \delay_measurement_inst.N_54_cascade_\ : std_logic;
signal \delay_measurement_inst.tr_syncZ0Z_1\ : std_logic;
signal \delay_measurement_inst.tr_stateZ0Z_0\ : std_logic;
signal \delay_measurement_inst.tr_prevZ0\ : std_logic;
signal \delay_measurement_inst.hc_stateZ0Z_0\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_14\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_9\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_32\ : std_logic;
signal \delay_measurement_inst.N_54_i\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_8\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_1\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_10\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_4\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_18\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_17\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_6\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_13\ : std_logic;
signal \delay_measurement_inst.N_109\ : std_logic;
signal \delay_measurement_inst.N_45\ : std_logic;
signal \delay_measurement_inst.N_107\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_10_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_10_16_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_17\ : std_logic;
signal \bfn_10_17_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.stoper_state_RNI10KLZ0Z_1\ : std_logic;
signal measured_delay_tr_3 : std_logic;
signal measured_delay_tr_18 : std_logic;
signal measured_delay_tr_4 : std_logic;
signal \delay_measurement_inst.N_129\ : std_logic;
signal \delay_measurement_inst.N_172\ : std_logic;
signal measured_delay_tr_2 : std_logic;
signal measured_delay_tr_10 : std_logic;
signal measured_delay_tr_11 : std_logic;
signal measured_delay_tr_13 : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_reset_i_a2_6\ : std_logic;
signal \delay_measurement_inst.N_132\ : std_logic;
signal \delay_measurement_inst.N_139\ : std_logic;
signal \delay_measurement_inst.N_134_i\ : std_logic;
signal \delay_measurement_inst.N_201_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_167\ : std_logic;
signal \delay_measurement_inst.N_170\ : std_logic;
signal \il_min_comp1_D2\ : std_logic;
signal \phase_controller_inst1.T01_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_0\ : std_logic;
signal \T12_c\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.tr_time_passed\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_inst1.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_60\ : std_logic;
signal \delay_measurement_inst.stop_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.start_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_181_i\ : std_logic;
signal \delay_measurement_inst.hc_prevZ0\ : std_logic;
signal \delay_measurement_inst.hc_syncZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_81\ : std_logic;
signal \delay_measurement_inst.N_54\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlt8_cascade_\ : std_logic;
signal measured_delay_hc_8 : std_logic;
signal measured_delay_hc_7 : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto9_cZ0_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_8_cascade_\ : std_logic;
signal measured_delay_hc_1 : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_2\ : std_logic;
signal measured_delay_hc_5 : std_logic;
signal measured_delay_hc_16 : std_logic;
signal measured_delay_hc_19 : std_logic;
signal measured_delay_hc_17 : std_logic;
signal measured_delay_hc_18 : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_start\ : std_logic;
signal measured_delay_hc_6 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ1Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal measured_delay_hc_9 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal measured_delay_hc_13 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlt15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_start\ : std_logic;
signal measured_delay_hc_10 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal measured_delay_hc_14 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0_cascade_\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_1\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_2\ : std_logic;
signal \delay_measurement_inst.N_201\ : std_logic;
signal measured_delay_tr_19 : std_logic;
signal \delay_measurement_inst.N_134_i_0\ : std_logic;
signal \delay_measurement_inst.elapsed_time_ns_1_RNI6L42C_31\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_0_o2_0_7_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_reset_i_a2_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_127\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_0_o2_0_6_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_0_o2_0_0_9\ : std_logic;
signal clk_12mhz : std_logic;
signal \GB_BUFFER_clk_12mhz_THRU_CO\ : std_logic;
signal delay_hc_d2 : std_logic;
signal \delay_measurement_inst.hc_syncZ0Z_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_15\ : std_logic;
signal \delay_measurement_inst.N_84\ : std_logic;
signal \delay_measurement_inst.N_40\ : std_logic;
signal measured_delay_hc_15 : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_12\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_31\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_11\ : std_logic;
signal \delay_measurement_inst.N_48\ : std_logic;
signal \delay_measurement_inst.N_54_i_0\ : std_logic;
signal \delay_measurement_inst.N_32_g\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_179_i_g\ : std_logic;
signal measured_delay_hc_2 : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto6Z0Z_0\ : std_logic;
signal measured_delay_hc_3 : std_logic;
signal measured_delay_hc_4 : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_4\ : std_logic;
signal measured_delay_hc_12 : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlt19_0_cascade_\ : std_logic;
signal measured_delay_hc_11 : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_9\ : std_logic;
signal \il_max_comp1_D1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\ : std_logic;
signal \bfn_12_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIGEUBZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\ : std_logic;
signal \bfn_12_16_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\ : std_logic;
signal \bfn_12_17_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\ : std_logic;
signal \bfn_12_18_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_7\ : std_logic;
signal \bfn_12_19_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_15\ : std_logic;
signal \bfn_12_20_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_23\ : std_logic;
signal \bfn_12_21_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_181_i_g\ : std_logic;
signal \il_max_comp1_D2\ : std_logic;
signal \phase_controller_inst1.N_108\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_1\ : std_logic;
signal s2_phy_c : std_logic;
signal \phase_controller_inst1.stateZ0Z_3\ : std_logic;
signal s1_phy_c : std_logic;
signal \pll_inst.red_c_i\ : std_logic;
signal delay_hc_input_c : std_logic;
signal delay_hc_d1 : std_logic;
signal \delay_measurement_inst.tr_syncZ0Z_0\ : std_logic;
signal \delay_measurement_inst.start_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_178_i\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_state_RNITN7VZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_inst1.start_timer_hc_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.N_112\ : std_logic;
signal \phase_controller_inst1.start_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_3\ : std_logic;
signal \bfn_13_19_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_11\ : std_logic;
signal \bfn_13_20_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_19\ : std_logic;
signal \bfn_13_21_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\ : std_logic;
signal \bfn_13_22_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_31\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_180_i_g\ : std_logic;
signal start_stop_c : std_logic;
signal \phase_controller_inst1.stateZ0Z_4\ : std_logic;
signal \phase_controller_inst1.N_110\ : std_logic;
signal delay_tr_input_c : std_logic;
signal delay_tr_d1 : std_logic;
signal \T23_c\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_60\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst1.hc_time_passed\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_100mhz : std_logic;
signal red_c_g : std_logic;

signal reset_wire : std_logic;
signal il_min_comp2_wire : std_logic;
signal s1_phy_wire : std_logic;
signal s4_phy_wire : std_logic;
signal start_stop_wire : std_logic;
signal il_max_comp2_wire : std_logic;
signal \T23_wire\ : std_logic;
signal pwm_output_wire : std_logic;
signal il_max_comp1_wire : std_logic;
signal il_min_comp1_wire : std_logic;
signal s2_phy_wire : std_logic;
signal s3_phy_wire : std_logic;
signal delay_hc_input_wire : std_logic;
signal \T12_wire\ : std_logic;
signal delay_tr_input_wire : std_logic;
signal rgb_r_wire : std_logic;
signal rgb_b_wire : std_logic;
signal rgb_g_wire : std_logic;
signal \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    reset_wire <= reset;
    il_min_comp2_wire <= il_min_comp2;
    s1_phy <= s1_phy_wire;
    s4_phy <= s4_phy_wire;
    start_stop_wire <= start_stop;
    il_max_comp2_wire <= il_max_comp2;
    T23 <= \T23_wire\;
    pwm_output <= pwm_output_wire;
    il_max_comp1_wire <= il_max_comp1;
    il_min_comp1_wire <= il_min_comp1;
    s2_phy <= s2_phy_wire;
    s3_phy <= s3_phy_wire;
    delay_hc_input_wire <= delay_hc_input;
    T12 <= \T12_wire\;
    delay_tr_input_wire <= delay_tr_input;
    rgb_r <= rgb_r_wire;
    rgb_b <= rgb_b_wire;
    rgb_g <= rgb_g_wire;
    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__17066\,
            RESETB => \N__18890\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => clk_100mhz
        );

    \reset_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__21831\,
            GLOBALBUFFEROUTPUT => red_c_g
        );

    \reset_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21833\,
            DIN => \N__21832\,
            DOUT => \N__21831\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__21833\,
            PADOUT => \N__21832\,
            PADIN => \N__21831\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21822\,
            DIN => \N__21821\,
            DOUT => \N__21820\,
            PACKAGEPIN => il_min_comp2_wire
        );

    \il_min_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__21822\,
            PADOUT => \N__21821\,
            PADIN => \N__21820\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s1_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21813\,
            DIN => \N__21812\,
            DOUT => \N__21811\,
            PACKAGEPIN => s1_phy_wire
        );

    \s1_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__21813\,
            PADOUT => \N__21812\,
            PADIN => \N__21811\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__18902\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s4_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21804\,
            DIN => \N__21803\,
            DOUT => \N__21802\,
            PACKAGEPIN => s4_phy_wire
        );

    \s4_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__21804\,
            PADOUT => \N__21803\,
            PADIN => \N__21802\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9728\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \start_stop_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21795\,
            DIN => \N__21794\,
            DOUT => \N__21793\,
            PACKAGEPIN => start_stop_wire
        );

    \start_stop_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__21795\,
            PADOUT => \N__21794\,
            PADIN => \N__21793\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => start_stop_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21786\,
            DIN => \N__21785\,
            DOUT => \N__21784\,
            PACKAGEPIN => il_max_comp2_wire
        );

    \il_max_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__21786\,
            PADOUT => \N__21785\,
            PADIN => \N__21784\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T23_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21777\,
            DIN => \N__21776\,
            DOUT => \N__21775\,
            PACKAGEPIN => \T23_wire\
        );

    \T23_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__21777\,
            PADOUT => \N__21776\,
            PADIN => \N__21775\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21416\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21768\,
            DIN => \N__21767\,
            DOUT => \N__21766\,
            PACKAGEPIN => pwm_output_wire
        );

    \pwm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__21768\,
            PADOUT => \N__21767\,
            PADIN => \N__21766\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21759\,
            DIN => \N__21758\,
            DOUT => \N__21757\,
            PACKAGEPIN => il_max_comp1_wire
        );

    \il_max_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__21759\,
            PADOUT => \N__21758\,
            PADIN => \N__21757\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21750\,
            DIN => \N__21749\,
            DOUT => \N__21748\,
            PACKAGEPIN => il_min_comp1_wire
        );

    \il_min_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__21750\,
            PADOUT => \N__21749\,
            PADIN => \N__21748\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s2_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21741\,
            DIN => \N__21740\,
            DOUT => \N__21739\,
            PACKAGEPIN => s2_phy_wire
        );

    \s2_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__21741\,
            PADOUT => \N__21740\,
            PADIN => \N__21739\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__18950\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s3_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21732\,
            DIN => \N__21731\,
            DOUT => \N__21730\,
            PACKAGEPIN => s3_phy_wire
        );

    \s3_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__21732\,
            PADOUT => \N__21731\,
            PADIN => \N__21730\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__13892\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_hc_input_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21723\,
            DIN => \N__21722\,
            DOUT => \N__21721\,
            PACKAGEPIN => delay_hc_input_wire
        );

    \delay_hc_input_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__21723\,
            PADOUT => \N__21722\,
            PADIN => \N__21721\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_hc_input_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T12_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21714\,
            DIN => \N__21713\,
            DOUT => \N__21712\,
            PACKAGEPIN => \T12_wire\
        );

    \T12_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__21714\,
            PADOUT => \N__21713\,
            PADIN => \N__21712\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__15176\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_tr_input_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21705\,
            DIN => \N__21704\,
            DOUT => \N__21703\,
            PACKAGEPIN => delay_tr_input_wire
        );

    \delay_tr_input_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__21705\,
            PADOUT => \N__21704\,
            PADIN => \N__21703\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_tr_input_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__5172\ : InMux
    port map (
            O => \N__21686\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__5171\ : CascadeMux
    port map (
            O => \N__21683\,
            I => \N__21672\
        );

    \I__5170\ : InMux
    port map (
            O => \N__21682\,
            I => \N__21667\
        );

    \I__5169\ : InMux
    port map (
            O => \N__21681\,
            I => \N__21661\
        );

    \I__5168\ : InMux
    port map (
            O => \N__21680\,
            I => \N__21658\
        );

    \I__5167\ : InMux
    port map (
            O => \N__21679\,
            I => \N__21653\
        );

    \I__5166\ : InMux
    port map (
            O => \N__21678\,
            I => \N__21653\
        );

    \I__5165\ : InMux
    port map (
            O => \N__21677\,
            I => \N__21646\
        );

    \I__5164\ : InMux
    port map (
            O => \N__21676\,
            I => \N__21646\
        );

    \I__5163\ : InMux
    port map (
            O => \N__21675\,
            I => \N__21646\
        );

    \I__5162\ : InMux
    port map (
            O => \N__21672\,
            I => \N__21639\
        );

    \I__5161\ : InMux
    port map (
            O => \N__21671\,
            I => \N__21639\
        );

    \I__5160\ : InMux
    port map (
            O => \N__21670\,
            I => \N__21639\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__21667\,
            I => \N__21636\
        );

    \I__5158\ : InMux
    port map (
            O => \N__21666\,
            I => \N__21633\
        );

    \I__5157\ : InMux
    port map (
            O => \N__21665\,
            I => \N__21628\
        );

    \I__5156\ : InMux
    port map (
            O => \N__21664\,
            I => \N__21628\
        );

    \I__5155\ : LocalMux
    port map (
            O => \N__21661\,
            I => \N__21625\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__21658\,
            I => \N__21620\
        );

    \I__5153\ : LocalMux
    port map (
            O => \N__21653\,
            I => \N__21620\
        );

    \I__5152\ : LocalMux
    port map (
            O => \N__21646\,
            I => \N__21609\
        );

    \I__5151\ : LocalMux
    port map (
            O => \N__21639\,
            I => \N__21609\
        );

    \I__5150\ : Span4Mux_v
    port map (
            O => \N__21636\,
            I => \N__21609\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__21633\,
            I => \N__21609\
        );

    \I__5148\ : LocalMux
    port map (
            O => \N__21628\,
            I => \N__21609\
        );

    \I__5147\ : Span4Mux_h
    port map (
            O => \N__21625\,
            I => \N__21606\
        );

    \I__5146\ : Span4Mux_v
    port map (
            O => \N__21620\,
            I => \N__21601\
        );

    \I__5145\ : Span4Mux_v
    port map (
            O => \N__21609\,
            I => \N__21601\
        );

    \I__5144\ : Odrv4
    port map (
            O => \N__21606\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__5143\ : Odrv4
    port map (
            O => \N__21601\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__5142\ : CEMux
    port map (
            O => \N__21596\,
            I => \N__21581\
        );

    \I__5141\ : CEMux
    port map (
            O => \N__21595\,
            I => \N__21581\
        );

    \I__5140\ : CEMux
    port map (
            O => \N__21594\,
            I => \N__21581\
        );

    \I__5139\ : CEMux
    port map (
            O => \N__21593\,
            I => \N__21581\
        );

    \I__5138\ : CEMux
    port map (
            O => \N__21592\,
            I => \N__21581\
        );

    \I__5137\ : GlobalMux
    port map (
            O => \N__21581\,
            I => \N__21578\
        );

    \I__5136\ : gio2CtrlBuf
    port map (
            O => \N__21578\,
            I => \delay_measurement_inst.delay_tr_timer.N_180_i_g\
        );

    \I__5135\ : InMux
    port map (
            O => \N__21575\,
            I => \N__21572\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__21572\,
            I => \N__21568\
        );

    \I__5133\ : InMux
    port map (
            O => \N__21571\,
            I => \N__21565\
        );

    \I__5132\ : Span4Mux_s1_v
    port map (
            O => \N__21568\,
            I => \N__21560\
        );

    \I__5131\ : LocalMux
    port map (
            O => \N__21565\,
            I => \N__21560\
        );

    \I__5130\ : Span4Mux_v
    port map (
            O => \N__21560\,
            I => \N__21557\
        );

    \I__5129\ : Span4Mux_h
    port map (
            O => \N__21557\,
            I => \N__21551\
        );

    \I__5128\ : InMux
    port map (
            O => \N__21556\,
            I => \N__21548\
        );

    \I__5127\ : CascadeMux
    port map (
            O => \N__21555\,
            I => \N__21545\
        );

    \I__5126\ : InMux
    port map (
            O => \N__21554\,
            I => \N__21542\
        );

    \I__5125\ : Span4Mux_v
    port map (
            O => \N__21551\,
            I => \N__21537\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__21548\,
            I => \N__21537\
        );

    \I__5123\ : InMux
    port map (
            O => \N__21545\,
            I => \N__21534\
        );

    \I__5122\ : LocalMux
    port map (
            O => \N__21542\,
            I => \N__21531\
        );

    \I__5121\ : Span4Mux_v
    port map (
            O => \N__21537\,
            I => \N__21527\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__21534\,
            I => \N__21524\
        );

    \I__5119\ : Span4Mux_v
    port map (
            O => \N__21531\,
            I => \N__21521\
        );

    \I__5118\ : InMux
    port map (
            O => \N__21530\,
            I => \N__21518\
        );

    \I__5117\ : Sp12to4
    port map (
            O => \N__21527\,
            I => \N__21513\
        );

    \I__5116\ : Span12Mux_s6_h
    port map (
            O => \N__21524\,
            I => \N__21513\
        );

    \I__5115\ : Span4Mux_h
    port map (
            O => \N__21521\,
            I => \N__21510\
        );

    \I__5114\ : LocalMux
    port map (
            O => \N__21518\,
            I => \N__21507\
        );

    \I__5113\ : Span12Mux_v
    port map (
            O => \N__21513\,
            I => \N__21504\
        );

    \I__5112\ : Sp12to4
    port map (
            O => \N__21510\,
            I => \N__21499\
        );

    \I__5111\ : Span12Mux_h
    port map (
            O => \N__21507\,
            I => \N__21499\
        );

    \I__5110\ : Span12Mux_h
    port map (
            O => \N__21504\,
            I => \N__21496\
        );

    \I__5109\ : Span12Mux_v
    port map (
            O => \N__21499\,
            I => \N__21493\
        );

    \I__5108\ : Odrv12
    port map (
            O => \N__21496\,
            I => start_stop_c
        );

    \I__5107\ : Odrv12
    port map (
            O => \N__21493\,
            I => start_stop_c
        );

    \I__5106\ : CascadeMux
    port map (
            O => \N__21488\,
            I => \N__21484\
        );

    \I__5105\ : InMux
    port map (
            O => \N__21487\,
            I => \N__21481\
        );

    \I__5104\ : InMux
    port map (
            O => \N__21484\,
            I => \N__21477\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__21481\,
            I => \N__21474\
        );

    \I__5102\ : InMux
    port map (
            O => \N__21480\,
            I => \N__21471\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__21477\,
            I => \N__21468\
        );

    \I__5100\ : Span4Mux_v
    port map (
            O => \N__21474\,
            I => \N__21465\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__21471\,
            I => \N__21460\
        );

    \I__5098\ : Span4Mux_v
    port map (
            O => \N__21468\,
            I => \N__21455\
        );

    \I__5097\ : Span4Mux_h
    port map (
            O => \N__21465\,
            I => \N__21455\
        );

    \I__5096\ : InMux
    port map (
            O => \N__21464\,
            I => \N__21452\
        );

    \I__5095\ : InMux
    port map (
            O => \N__21463\,
            I => \N__21449\
        );

    \I__5094\ : Odrv12
    port map (
            O => \N__21460\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__5093\ : Odrv4
    port map (
            O => \N__21455\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__21452\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__21449\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__5090\ : InMux
    port map (
            O => \N__21440\,
            I => \N__21437\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__21437\,
            I => \phase_controller_inst1.N_110\
        );

    \I__5088\ : InMux
    port map (
            O => \N__21434\,
            I => \N__21431\
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__21431\,
            I => \N__21428\
        );

    \I__5086\ : Span4Mux_v
    port map (
            O => \N__21428\,
            I => \N__21425\
        );

    \I__5085\ : Odrv4
    port map (
            O => \N__21425\,
            I => delay_tr_input_c
        );

    \I__5084\ : InMux
    port map (
            O => \N__21422\,
            I => \N__21419\
        );

    \I__5083\ : LocalMux
    port map (
            O => \N__21419\,
            I => delay_tr_d1
        );

    \I__5082\ : IoInMux
    port map (
            O => \N__21416\,
            I => \N__21413\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__21413\,
            I => \N__21410\
        );

    \I__5080\ : Span4Mux_s3_v
    port map (
            O => \N__21410\,
            I => \N__21407\
        );

    \I__5079\ : Span4Mux_h
    port map (
            O => \N__21407\,
            I => \N__21404\
        );

    \I__5078\ : Sp12to4
    port map (
            O => \N__21404\,
            I => \N__21401\
        );

    \I__5077\ : Span12Mux_v
    port map (
            O => \N__21401\,
            I => \N__21397\
        );

    \I__5076\ : InMux
    port map (
            O => \N__21400\,
            I => \N__21394\
        );

    \I__5075\ : Odrv12
    port map (
            O => \N__21397\,
            I => \T23_c\
        );

    \I__5074\ : LocalMux
    port map (
            O => \N__21394\,
            I => \T23_c\
        );

    \I__5073\ : CascadeMux
    port map (
            O => \N__21389\,
            I => \N__21384\
        );

    \I__5072\ : CascadeMux
    port map (
            O => \N__21388\,
            I => \N__21381\
        );

    \I__5071\ : CascadeMux
    port map (
            O => \N__21387\,
            I => \N__21378\
        );

    \I__5070\ : InMux
    port map (
            O => \N__21384\,
            I => \N__21360\
        );

    \I__5069\ : InMux
    port map (
            O => \N__21381\,
            I => \N__21360\
        );

    \I__5068\ : InMux
    port map (
            O => \N__21378\,
            I => \N__21360\
        );

    \I__5067\ : InMux
    port map (
            O => \N__21377\,
            I => \N__21357\
        );

    \I__5066\ : InMux
    port map (
            O => \N__21376\,
            I => \N__21354\
        );

    \I__5065\ : InMux
    port map (
            O => \N__21375\,
            I => \N__21351\
        );

    \I__5064\ : CascadeMux
    port map (
            O => \N__21374\,
            I => \N__21340\
        );

    \I__5063\ : InMux
    port map (
            O => \N__21373\,
            I => \N__21323\
        );

    \I__5062\ : InMux
    port map (
            O => \N__21372\,
            I => \N__21323\
        );

    \I__5061\ : InMux
    port map (
            O => \N__21371\,
            I => \N__21323\
        );

    \I__5060\ : InMux
    port map (
            O => \N__21370\,
            I => \N__21323\
        );

    \I__5059\ : InMux
    port map (
            O => \N__21369\,
            I => \N__21323\
        );

    \I__5058\ : InMux
    port map (
            O => \N__21368\,
            I => \N__21323\
        );

    \I__5057\ : InMux
    port map (
            O => \N__21367\,
            I => \N__21323\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__21360\,
            I => \N__21318\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__21357\,
            I => \N__21318\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__21354\,
            I => \N__21313\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__21351\,
            I => \N__21313\
        );

    \I__5052\ : InMux
    port map (
            O => \N__21350\,
            I => \N__21300\
        );

    \I__5051\ : InMux
    port map (
            O => \N__21349\,
            I => \N__21300\
        );

    \I__5050\ : InMux
    port map (
            O => \N__21348\,
            I => \N__21300\
        );

    \I__5049\ : InMux
    port map (
            O => \N__21347\,
            I => \N__21300\
        );

    \I__5048\ : InMux
    port map (
            O => \N__21346\,
            I => \N__21300\
        );

    \I__5047\ : InMux
    port map (
            O => \N__21345\,
            I => \N__21287\
        );

    \I__5046\ : InMux
    port map (
            O => \N__21344\,
            I => \N__21287\
        );

    \I__5045\ : InMux
    port map (
            O => \N__21343\,
            I => \N__21287\
        );

    \I__5044\ : InMux
    port map (
            O => \N__21340\,
            I => \N__21287\
        );

    \I__5043\ : InMux
    port map (
            O => \N__21339\,
            I => \N__21287\
        );

    \I__5042\ : InMux
    port map (
            O => \N__21338\,
            I => \N__21287\
        );

    \I__5041\ : LocalMux
    port map (
            O => \N__21323\,
            I => \N__21282\
        );

    \I__5040\ : Span4Mux_h
    port map (
            O => \N__21318\,
            I => \N__21282\
        );

    \I__5039\ : Span4Mux_v
    port map (
            O => \N__21313\,
            I => \N__21279\
        );

    \I__5038\ : InMux
    port map (
            O => \N__21312\,
            I => \N__21274\
        );

    \I__5037\ : InMux
    port map (
            O => \N__21311\,
            I => \N__21274\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__21300\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__21287\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__5034\ : Odrv4
    port map (
            O => \N__21282\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__5033\ : Odrv4
    port map (
            O => \N__21279\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__21274\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__5031\ : CascadeMux
    port map (
            O => \N__21263\,
            I => \N__21260\
        );

    \I__5030\ : InMux
    port map (
            O => \N__21260\,
            I => \N__21257\
        );

    \I__5029\ : LocalMux
    port map (
            O => \N__21257\,
            I => \phase_controller_inst1.stoper_hc.N_60\
        );

    \I__5028\ : InMux
    port map (
            O => \N__21254\,
            I => \N__21251\
        );

    \I__5027\ : LocalMux
    port map (
            O => \N__21251\,
            I => \N__21243\
        );

    \I__5026\ : InMux
    port map (
            O => \N__21250\,
            I => \N__21232\
        );

    \I__5025\ : InMux
    port map (
            O => \N__21249\,
            I => \N__21232\
        );

    \I__5024\ : InMux
    port map (
            O => \N__21248\,
            I => \N__21232\
        );

    \I__5023\ : InMux
    port map (
            O => \N__21247\,
            I => \N__21232\
        );

    \I__5022\ : InMux
    port map (
            O => \N__21246\,
            I => \N__21232\
        );

    \I__5021\ : Odrv12
    port map (
            O => \N__21243\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__5020\ : LocalMux
    port map (
            O => \N__21232\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__5019\ : InMux
    port map (
            O => \N__21227\,
            I => \N__21223\
        );

    \I__5018\ : InMux
    port map (
            O => \N__21226\,
            I => \N__21220\
        );

    \I__5017\ : LocalMux
    port map (
            O => \N__21223\,
            I => \N__21215\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__21220\,
            I => \N__21215\
        );

    \I__5015\ : Span4Mux_h
    port map (
            O => \N__21215\,
            I => \N__21211\
        );

    \I__5014\ : InMux
    port map (
            O => \N__21214\,
            I => \N__21207\
        );

    \I__5013\ : Span4Mux_v
    port map (
            O => \N__21211\,
            I => \N__21204\
        );

    \I__5012\ : InMux
    port map (
            O => \N__21210\,
            I => \N__21201\
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__21207\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__5010\ : Odrv4
    port map (
            O => \N__21204\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__21201\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__5008\ : ClkMux
    port map (
            O => \N__21194\,
            I => \N__20906\
        );

    \I__5007\ : ClkMux
    port map (
            O => \N__21193\,
            I => \N__20906\
        );

    \I__5006\ : ClkMux
    port map (
            O => \N__21192\,
            I => \N__20906\
        );

    \I__5005\ : ClkMux
    port map (
            O => \N__21191\,
            I => \N__20906\
        );

    \I__5004\ : ClkMux
    port map (
            O => \N__21190\,
            I => \N__20906\
        );

    \I__5003\ : ClkMux
    port map (
            O => \N__21189\,
            I => \N__20906\
        );

    \I__5002\ : ClkMux
    port map (
            O => \N__21188\,
            I => \N__20906\
        );

    \I__5001\ : ClkMux
    port map (
            O => \N__21187\,
            I => \N__20906\
        );

    \I__5000\ : ClkMux
    port map (
            O => \N__21186\,
            I => \N__20906\
        );

    \I__4999\ : ClkMux
    port map (
            O => \N__21185\,
            I => \N__20906\
        );

    \I__4998\ : ClkMux
    port map (
            O => \N__21184\,
            I => \N__20906\
        );

    \I__4997\ : ClkMux
    port map (
            O => \N__21183\,
            I => \N__20906\
        );

    \I__4996\ : ClkMux
    port map (
            O => \N__21182\,
            I => \N__20906\
        );

    \I__4995\ : ClkMux
    port map (
            O => \N__21181\,
            I => \N__20906\
        );

    \I__4994\ : ClkMux
    port map (
            O => \N__21180\,
            I => \N__20906\
        );

    \I__4993\ : ClkMux
    port map (
            O => \N__21179\,
            I => \N__20906\
        );

    \I__4992\ : ClkMux
    port map (
            O => \N__21178\,
            I => \N__20906\
        );

    \I__4991\ : ClkMux
    port map (
            O => \N__21177\,
            I => \N__20906\
        );

    \I__4990\ : ClkMux
    port map (
            O => \N__21176\,
            I => \N__20906\
        );

    \I__4989\ : ClkMux
    port map (
            O => \N__21175\,
            I => \N__20906\
        );

    \I__4988\ : ClkMux
    port map (
            O => \N__21174\,
            I => \N__20906\
        );

    \I__4987\ : ClkMux
    port map (
            O => \N__21173\,
            I => \N__20906\
        );

    \I__4986\ : ClkMux
    port map (
            O => \N__21172\,
            I => \N__20906\
        );

    \I__4985\ : ClkMux
    port map (
            O => \N__21171\,
            I => \N__20906\
        );

    \I__4984\ : ClkMux
    port map (
            O => \N__21170\,
            I => \N__20906\
        );

    \I__4983\ : ClkMux
    port map (
            O => \N__21169\,
            I => \N__20906\
        );

    \I__4982\ : ClkMux
    port map (
            O => \N__21168\,
            I => \N__20906\
        );

    \I__4981\ : ClkMux
    port map (
            O => \N__21167\,
            I => \N__20906\
        );

    \I__4980\ : ClkMux
    port map (
            O => \N__21166\,
            I => \N__20906\
        );

    \I__4979\ : ClkMux
    port map (
            O => \N__21165\,
            I => \N__20906\
        );

    \I__4978\ : ClkMux
    port map (
            O => \N__21164\,
            I => \N__20906\
        );

    \I__4977\ : ClkMux
    port map (
            O => \N__21163\,
            I => \N__20906\
        );

    \I__4976\ : ClkMux
    port map (
            O => \N__21162\,
            I => \N__20906\
        );

    \I__4975\ : ClkMux
    port map (
            O => \N__21161\,
            I => \N__20906\
        );

    \I__4974\ : ClkMux
    port map (
            O => \N__21160\,
            I => \N__20906\
        );

    \I__4973\ : ClkMux
    port map (
            O => \N__21159\,
            I => \N__20906\
        );

    \I__4972\ : ClkMux
    port map (
            O => \N__21158\,
            I => \N__20906\
        );

    \I__4971\ : ClkMux
    port map (
            O => \N__21157\,
            I => \N__20906\
        );

    \I__4970\ : ClkMux
    port map (
            O => \N__21156\,
            I => \N__20906\
        );

    \I__4969\ : ClkMux
    port map (
            O => \N__21155\,
            I => \N__20906\
        );

    \I__4968\ : ClkMux
    port map (
            O => \N__21154\,
            I => \N__20906\
        );

    \I__4967\ : ClkMux
    port map (
            O => \N__21153\,
            I => \N__20906\
        );

    \I__4966\ : ClkMux
    port map (
            O => \N__21152\,
            I => \N__20906\
        );

    \I__4965\ : ClkMux
    port map (
            O => \N__21151\,
            I => \N__20906\
        );

    \I__4964\ : ClkMux
    port map (
            O => \N__21150\,
            I => \N__20906\
        );

    \I__4963\ : ClkMux
    port map (
            O => \N__21149\,
            I => \N__20906\
        );

    \I__4962\ : ClkMux
    port map (
            O => \N__21148\,
            I => \N__20906\
        );

    \I__4961\ : ClkMux
    port map (
            O => \N__21147\,
            I => \N__20906\
        );

    \I__4960\ : ClkMux
    port map (
            O => \N__21146\,
            I => \N__20906\
        );

    \I__4959\ : ClkMux
    port map (
            O => \N__21145\,
            I => \N__20906\
        );

    \I__4958\ : ClkMux
    port map (
            O => \N__21144\,
            I => \N__20906\
        );

    \I__4957\ : ClkMux
    port map (
            O => \N__21143\,
            I => \N__20906\
        );

    \I__4956\ : ClkMux
    port map (
            O => \N__21142\,
            I => \N__20906\
        );

    \I__4955\ : ClkMux
    port map (
            O => \N__21141\,
            I => \N__20906\
        );

    \I__4954\ : ClkMux
    port map (
            O => \N__21140\,
            I => \N__20906\
        );

    \I__4953\ : ClkMux
    port map (
            O => \N__21139\,
            I => \N__20906\
        );

    \I__4952\ : ClkMux
    port map (
            O => \N__21138\,
            I => \N__20906\
        );

    \I__4951\ : ClkMux
    port map (
            O => \N__21137\,
            I => \N__20906\
        );

    \I__4950\ : ClkMux
    port map (
            O => \N__21136\,
            I => \N__20906\
        );

    \I__4949\ : ClkMux
    port map (
            O => \N__21135\,
            I => \N__20906\
        );

    \I__4948\ : ClkMux
    port map (
            O => \N__21134\,
            I => \N__20906\
        );

    \I__4947\ : ClkMux
    port map (
            O => \N__21133\,
            I => \N__20906\
        );

    \I__4946\ : ClkMux
    port map (
            O => \N__21132\,
            I => \N__20906\
        );

    \I__4945\ : ClkMux
    port map (
            O => \N__21131\,
            I => \N__20906\
        );

    \I__4944\ : ClkMux
    port map (
            O => \N__21130\,
            I => \N__20906\
        );

    \I__4943\ : ClkMux
    port map (
            O => \N__21129\,
            I => \N__20906\
        );

    \I__4942\ : ClkMux
    port map (
            O => \N__21128\,
            I => \N__20906\
        );

    \I__4941\ : ClkMux
    port map (
            O => \N__21127\,
            I => \N__20906\
        );

    \I__4940\ : ClkMux
    port map (
            O => \N__21126\,
            I => \N__20906\
        );

    \I__4939\ : ClkMux
    port map (
            O => \N__21125\,
            I => \N__20906\
        );

    \I__4938\ : ClkMux
    port map (
            O => \N__21124\,
            I => \N__20906\
        );

    \I__4937\ : ClkMux
    port map (
            O => \N__21123\,
            I => \N__20906\
        );

    \I__4936\ : ClkMux
    port map (
            O => \N__21122\,
            I => \N__20906\
        );

    \I__4935\ : ClkMux
    port map (
            O => \N__21121\,
            I => \N__20906\
        );

    \I__4934\ : ClkMux
    port map (
            O => \N__21120\,
            I => \N__20906\
        );

    \I__4933\ : ClkMux
    port map (
            O => \N__21119\,
            I => \N__20906\
        );

    \I__4932\ : ClkMux
    port map (
            O => \N__21118\,
            I => \N__20906\
        );

    \I__4931\ : ClkMux
    port map (
            O => \N__21117\,
            I => \N__20906\
        );

    \I__4930\ : ClkMux
    port map (
            O => \N__21116\,
            I => \N__20906\
        );

    \I__4929\ : ClkMux
    port map (
            O => \N__21115\,
            I => \N__20906\
        );

    \I__4928\ : ClkMux
    port map (
            O => \N__21114\,
            I => \N__20906\
        );

    \I__4927\ : ClkMux
    port map (
            O => \N__21113\,
            I => \N__20906\
        );

    \I__4926\ : ClkMux
    port map (
            O => \N__21112\,
            I => \N__20906\
        );

    \I__4925\ : ClkMux
    port map (
            O => \N__21111\,
            I => \N__20906\
        );

    \I__4924\ : ClkMux
    port map (
            O => \N__21110\,
            I => \N__20906\
        );

    \I__4923\ : ClkMux
    port map (
            O => \N__21109\,
            I => \N__20906\
        );

    \I__4922\ : ClkMux
    port map (
            O => \N__21108\,
            I => \N__20906\
        );

    \I__4921\ : ClkMux
    port map (
            O => \N__21107\,
            I => \N__20906\
        );

    \I__4920\ : ClkMux
    port map (
            O => \N__21106\,
            I => \N__20906\
        );

    \I__4919\ : ClkMux
    port map (
            O => \N__21105\,
            I => \N__20906\
        );

    \I__4918\ : ClkMux
    port map (
            O => \N__21104\,
            I => \N__20906\
        );

    \I__4917\ : ClkMux
    port map (
            O => \N__21103\,
            I => \N__20906\
        );

    \I__4916\ : ClkMux
    port map (
            O => \N__21102\,
            I => \N__20906\
        );

    \I__4915\ : ClkMux
    port map (
            O => \N__21101\,
            I => \N__20906\
        );

    \I__4914\ : ClkMux
    port map (
            O => \N__21100\,
            I => \N__20906\
        );

    \I__4913\ : ClkMux
    port map (
            O => \N__21099\,
            I => \N__20906\
        );

    \I__4912\ : GlobalMux
    port map (
            O => \N__20906\,
            I => clk_100mhz
        );

    \I__4911\ : CascadeMux
    port map (
            O => \N__20903\,
            I => \N__20895\
        );

    \I__4910\ : InMux
    port map (
            O => \N__20902\,
            I => \N__20886\
        );

    \I__4909\ : InMux
    port map (
            O => \N__20901\,
            I => \N__20883\
        );

    \I__4908\ : InMux
    port map (
            O => \N__20900\,
            I => \N__20880\
        );

    \I__4907\ : InMux
    port map (
            O => \N__20899\,
            I => \N__20877\
        );

    \I__4906\ : InMux
    port map (
            O => \N__20898\,
            I => \N__20874\
        );

    \I__4905\ : InMux
    port map (
            O => \N__20895\,
            I => \N__20869\
        );

    \I__4904\ : InMux
    port map (
            O => \N__20894\,
            I => \N__20869\
        );

    \I__4903\ : InMux
    port map (
            O => \N__20893\,
            I => \N__20866\
        );

    \I__4902\ : InMux
    port map (
            O => \N__20892\,
            I => \N__20863\
        );

    \I__4901\ : InMux
    port map (
            O => \N__20891\,
            I => \N__20856\
        );

    \I__4900\ : InMux
    port map (
            O => \N__20890\,
            I => \N__20856\
        );

    \I__4899\ : InMux
    port map (
            O => \N__20889\,
            I => \N__20856\
        );

    \I__4898\ : LocalMux
    port map (
            O => \N__20886\,
            I => \N__20853\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__20883\,
            I => \N__20850\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__20880\,
            I => \N__20847\
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__20877\,
            I => \N__20840\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__20874\,
            I => \N__20815\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__20869\,
            I => \N__20773\
        );

    \I__4892\ : LocalMux
    port map (
            O => \N__20866\,
            I => \N__20770\
        );

    \I__4891\ : LocalMux
    port map (
            O => \N__20863\,
            I => \N__20766\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__20856\,
            I => \N__20763\
        );

    \I__4889\ : Glb2LocalMux
    port map (
            O => \N__20853\,
            I => \N__20597\
        );

    \I__4888\ : Glb2LocalMux
    port map (
            O => \N__20850\,
            I => \N__20597\
        );

    \I__4887\ : Glb2LocalMux
    port map (
            O => \N__20847\,
            I => \N__20597\
        );

    \I__4886\ : SRMux
    port map (
            O => \N__20846\,
            I => \N__20597\
        );

    \I__4885\ : SRMux
    port map (
            O => \N__20845\,
            I => \N__20597\
        );

    \I__4884\ : SRMux
    port map (
            O => \N__20844\,
            I => \N__20597\
        );

    \I__4883\ : SRMux
    port map (
            O => \N__20843\,
            I => \N__20597\
        );

    \I__4882\ : Glb2LocalMux
    port map (
            O => \N__20840\,
            I => \N__20597\
        );

    \I__4881\ : SRMux
    port map (
            O => \N__20839\,
            I => \N__20597\
        );

    \I__4880\ : SRMux
    port map (
            O => \N__20838\,
            I => \N__20597\
        );

    \I__4879\ : SRMux
    port map (
            O => \N__20837\,
            I => \N__20597\
        );

    \I__4878\ : SRMux
    port map (
            O => \N__20836\,
            I => \N__20597\
        );

    \I__4877\ : SRMux
    port map (
            O => \N__20835\,
            I => \N__20597\
        );

    \I__4876\ : SRMux
    port map (
            O => \N__20834\,
            I => \N__20597\
        );

    \I__4875\ : SRMux
    port map (
            O => \N__20833\,
            I => \N__20597\
        );

    \I__4874\ : SRMux
    port map (
            O => \N__20832\,
            I => \N__20597\
        );

    \I__4873\ : SRMux
    port map (
            O => \N__20831\,
            I => \N__20597\
        );

    \I__4872\ : SRMux
    port map (
            O => \N__20830\,
            I => \N__20597\
        );

    \I__4871\ : SRMux
    port map (
            O => \N__20829\,
            I => \N__20597\
        );

    \I__4870\ : SRMux
    port map (
            O => \N__20828\,
            I => \N__20597\
        );

    \I__4869\ : SRMux
    port map (
            O => \N__20827\,
            I => \N__20597\
        );

    \I__4868\ : SRMux
    port map (
            O => \N__20826\,
            I => \N__20597\
        );

    \I__4867\ : SRMux
    port map (
            O => \N__20825\,
            I => \N__20597\
        );

    \I__4866\ : SRMux
    port map (
            O => \N__20824\,
            I => \N__20597\
        );

    \I__4865\ : SRMux
    port map (
            O => \N__20823\,
            I => \N__20597\
        );

    \I__4864\ : SRMux
    port map (
            O => \N__20822\,
            I => \N__20597\
        );

    \I__4863\ : SRMux
    port map (
            O => \N__20821\,
            I => \N__20597\
        );

    \I__4862\ : SRMux
    port map (
            O => \N__20820\,
            I => \N__20597\
        );

    \I__4861\ : SRMux
    port map (
            O => \N__20819\,
            I => \N__20597\
        );

    \I__4860\ : SRMux
    port map (
            O => \N__20818\,
            I => \N__20597\
        );

    \I__4859\ : Glb2LocalMux
    port map (
            O => \N__20815\,
            I => \N__20597\
        );

    \I__4858\ : SRMux
    port map (
            O => \N__20814\,
            I => \N__20597\
        );

    \I__4857\ : SRMux
    port map (
            O => \N__20813\,
            I => \N__20597\
        );

    \I__4856\ : SRMux
    port map (
            O => \N__20812\,
            I => \N__20597\
        );

    \I__4855\ : SRMux
    port map (
            O => \N__20811\,
            I => \N__20597\
        );

    \I__4854\ : SRMux
    port map (
            O => \N__20810\,
            I => \N__20597\
        );

    \I__4853\ : SRMux
    port map (
            O => \N__20809\,
            I => \N__20597\
        );

    \I__4852\ : SRMux
    port map (
            O => \N__20808\,
            I => \N__20597\
        );

    \I__4851\ : SRMux
    port map (
            O => \N__20807\,
            I => \N__20597\
        );

    \I__4850\ : SRMux
    port map (
            O => \N__20806\,
            I => \N__20597\
        );

    \I__4849\ : SRMux
    port map (
            O => \N__20805\,
            I => \N__20597\
        );

    \I__4848\ : SRMux
    port map (
            O => \N__20804\,
            I => \N__20597\
        );

    \I__4847\ : SRMux
    port map (
            O => \N__20803\,
            I => \N__20597\
        );

    \I__4846\ : SRMux
    port map (
            O => \N__20802\,
            I => \N__20597\
        );

    \I__4845\ : SRMux
    port map (
            O => \N__20801\,
            I => \N__20597\
        );

    \I__4844\ : SRMux
    port map (
            O => \N__20800\,
            I => \N__20597\
        );

    \I__4843\ : SRMux
    port map (
            O => \N__20799\,
            I => \N__20597\
        );

    \I__4842\ : SRMux
    port map (
            O => \N__20798\,
            I => \N__20597\
        );

    \I__4841\ : SRMux
    port map (
            O => \N__20797\,
            I => \N__20597\
        );

    \I__4840\ : SRMux
    port map (
            O => \N__20796\,
            I => \N__20597\
        );

    \I__4839\ : SRMux
    port map (
            O => \N__20795\,
            I => \N__20597\
        );

    \I__4838\ : SRMux
    port map (
            O => \N__20794\,
            I => \N__20597\
        );

    \I__4837\ : SRMux
    port map (
            O => \N__20793\,
            I => \N__20597\
        );

    \I__4836\ : SRMux
    port map (
            O => \N__20792\,
            I => \N__20597\
        );

    \I__4835\ : SRMux
    port map (
            O => \N__20791\,
            I => \N__20597\
        );

    \I__4834\ : SRMux
    port map (
            O => \N__20790\,
            I => \N__20597\
        );

    \I__4833\ : SRMux
    port map (
            O => \N__20789\,
            I => \N__20597\
        );

    \I__4832\ : SRMux
    port map (
            O => \N__20788\,
            I => \N__20597\
        );

    \I__4831\ : SRMux
    port map (
            O => \N__20787\,
            I => \N__20597\
        );

    \I__4830\ : SRMux
    port map (
            O => \N__20786\,
            I => \N__20597\
        );

    \I__4829\ : SRMux
    port map (
            O => \N__20785\,
            I => \N__20597\
        );

    \I__4828\ : SRMux
    port map (
            O => \N__20784\,
            I => \N__20597\
        );

    \I__4827\ : SRMux
    port map (
            O => \N__20783\,
            I => \N__20597\
        );

    \I__4826\ : SRMux
    port map (
            O => \N__20782\,
            I => \N__20597\
        );

    \I__4825\ : SRMux
    port map (
            O => \N__20781\,
            I => \N__20597\
        );

    \I__4824\ : SRMux
    port map (
            O => \N__20780\,
            I => \N__20597\
        );

    \I__4823\ : SRMux
    port map (
            O => \N__20779\,
            I => \N__20597\
        );

    \I__4822\ : SRMux
    port map (
            O => \N__20778\,
            I => \N__20597\
        );

    \I__4821\ : SRMux
    port map (
            O => \N__20777\,
            I => \N__20597\
        );

    \I__4820\ : SRMux
    port map (
            O => \N__20776\,
            I => \N__20597\
        );

    \I__4819\ : Glb2LocalMux
    port map (
            O => \N__20773\,
            I => \N__20597\
        );

    \I__4818\ : Glb2LocalMux
    port map (
            O => \N__20770\,
            I => \N__20597\
        );

    \I__4817\ : SRMux
    port map (
            O => \N__20769\,
            I => \N__20597\
        );

    \I__4816\ : Glb2LocalMux
    port map (
            O => \N__20766\,
            I => \N__20597\
        );

    \I__4815\ : Glb2LocalMux
    port map (
            O => \N__20763\,
            I => \N__20597\
        );

    \I__4814\ : SRMux
    port map (
            O => \N__20762\,
            I => \N__20597\
        );

    \I__4813\ : SRMux
    port map (
            O => \N__20761\,
            I => \N__20597\
        );

    \I__4812\ : SRMux
    port map (
            O => \N__20760\,
            I => \N__20597\
        );

    \I__4811\ : SRMux
    port map (
            O => \N__20759\,
            I => \N__20597\
        );

    \I__4810\ : SRMux
    port map (
            O => \N__20758\,
            I => \N__20597\
        );

    \I__4809\ : GlobalMux
    port map (
            O => \N__20597\,
            I => \N__20594\
        );

    \I__4808\ : gio2CtrlBuf
    port map (
            O => \N__20594\,
            I => red_c_g
        );

    \I__4807\ : CascadeMux
    port map (
            O => \N__20591\,
            I => \N__20586\
        );

    \I__4806\ : InMux
    port map (
            O => \N__20590\,
            I => \N__20583\
        );

    \I__4805\ : InMux
    port map (
            O => \N__20589\,
            I => \N__20580\
        );

    \I__4804\ : InMux
    port map (
            O => \N__20586\,
            I => \N__20577\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__20583\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__4802\ : LocalMux
    port map (
            O => \N__20580\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__20577\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__4800\ : CascadeMux
    port map (
            O => \N__20570\,
            I => \N__20567\
        );

    \I__4799\ : InMux
    port map (
            O => \N__20567\,
            I => \N__20564\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__20564\,
            I => \N__20561\
        );

    \I__4797\ : Odrv4
    port map (
            O => \N__20561\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__4796\ : InMux
    port map (
            O => \N__20558\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__4795\ : CascadeMux
    port map (
            O => \N__20555\,
            I => \N__20550\
        );

    \I__4794\ : InMux
    port map (
            O => \N__20554\,
            I => \N__20547\
        );

    \I__4793\ : InMux
    port map (
            O => \N__20553\,
            I => \N__20544\
        );

    \I__4792\ : InMux
    port map (
            O => \N__20550\,
            I => \N__20541\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__20547\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__20544\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__20541\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__4788\ : InMux
    port map (
            O => \N__20534\,
            I => \N__20531\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__20531\,
            I => \N__20528\
        );

    \I__4786\ : Span4Mux_h
    port map (
            O => \N__20528\,
            I => \N__20525\
        );

    \I__4785\ : Odrv4
    port map (
            O => \N__20525\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__4784\ : InMux
    port map (
            O => \N__20522\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__4783\ : CascadeMux
    port map (
            O => \N__20519\,
            I => \N__20514\
        );

    \I__4782\ : InMux
    port map (
            O => \N__20518\,
            I => \N__20511\
        );

    \I__4781\ : InMux
    port map (
            O => \N__20517\,
            I => \N__20508\
        );

    \I__4780\ : InMux
    port map (
            O => \N__20514\,
            I => \N__20505\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__20511\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__4778\ : LocalMux
    port map (
            O => \N__20508\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__20505\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__4776\ : InMux
    port map (
            O => \N__20498\,
            I => \N__20495\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__20495\,
            I => \N__20492\
        );

    \I__4774\ : Odrv4
    port map (
            O => \N__20492\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__4773\ : InMux
    port map (
            O => \N__20489\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__4772\ : CascadeMux
    port map (
            O => \N__20486\,
            I => \N__20481\
        );

    \I__4771\ : InMux
    port map (
            O => \N__20485\,
            I => \N__20478\
        );

    \I__4770\ : InMux
    port map (
            O => \N__20484\,
            I => \N__20475\
        );

    \I__4769\ : InMux
    port map (
            O => \N__20481\,
            I => \N__20472\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__20478\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__20475\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__20472\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__4765\ : InMux
    port map (
            O => \N__20465\,
            I => \N__20462\
        );

    \I__4764\ : LocalMux
    port map (
            O => \N__20462\,
            I => \N__20459\
        );

    \I__4763\ : Odrv4
    port map (
            O => \N__20459\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__4762\ : InMux
    port map (
            O => \N__20456\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__4761\ : CascadeMux
    port map (
            O => \N__20453\,
            I => \N__20448\
        );

    \I__4760\ : InMux
    port map (
            O => \N__20452\,
            I => \N__20445\
        );

    \I__4759\ : InMux
    port map (
            O => \N__20451\,
            I => \N__20442\
        );

    \I__4758\ : InMux
    port map (
            O => \N__20448\,
            I => \N__20439\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__20445\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__4756\ : LocalMux
    port map (
            O => \N__20442\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__4755\ : LocalMux
    port map (
            O => \N__20439\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__4754\ : InMux
    port map (
            O => \N__20432\,
            I => \N__20429\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__20429\,
            I => \N__20426\
        );

    \I__4752\ : Span4Mux_v
    port map (
            O => \N__20426\,
            I => \N__20423\
        );

    \I__4751\ : Odrv4
    port map (
            O => \N__20423\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__4750\ : InMux
    port map (
            O => \N__20420\,
            I => \bfn_13_22_0_\
        );

    \I__4749\ : CascadeMux
    port map (
            O => \N__20417\,
            I => \N__20412\
        );

    \I__4748\ : InMux
    port map (
            O => \N__20416\,
            I => \N__20409\
        );

    \I__4747\ : InMux
    port map (
            O => \N__20415\,
            I => \N__20406\
        );

    \I__4746\ : InMux
    port map (
            O => \N__20412\,
            I => \N__20403\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__20409\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__20406\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__20403\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__4742\ : CascadeMux
    port map (
            O => \N__20396\,
            I => \N__20393\
        );

    \I__4741\ : InMux
    port map (
            O => \N__20393\,
            I => \N__20390\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__20390\,
            I => \N__20387\
        );

    \I__4739\ : Span4Mux_v
    port map (
            O => \N__20387\,
            I => \N__20384\
        );

    \I__4738\ : Odrv4
    port map (
            O => \N__20384\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__4737\ : InMux
    port map (
            O => \N__20381\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__4736\ : CascadeMux
    port map (
            O => \N__20378\,
            I => \N__20373\
        );

    \I__4735\ : InMux
    port map (
            O => \N__20377\,
            I => \N__20370\
        );

    \I__4734\ : InMux
    port map (
            O => \N__20376\,
            I => \N__20367\
        );

    \I__4733\ : InMux
    port map (
            O => \N__20373\,
            I => \N__20364\
        );

    \I__4732\ : LocalMux
    port map (
            O => \N__20370\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__4731\ : LocalMux
    port map (
            O => \N__20367\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__20364\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__4729\ : CascadeMux
    port map (
            O => \N__20357\,
            I => \N__20353\
        );

    \I__4728\ : InMux
    port map (
            O => \N__20356\,
            I => \N__20350\
        );

    \I__4727\ : InMux
    port map (
            O => \N__20353\,
            I => \N__20347\
        );

    \I__4726\ : LocalMux
    port map (
            O => \N__20350\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__20347\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__4724\ : InMux
    port map (
            O => \N__20342\,
            I => \N__20339\
        );

    \I__4723\ : LocalMux
    port map (
            O => \N__20339\,
            I => \N__20336\
        );

    \I__4722\ : Odrv4
    port map (
            O => \N__20336\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__4721\ : InMux
    port map (
            O => \N__20333\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__4720\ : CascadeMux
    port map (
            O => \N__20330\,
            I => \N__20325\
        );

    \I__4719\ : InMux
    port map (
            O => \N__20329\,
            I => \N__20322\
        );

    \I__4718\ : InMux
    port map (
            O => \N__20328\,
            I => \N__20319\
        );

    \I__4717\ : InMux
    port map (
            O => \N__20325\,
            I => \N__20316\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__20322\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__4715\ : LocalMux
    port map (
            O => \N__20319\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__20316\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__4713\ : CascadeMux
    port map (
            O => \N__20309\,
            I => \N__20305\
        );

    \I__4712\ : InMux
    port map (
            O => \N__20308\,
            I => \N__20302\
        );

    \I__4711\ : InMux
    port map (
            O => \N__20305\,
            I => \N__20299\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__20302\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__20299\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__4708\ : InMux
    port map (
            O => \N__20294\,
            I => \N__20291\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__20291\,
            I => \N__20288\
        );

    \I__4706\ : Odrv4
    port map (
            O => \N__20288\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\
        );

    \I__4705\ : InMux
    port map (
            O => \N__20285\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__4704\ : CascadeMux
    port map (
            O => \N__20282\,
            I => \N__20277\
        );

    \I__4703\ : InMux
    port map (
            O => \N__20281\,
            I => \N__20274\
        );

    \I__4702\ : InMux
    port map (
            O => \N__20280\,
            I => \N__20271\
        );

    \I__4701\ : InMux
    port map (
            O => \N__20277\,
            I => \N__20268\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__20274\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__20271\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__4698\ : LocalMux
    port map (
            O => \N__20268\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__4697\ : CascadeMux
    port map (
            O => \N__20261\,
            I => \N__20253\
        );

    \I__4696\ : InMux
    port map (
            O => \N__20260\,
            I => \N__20250\
        );

    \I__4695\ : InMux
    port map (
            O => \N__20259\,
            I => \N__20247\
        );

    \I__4694\ : InMux
    port map (
            O => \N__20258\,
            I => \N__20240\
        );

    \I__4693\ : InMux
    port map (
            O => \N__20257\,
            I => \N__20240\
        );

    \I__4692\ : InMux
    port map (
            O => \N__20256\,
            I => \N__20240\
        );

    \I__4691\ : InMux
    port map (
            O => \N__20253\,
            I => \N__20237\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__20250\,
            I => \N__20232\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__20247\,
            I => \N__20232\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__20240\,
            I => \N__20229\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__20237\,
            I => \N__20224\
        );

    \I__4686\ : Span4Mux_v
    port map (
            O => \N__20232\,
            I => \N__20224\
        );

    \I__4685\ : Span4Mux_v
    port map (
            O => \N__20229\,
            I => \N__20221\
        );

    \I__4684\ : Span4Mux_h
    port map (
            O => \N__20224\,
            I => \N__20218\
        );

    \I__4683\ : Odrv4
    port map (
            O => \N__20221\,
            I => \delay_measurement_inst.elapsed_time_tr_15\
        );

    \I__4682\ : Odrv4
    port map (
            O => \N__20218\,
            I => \delay_measurement_inst.elapsed_time_tr_15\
        );

    \I__4681\ : InMux
    port map (
            O => \N__20213\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__4680\ : CascadeMux
    port map (
            O => \N__20210\,
            I => \N__20205\
        );

    \I__4679\ : InMux
    port map (
            O => \N__20209\,
            I => \N__20202\
        );

    \I__4678\ : InMux
    port map (
            O => \N__20208\,
            I => \N__20199\
        );

    \I__4677\ : InMux
    port map (
            O => \N__20205\,
            I => \N__20196\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__20202\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__4675\ : LocalMux
    port map (
            O => \N__20199\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__20196\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__4673\ : InMux
    port map (
            O => \N__20189\,
            I => \N__20184\
        );

    \I__4672\ : InMux
    port map (
            O => \N__20188\,
            I => \N__20181\
        );

    \I__4671\ : InMux
    port map (
            O => \N__20187\,
            I => \N__20178\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__20184\,
            I => \N__20173\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__20181\,
            I => \N__20173\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__20178\,
            I => \N__20170\
        );

    \I__4667\ : Span4Mux_v
    port map (
            O => \N__20173\,
            I => \N__20167\
        );

    \I__4666\ : Span4Mux_v
    port map (
            O => \N__20170\,
            I => \N__20164\
        );

    \I__4665\ : Span4Mux_h
    port map (
            O => \N__20167\,
            I => \N__20161\
        );

    \I__4664\ : Odrv4
    port map (
            O => \N__20164\,
            I => \delay_measurement_inst.elapsed_time_tr_16\
        );

    \I__4663\ : Odrv4
    port map (
            O => \N__20161\,
            I => \delay_measurement_inst.elapsed_time_tr_16\
        );

    \I__4662\ : InMux
    port map (
            O => \N__20156\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__4661\ : CascadeMux
    port map (
            O => \N__20153\,
            I => \N__20148\
        );

    \I__4660\ : InMux
    port map (
            O => \N__20152\,
            I => \N__20145\
        );

    \I__4659\ : InMux
    port map (
            O => \N__20151\,
            I => \N__20142\
        );

    \I__4658\ : InMux
    port map (
            O => \N__20148\,
            I => \N__20139\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__20145\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__20142\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__4655\ : LocalMux
    port map (
            O => \N__20139\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__4654\ : InMux
    port map (
            O => \N__20132\,
            I => \N__20125\
        );

    \I__4653\ : InMux
    port map (
            O => \N__20131\,
            I => \N__20125\
        );

    \I__4652\ : InMux
    port map (
            O => \N__20130\,
            I => \N__20122\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__20125\,
            I => \N__20119\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__20122\,
            I => \N__20116\
        );

    \I__4649\ : Span4Mux_h
    port map (
            O => \N__20119\,
            I => \N__20113\
        );

    \I__4648\ : Odrv12
    port map (
            O => \N__20116\,
            I => \delay_measurement_inst.elapsed_time_tr_17\
        );

    \I__4647\ : Odrv4
    port map (
            O => \N__20113\,
            I => \delay_measurement_inst.elapsed_time_tr_17\
        );

    \I__4646\ : InMux
    port map (
            O => \N__20108\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__4645\ : CascadeMux
    port map (
            O => \N__20105\,
            I => \N__20100\
        );

    \I__4644\ : InMux
    port map (
            O => \N__20104\,
            I => \N__20097\
        );

    \I__4643\ : InMux
    port map (
            O => \N__20103\,
            I => \N__20094\
        );

    \I__4642\ : InMux
    port map (
            O => \N__20100\,
            I => \N__20091\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__20097\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__20094\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__20091\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__4638\ : CascadeMux
    port map (
            O => \N__20084\,
            I => \N__20080\
        );

    \I__4637\ : CascadeMux
    port map (
            O => \N__20083\,
            I => \N__20077\
        );

    \I__4636\ : InMux
    port map (
            O => \N__20080\,
            I => \N__20073\
        );

    \I__4635\ : InMux
    port map (
            O => \N__20077\,
            I => \N__20070\
        );

    \I__4634\ : InMux
    port map (
            O => \N__20076\,
            I => \N__20067\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__20073\,
            I => \N__20062\
        );

    \I__4632\ : LocalMux
    port map (
            O => \N__20070\,
            I => \N__20062\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__20067\,
            I => \N__20059\
        );

    \I__4630\ : Span4Mux_h
    port map (
            O => \N__20062\,
            I => \N__20056\
        );

    \I__4629\ : Odrv4
    port map (
            O => \N__20059\,
            I => \delay_measurement_inst.elapsed_time_tr_18\
        );

    \I__4628\ : Odrv4
    port map (
            O => \N__20056\,
            I => \delay_measurement_inst.elapsed_time_tr_18\
        );

    \I__4627\ : InMux
    port map (
            O => \N__20051\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__4626\ : CascadeMux
    port map (
            O => \N__20048\,
            I => \N__20043\
        );

    \I__4625\ : InMux
    port map (
            O => \N__20047\,
            I => \N__20040\
        );

    \I__4624\ : InMux
    port map (
            O => \N__20046\,
            I => \N__20037\
        );

    \I__4623\ : InMux
    port map (
            O => \N__20043\,
            I => \N__20034\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__20040\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__20037\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__20034\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__4619\ : InMux
    port map (
            O => \N__20027\,
            I => \N__20023\
        );

    \I__4618\ : CascadeMux
    port map (
            O => \N__20026\,
            I => \N__20019\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__20023\,
            I => \N__20016\
        );

    \I__4616\ : InMux
    port map (
            O => \N__20022\,
            I => \N__20011\
        );

    \I__4615\ : InMux
    port map (
            O => \N__20019\,
            I => \N__20011\
        );

    \I__4614\ : Span4Mux_v
    port map (
            O => \N__20016\,
            I => \N__20006\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__20011\,
            I => \N__20006\
        );

    \I__4612\ : Odrv4
    port map (
            O => \N__20006\,
            I => \delay_measurement_inst.elapsed_time_tr_19\
        );

    \I__4611\ : InMux
    port map (
            O => \N__20003\,
            I => \bfn_13_21_0_\
        );

    \I__4610\ : CascadeMux
    port map (
            O => \N__20000\,
            I => \N__19995\
        );

    \I__4609\ : InMux
    port map (
            O => \N__19999\,
            I => \N__19992\
        );

    \I__4608\ : InMux
    port map (
            O => \N__19998\,
            I => \N__19989\
        );

    \I__4607\ : InMux
    port map (
            O => \N__19995\,
            I => \N__19986\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__19992\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__19989\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__4604\ : LocalMux
    port map (
            O => \N__19986\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__4603\ : CascadeMux
    port map (
            O => \N__19979\,
            I => \N__19976\
        );

    \I__4602\ : InMux
    port map (
            O => \N__19976\,
            I => \N__19973\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__19973\,
            I => \N__19970\
        );

    \I__4600\ : Odrv12
    port map (
            O => \N__19970\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__4599\ : InMux
    port map (
            O => \N__19967\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__4598\ : CascadeMux
    port map (
            O => \N__19964\,
            I => \N__19959\
        );

    \I__4597\ : InMux
    port map (
            O => \N__19963\,
            I => \N__19956\
        );

    \I__4596\ : InMux
    port map (
            O => \N__19962\,
            I => \N__19953\
        );

    \I__4595\ : InMux
    port map (
            O => \N__19959\,
            I => \N__19950\
        );

    \I__4594\ : LocalMux
    port map (
            O => \N__19956\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__19953\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__19950\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__4591\ : InMux
    port map (
            O => \N__19943\,
            I => \N__19940\
        );

    \I__4590\ : LocalMux
    port map (
            O => \N__19940\,
            I => \N__19937\
        );

    \I__4589\ : Odrv4
    port map (
            O => \N__19937\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__4588\ : InMux
    port map (
            O => \N__19934\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__4587\ : CascadeMux
    port map (
            O => \N__19931\,
            I => \N__19926\
        );

    \I__4586\ : InMux
    port map (
            O => \N__19930\,
            I => \N__19923\
        );

    \I__4585\ : InMux
    port map (
            O => \N__19929\,
            I => \N__19920\
        );

    \I__4584\ : InMux
    port map (
            O => \N__19926\,
            I => \N__19917\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__19923\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__19920\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__19917\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__4580\ : InMux
    port map (
            O => \N__19910\,
            I => \N__19907\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__19907\,
            I => \N__19904\
        );

    \I__4578\ : Odrv12
    port map (
            O => \N__19904\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__4577\ : InMux
    port map (
            O => \N__19901\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__4576\ : CascadeMux
    port map (
            O => \N__19898\,
            I => \N__19895\
        );

    \I__4575\ : InMux
    port map (
            O => \N__19895\,
            I => \N__19892\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__19892\,
            I => \N__19888\
        );

    \I__4573\ : InMux
    port map (
            O => \N__19891\,
            I => \N__19885\
        );

    \I__4572\ : Span4Mux_h
    port map (
            O => \N__19888\,
            I => \N__19882\
        );

    \I__4571\ : LocalMux
    port map (
            O => \N__19885\,
            I => \N__19879\
        );

    \I__4570\ : Odrv4
    port map (
            O => \N__19882\,
            I => \delay_measurement_inst.elapsed_time_tr_7\
        );

    \I__4569\ : Odrv12
    port map (
            O => \N__19879\,
            I => \delay_measurement_inst.elapsed_time_tr_7\
        );

    \I__4568\ : InMux
    port map (
            O => \N__19874\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__4567\ : CascadeMux
    port map (
            O => \N__19871\,
            I => \N__19866\
        );

    \I__4566\ : InMux
    port map (
            O => \N__19870\,
            I => \N__19863\
        );

    \I__4565\ : InMux
    port map (
            O => \N__19869\,
            I => \N__19860\
        );

    \I__4564\ : InMux
    port map (
            O => \N__19866\,
            I => \N__19857\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__19863\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__19860\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__19857\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__4560\ : InMux
    port map (
            O => \N__19850\,
            I => \N__19847\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__19847\,
            I => \N__19844\
        );

    \I__4558\ : Span4Mux_h
    port map (
            O => \N__19844\,
            I => \N__19840\
        );

    \I__4557\ : InMux
    port map (
            O => \N__19843\,
            I => \N__19837\
        );

    \I__4556\ : Span4Mux_v
    port map (
            O => \N__19840\,
            I => \N__19834\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__19837\,
            I => \N__19831\
        );

    \I__4554\ : Odrv4
    port map (
            O => \N__19834\,
            I => \delay_measurement_inst.elapsed_time_tr_8\
        );

    \I__4553\ : Odrv12
    port map (
            O => \N__19831\,
            I => \delay_measurement_inst.elapsed_time_tr_8\
        );

    \I__4552\ : InMux
    port map (
            O => \N__19826\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__4551\ : CascadeMux
    port map (
            O => \N__19823\,
            I => \N__19818\
        );

    \I__4550\ : InMux
    port map (
            O => \N__19822\,
            I => \N__19815\
        );

    \I__4549\ : InMux
    port map (
            O => \N__19821\,
            I => \N__19812\
        );

    \I__4548\ : InMux
    port map (
            O => \N__19818\,
            I => \N__19809\
        );

    \I__4547\ : LocalMux
    port map (
            O => \N__19815\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__19812\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__19809\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__4544\ : InMux
    port map (
            O => \N__19802\,
            I => \N__19798\
        );

    \I__4543\ : CascadeMux
    port map (
            O => \N__19801\,
            I => \N__19794\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__19798\,
            I => \N__19791\
        );

    \I__4541\ : InMux
    port map (
            O => \N__19797\,
            I => \N__19788\
        );

    \I__4540\ : InMux
    port map (
            O => \N__19794\,
            I => \N__19785\
        );

    \I__4539\ : Span4Mux_v
    port map (
            O => \N__19791\,
            I => \N__19778\
        );

    \I__4538\ : LocalMux
    port map (
            O => \N__19788\,
            I => \N__19778\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__19785\,
            I => \N__19778\
        );

    \I__4536\ : Span4Mux_h
    port map (
            O => \N__19778\,
            I => \N__19775\
        );

    \I__4535\ : Odrv4
    port map (
            O => \N__19775\,
            I => \delay_measurement_inst.elapsed_time_tr_9\
        );

    \I__4534\ : InMux
    port map (
            O => \N__19772\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__4533\ : CascadeMux
    port map (
            O => \N__19769\,
            I => \N__19764\
        );

    \I__4532\ : InMux
    port map (
            O => \N__19768\,
            I => \N__19761\
        );

    \I__4531\ : InMux
    port map (
            O => \N__19767\,
            I => \N__19758\
        );

    \I__4530\ : InMux
    port map (
            O => \N__19764\,
            I => \N__19755\
        );

    \I__4529\ : LocalMux
    port map (
            O => \N__19761\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__19758\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__19755\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__4526\ : InMux
    port map (
            O => \N__19748\,
            I => \N__19745\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__19745\,
            I => \N__19741\
        );

    \I__4524\ : InMux
    port map (
            O => \N__19744\,
            I => \N__19738\
        );

    \I__4523\ : Span4Mux_v
    port map (
            O => \N__19741\,
            I => \N__19733\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__19738\,
            I => \N__19733\
        );

    \I__4521\ : Span4Mux_h
    port map (
            O => \N__19733\,
            I => \N__19730\
        );

    \I__4520\ : Odrv4
    port map (
            O => \N__19730\,
            I => \delay_measurement_inst.elapsed_time_tr_10\
        );

    \I__4519\ : InMux
    port map (
            O => \N__19727\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__4518\ : CascadeMux
    port map (
            O => \N__19724\,
            I => \N__19719\
        );

    \I__4517\ : InMux
    port map (
            O => \N__19723\,
            I => \N__19716\
        );

    \I__4516\ : InMux
    port map (
            O => \N__19722\,
            I => \N__19713\
        );

    \I__4515\ : InMux
    port map (
            O => \N__19719\,
            I => \N__19710\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__19716\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__19713\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__19710\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__4511\ : InMux
    port map (
            O => \N__19703\,
            I => \N__19699\
        );

    \I__4510\ : InMux
    port map (
            O => \N__19702\,
            I => \N__19696\
        );

    \I__4509\ : LocalMux
    port map (
            O => \N__19699\,
            I => \N__19693\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__19696\,
            I => \N__19690\
        );

    \I__4507\ : Span4Mux_h
    port map (
            O => \N__19693\,
            I => \N__19687\
        );

    \I__4506\ : Odrv12
    port map (
            O => \N__19690\,
            I => \delay_measurement_inst.elapsed_time_tr_11\
        );

    \I__4505\ : Odrv4
    port map (
            O => \N__19687\,
            I => \delay_measurement_inst.elapsed_time_tr_11\
        );

    \I__4504\ : InMux
    port map (
            O => \N__19682\,
            I => \bfn_13_20_0_\
        );

    \I__4503\ : CascadeMux
    port map (
            O => \N__19679\,
            I => \N__19674\
        );

    \I__4502\ : InMux
    port map (
            O => \N__19678\,
            I => \N__19671\
        );

    \I__4501\ : InMux
    port map (
            O => \N__19677\,
            I => \N__19668\
        );

    \I__4500\ : InMux
    port map (
            O => \N__19674\,
            I => \N__19665\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__19671\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__19668\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__19665\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__4496\ : InMux
    port map (
            O => \N__19658\,
            I => \N__19654\
        );

    \I__4495\ : InMux
    port map (
            O => \N__19657\,
            I => \N__19651\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__19654\,
            I => \N__19648\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__19651\,
            I => \N__19645\
        );

    \I__4492\ : Span4Mux_h
    port map (
            O => \N__19648\,
            I => \N__19642\
        );

    \I__4491\ : Odrv12
    port map (
            O => \N__19645\,
            I => \delay_measurement_inst.elapsed_time_tr_12\
        );

    \I__4490\ : Odrv4
    port map (
            O => \N__19642\,
            I => \delay_measurement_inst.elapsed_time_tr_12\
        );

    \I__4489\ : InMux
    port map (
            O => \N__19637\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__4488\ : CascadeMux
    port map (
            O => \N__19634\,
            I => \N__19629\
        );

    \I__4487\ : InMux
    port map (
            O => \N__19633\,
            I => \N__19626\
        );

    \I__4486\ : InMux
    port map (
            O => \N__19632\,
            I => \N__19623\
        );

    \I__4485\ : InMux
    port map (
            O => \N__19629\,
            I => \N__19620\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__19626\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__4483\ : LocalMux
    port map (
            O => \N__19623\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__19620\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__4481\ : CascadeMux
    port map (
            O => \N__19613\,
            I => \N__19609\
        );

    \I__4480\ : InMux
    port map (
            O => \N__19612\,
            I => \N__19606\
        );

    \I__4479\ : InMux
    port map (
            O => \N__19609\,
            I => \N__19603\
        );

    \I__4478\ : LocalMux
    port map (
            O => \N__19606\,
            I => \N__19600\
        );

    \I__4477\ : LocalMux
    port map (
            O => \N__19603\,
            I => \N__19597\
        );

    \I__4476\ : Span4Mux_h
    port map (
            O => \N__19600\,
            I => \N__19594\
        );

    \I__4475\ : Span4Mux_h
    port map (
            O => \N__19597\,
            I => \N__19591\
        );

    \I__4474\ : Odrv4
    port map (
            O => \N__19594\,
            I => \delay_measurement_inst.elapsed_time_tr_13\
        );

    \I__4473\ : Odrv4
    port map (
            O => \N__19591\,
            I => \delay_measurement_inst.elapsed_time_tr_13\
        );

    \I__4472\ : InMux
    port map (
            O => \N__19586\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__4471\ : CascadeMux
    port map (
            O => \N__19583\,
            I => \N__19578\
        );

    \I__4470\ : InMux
    port map (
            O => \N__19582\,
            I => \N__19575\
        );

    \I__4469\ : InMux
    port map (
            O => \N__19581\,
            I => \N__19572\
        );

    \I__4468\ : InMux
    port map (
            O => \N__19578\,
            I => \N__19569\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__19575\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__19572\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__19569\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__4464\ : CascadeMux
    port map (
            O => \N__19562\,
            I => \N__19559\
        );

    \I__4463\ : InMux
    port map (
            O => \N__19559\,
            I => \N__19553\
        );

    \I__4462\ : InMux
    port map (
            O => \N__19558\,
            I => \N__19548\
        );

    \I__4461\ : InMux
    port map (
            O => \N__19557\,
            I => \N__19548\
        );

    \I__4460\ : InMux
    port map (
            O => \N__19556\,
            I => \N__19545\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__19553\,
            I => \N__19540\
        );

    \I__4458\ : LocalMux
    port map (
            O => \N__19548\,
            I => \N__19540\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__19545\,
            I => \N__19537\
        );

    \I__4456\ : Span4Mux_h
    port map (
            O => \N__19540\,
            I => \N__19534\
        );

    \I__4455\ : Odrv12
    port map (
            O => \N__19537\,
            I => \delay_measurement_inst.elapsed_time_tr_14\
        );

    \I__4454\ : Odrv4
    port map (
            O => \N__19534\,
            I => \delay_measurement_inst.elapsed_time_tr_14\
        );

    \I__4453\ : InMux
    port map (
            O => \N__19529\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__4452\ : InMux
    port map (
            O => \N__19526\,
            I => \N__19523\
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__19523\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\
        );

    \I__4450\ : InMux
    port map (
            O => \N__19520\,
            I => \N__19516\
        );

    \I__4449\ : InMux
    port map (
            O => \N__19519\,
            I => \N__19513\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__19516\,
            I => \N__19510\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__19513\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__4446\ : Odrv4
    port map (
            O => \N__19510\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__4445\ : InMux
    port map (
            O => \N__19505\,
            I => \N__19501\
        );

    \I__4444\ : CascadeMux
    port map (
            O => \N__19504\,
            I => \N__19497\
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__19501\,
            I => \N__19494\
        );

    \I__4442\ : InMux
    port map (
            O => \N__19500\,
            I => \N__19491\
        );

    \I__4441\ : InMux
    port map (
            O => \N__19497\,
            I => \N__19488\
        );

    \I__4440\ : Span4Mux_v
    port map (
            O => \N__19494\,
            I => \N__19485\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__19491\,
            I => \N__19481\
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__19488\,
            I => \N__19476\
        );

    \I__4437\ : Span4Mux_h
    port map (
            O => \N__19485\,
            I => \N__19476\
        );

    \I__4436\ : InMux
    port map (
            O => \N__19484\,
            I => \N__19473\
        );

    \I__4435\ : Span4Mux_v
    port map (
            O => \N__19481\,
            I => \N__19470\
        );

    \I__4434\ : Odrv4
    port map (
            O => \N__19476\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__4433\ : LocalMux
    port map (
            O => \N__19473\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__4432\ : Odrv4
    port map (
            O => \N__19470\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__4431\ : CascadeMux
    port map (
            O => \N__19463\,
            I => \N__19452\
        );

    \I__4430\ : CascadeMux
    port map (
            O => \N__19462\,
            I => \N__19449\
        );

    \I__4429\ : CascadeMux
    port map (
            O => \N__19461\,
            I => \N__19446\
        );

    \I__4428\ : CascadeMux
    port map (
            O => \N__19460\,
            I => \N__19442\
        );

    \I__4427\ : InMux
    port map (
            O => \N__19459\,
            I => \N__19439\
        );

    \I__4426\ : InMux
    port map (
            O => \N__19458\,
            I => \N__19417\
        );

    \I__4425\ : InMux
    port map (
            O => \N__19457\,
            I => \N__19417\
        );

    \I__4424\ : InMux
    port map (
            O => \N__19456\,
            I => \N__19417\
        );

    \I__4423\ : InMux
    port map (
            O => \N__19455\,
            I => \N__19417\
        );

    \I__4422\ : InMux
    port map (
            O => \N__19452\,
            I => \N__19417\
        );

    \I__4421\ : InMux
    port map (
            O => \N__19449\,
            I => \N__19417\
        );

    \I__4420\ : InMux
    port map (
            O => \N__19446\,
            I => \N__19417\
        );

    \I__4419\ : InMux
    port map (
            O => \N__19445\,
            I => \N__19414\
        );

    \I__4418\ : InMux
    port map (
            O => \N__19442\,
            I => \N__19411\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__19439\,
            I => \N__19408\
        );

    \I__4416\ : CascadeMux
    port map (
            O => \N__19438\,
            I => \N__19404\
        );

    \I__4415\ : CascadeMux
    port map (
            O => \N__19437\,
            I => \N__19401\
        );

    \I__4414\ : CascadeMux
    port map (
            O => \N__19436\,
            I => \N__19398\
        );

    \I__4413\ : CascadeMux
    port map (
            O => \N__19435\,
            I => \N__19395\
        );

    \I__4412\ : CascadeMux
    port map (
            O => \N__19434\,
            I => \N__19389\
        );

    \I__4411\ : CascadeMux
    port map (
            O => \N__19433\,
            I => \N__19386\
        );

    \I__4410\ : CascadeMux
    port map (
            O => \N__19432\,
            I => \N__19383\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__19417\,
            I => \N__19378\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__19414\,
            I => \N__19375\
        );

    \I__4407\ : LocalMux
    port map (
            O => \N__19411\,
            I => \N__19370\
        );

    \I__4406\ : Span4Mux_v
    port map (
            O => \N__19408\,
            I => \N__19370\
        );

    \I__4405\ : InMux
    port map (
            O => \N__19407\,
            I => \N__19353\
        );

    \I__4404\ : InMux
    port map (
            O => \N__19404\,
            I => \N__19353\
        );

    \I__4403\ : InMux
    port map (
            O => \N__19401\,
            I => \N__19353\
        );

    \I__4402\ : InMux
    port map (
            O => \N__19398\,
            I => \N__19353\
        );

    \I__4401\ : InMux
    port map (
            O => \N__19395\,
            I => \N__19353\
        );

    \I__4400\ : InMux
    port map (
            O => \N__19394\,
            I => \N__19353\
        );

    \I__4399\ : InMux
    port map (
            O => \N__19393\,
            I => \N__19353\
        );

    \I__4398\ : InMux
    port map (
            O => \N__19392\,
            I => \N__19353\
        );

    \I__4397\ : InMux
    port map (
            O => \N__19389\,
            I => \N__19342\
        );

    \I__4396\ : InMux
    port map (
            O => \N__19386\,
            I => \N__19342\
        );

    \I__4395\ : InMux
    port map (
            O => \N__19383\,
            I => \N__19342\
        );

    \I__4394\ : InMux
    port map (
            O => \N__19382\,
            I => \N__19342\
        );

    \I__4393\ : InMux
    port map (
            O => \N__19381\,
            I => \N__19342\
        );

    \I__4392\ : Span4Mux_h
    port map (
            O => \N__19378\,
            I => \N__19339\
        );

    \I__4391\ : Span4Mux_v
    port map (
            O => \N__19375\,
            I => \N__19334\
        );

    \I__4390\ : Span4Mux_h
    port map (
            O => \N__19370\,
            I => \N__19334\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__19353\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__19342\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__4387\ : Odrv4
    port map (
            O => \N__19339\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__4386\ : Odrv4
    port map (
            O => \N__19334\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__4385\ : InMux
    port map (
            O => \N__19325\,
            I => \N__19322\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__19322\,
            I => \N__19319\
        );

    \I__4383\ : Span4Mux_v
    port map (
            O => \N__19319\,
            I => \N__19316\
        );

    \I__4382\ : Odrv4
    port map (
            O => \N__19316\,
            I => \phase_controller_inst1.start_timer_hc_0_sqmuxa\
        );

    \I__4381\ : InMux
    port map (
            O => \N__19313\,
            I => \N__19310\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__19310\,
            I => \phase_controller_inst1.N_112\
        );

    \I__4379\ : InMux
    port map (
            O => \N__19307\,
            I => \N__19286\
        );

    \I__4378\ : InMux
    port map (
            O => \N__19306\,
            I => \N__19286\
        );

    \I__4377\ : InMux
    port map (
            O => \N__19305\,
            I => \N__19286\
        );

    \I__4376\ : InMux
    port map (
            O => \N__19304\,
            I => \N__19286\
        );

    \I__4375\ : InMux
    port map (
            O => \N__19303\,
            I => \N__19286\
        );

    \I__4374\ : InMux
    port map (
            O => \N__19302\,
            I => \N__19286\
        );

    \I__4373\ : InMux
    port map (
            O => \N__19301\,
            I => \N__19286\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__19286\,
            I => \N__19269\
        );

    \I__4371\ : InMux
    port map (
            O => \N__19285\,
            I => \N__19260\
        );

    \I__4370\ : InMux
    port map (
            O => \N__19284\,
            I => \N__19260\
        );

    \I__4369\ : InMux
    port map (
            O => \N__19283\,
            I => \N__19260\
        );

    \I__4368\ : InMux
    port map (
            O => \N__19282\,
            I => \N__19260\
        );

    \I__4367\ : InMux
    port map (
            O => \N__19281\,
            I => \N__19257\
        );

    \I__4366\ : InMux
    port map (
            O => \N__19280\,
            I => \N__19240\
        );

    \I__4365\ : InMux
    port map (
            O => \N__19279\,
            I => \N__19240\
        );

    \I__4364\ : InMux
    port map (
            O => \N__19278\,
            I => \N__19240\
        );

    \I__4363\ : InMux
    port map (
            O => \N__19277\,
            I => \N__19240\
        );

    \I__4362\ : InMux
    port map (
            O => \N__19276\,
            I => \N__19240\
        );

    \I__4361\ : InMux
    port map (
            O => \N__19275\,
            I => \N__19240\
        );

    \I__4360\ : InMux
    port map (
            O => \N__19274\,
            I => \N__19240\
        );

    \I__4359\ : InMux
    port map (
            O => \N__19273\,
            I => \N__19240\
        );

    \I__4358\ : CascadeMux
    port map (
            O => \N__19272\,
            I => \N__19235\
        );

    \I__4357\ : Span4Mux_h
    port map (
            O => \N__19269\,
            I => \N__19232\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__19260\,
            I => \N__19227\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__19257\,
            I => \N__19227\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__19240\,
            I => \N__19224\
        );

    \I__4353\ : InMux
    port map (
            O => \N__19239\,
            I => \N__19220\
        );

    \I__4352\ : InMux
    port map (
            O => \N__19238\,
            I => \N__19217\
        );

    \I__4351\ : InMux
    port map (
            O => \N__19235\,
            I => \N__19214\
        );

    \I__4350\ : Span4Mux_v
    port map (
            O => \N__19232\,
            I => \N__19211\
        );

    \I__4349\ : Span4Mux_h
    port map (
            O => \N__19227\,
            I => \N__19208\
        );

    \I__4348\ : Span4Mux_h
    port map (
            O => \N__19224\,
            I => \N__19205\
        );

    \I__4347\ : InMux
    port map (
            O => \N__19223\,
            I => \N__19202\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__19220\,
            I => \N__19197\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__19217\,
            I => \N__19197\
        );

    \I__4344\ : LocalMux
    port map (
            O => \N__19214\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__4343\ : Odrv4
    port map (
            O => \N__19211\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__4342\ : Odrv4
    port map (
            O => \N__19208\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__4341\ : Odrv4
    port map (
            O => \N__19205\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__19202\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__4339\ : Odrv4
    port map (
            O => \N__19197\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__4338\ : InMux
    port map (
            O => \N__19184\,
            I => \N__19179\
        );

    \I__4337\ : InMux
    port map (
            O => \N__19183\,
            I => \N__19176\
        );

    \I__4336\ : InMux
    port map (
            O => \N__19182\,
            I => \N__19173\
        );

    \I__4335\ : LocalMux
    port map (
            O => \N__19179\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__19176\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__19173\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__4332\ : InMux
    port map (
            O => \N__19166\,
            I => \N__19162\
        );

    \I__4331\ : InMux
    port map (
            O => \N__19165\,
            I => \N__19159\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__19162\,
            I => \N__19156\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__19159\,
            I => \N__19153\
        );

    \I__4328\ : Span4Mux_h
    port map (
            O => \N__19156\,
            I => \N__19150\
        );

    \I__4327\ : Span4Mux_h
    port map (
            O => \N__19153\,
            I => \N__19147\
        );

    \I__4326\ : Odrv4
    port map (
            O => \N__19150\,
            I => \delay_measurement_inst.elapsed_time_tr_3\
        );

    \I__4325\ : Odrv4
    port map (
            O => \N__19147\,
            I => \delay_measurement_inst.elapsed_time_tr_3\
        );

    \I__4324\ : InMux
    port map (
            O => \N__19142\,
            I => \N__19137\
        );

    \I__4323\ : InMux
    port map (
            O => \N__19141\,
            I => \N__19134\
        );

    \I__4322\ : InMux
    port map (
            O => \N__19140\,
            I => \N__19131\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__19137\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__19134\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__19131\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__4318\ : CascadeMux
    port map (
            O => \N__19124\,
            I => \N__19121\
        );

    \I__4317\ : InMux
    port map (
            O => \N__19121\,
            I => \N__19117\
        );

    \I__4316\ : InMux
    port map (
            O => \N__19120\,
            I => \N__19114\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__19117\,
            I => \N__19111\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__19114\,
            I => \N__19108\
        );

    \I__4313\ : Span4Mux_h
    port map (
            O => \N__19111\,
            I => \N__19105\
        );

    \I__4312\ : Span4Mux_h
    port map (
            O => \N__19108\,
            I => \N__19102\
        );

    \I__4311\ : Odrv4
    port map (
            O => \N__19105\,
            I => \delay_measurement_inst.elapsed_time_tr_4\
        );

    \I__4310\ : Odrv4
    port map (
            O => \N__19102\,
            I => \delay_measurement_inst.elapsed_time_tr_4\
        );

    \I__4309\ : InMux
    port map (
            O => \N__19097\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__4308\ : CascadeMux
    port map (
            O => \N__19094\,
            I => \N__19089\
        );

    \I__4307\ : InMux
    port map (
            O => \N__19093\,
            I => \N__19086\
        );

    \I__4306\ : InMux
    port map (
            O => \N__19092\,
            I => \N__19083\
        );

    \I__4305\ : InMux
    port map (
            O => \N__19089\,
            I => \N__19080\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__19086\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__19083\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__4302\ : LocalMux
    port map (
            O => \N__19080\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__4301\ : InMux
    port map (
            O => \N__19073\,
            I => \N__19069\
        );

    \I__4300\ : InMux
    port map (
            O => \N__19072\,
            I => \N__19066\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__19069\,
            I => \N__19063\
        );

    \I__4298\ : LocalMux
    port map (
            O => \N__19066\,
            I => \N__19060\
        );

    \I__4297\ : Span4Mux_h
    port map (
            O => \N__19063\,
            I => \N__19057\
        );

    \I__4296\ : Span4Mux_v
    port map (
            O => \N__19060\,
            I => \N__19054\
        );

    \I__4295\ : Odrv4
    port map (
            O => \N__19057\,
            I => \delay_measurement_inst.elapsed_time_tr_5\
        );

    \I__4294\ : Odrv4
    port map (
            O => \N__19054\,
            I => \delay_measurement_inst.elapsed_time_tr_5\
        );

    \I__4293\ : InMux
    port map (
            O => \N__19049\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__4292\ : CascadeMux
    port map (
            O => \N__19046\,
            I => \N__19041\
        );

    \I__4291\ : InMux
    port map (
            O => \N__19045\,
            I => \N__19038\
        );

    \I__4290\ : InMux
    port map (
            O => \N__19044\,
            I => \N__19035\
        );

    \I__4289\ : InMux
    port map (
            O => \N__19041\,
            I => \N__19032\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__19038\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__4287\ : LocalMux
    port map (
            O => \N__19035\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__19032\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__4285\ : InMux
    port map (
            O => \N__19025\,
            I => \N__19022\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__19022\,
            I => \N__19018\
        );

    \I__4283\ : InMux
    port map (
            O => \N__19021\,
            I => \N__19015\
        );

    \I__4282\ : Span4Mux_h
    port map (
            O => \N__19018\,
            I => \N__19012\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__19015\,
            I => \N__19009\
        );

    \I__4280\ : Odrv4
    port map (
            O => \N__19012\,
            I => \delay_measurement_inst.elapsed_time_tr_6\
        );

    \I__4279\ : Odrv12
    port map (
            O => \N__19009\,
            I => \delay_measurement_inst.elapsed_time_tr_6\
        );

    \I__4278\ : InMux
    port map (
            O => \N__19004\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__4277\ : CascadeMux
    port map (
            O => \N__19001\,
            I => \N__18996\
        );

    \I__4276\ : InMux
    port map (
            O => \N__19000\,
            I => \N__18993\
        );

    \I__4275\ : InMux
    port map (
            O => \N__18999\,
            I => \N__18990\
        );

    \I__4274\ : InMux
    port map (
            O => \N__18996\,
            I => \N__18987\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__18993\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__18990\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__18987\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__4270\ : InMux
    port map (
            O => \N__18980\,
            I => \N__18977\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__18977\,
            I => \N__18973\
        );

    \I__4268\ : InMux
    port map (
            O => \N__18976\,
            I => \N__18970\
        );

    \I__4267\ : Span4Mux_h
    port map (
            O => \N__18973\,
            I => \N__18963\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__18970\,
            I => \N__18963\
        );

    \I__4265\ : InMux
    port map (
            O => \N__18969\,
            I => \N__18960\
        );

    \I__4264\ : InMux
    port map (
            O => \N__18968\,
            I => \N__18957\
        );

    \I__4263\ : Odrv4
    port map (
            O => \N__18963\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__18960\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__18957\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__4260\ : IoInMux
    port map (
            O => \N__18950\,
            I => \N__18947\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__18947\,
            I => \N__18944\
        );

    \I__4258\ : Span4Mux_s2_v
    port map (
            O => \N__18944\,
            I => \N__18941\
        );

    \I__4257\ : Odrv4
    port map (
            O => \N__18941\,
            I => s2_phy_c
        );

    \I__4256\ : InMux
    port map (
            O => \N__18938\,
            I => \N__18933\
        );

    \I__4255\ : CascadeMux
    port map (
            O => \N__18937\,
            I => \N__18930\
        );

    \I__4254\ : CascadeMux
    port map (
            O => \N__18936\,
            I => \N__18927\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__18933\,
            I => \N__18924\
        );

    \I__4252\ : InMux
    port map (
            O => \N__18930\,
            I => \N__18921\
        );

    \I__4251\ : InMux
    port map (
            O => \N__18927\,
            I => \N__18917\
        );

    \I__4250\ : Span4Mux_v
    port map (
            O => \N__18924\,
            I => \N__18912\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__18921\,
            I => \N__18912\
        );

    \I__4248\ : InMux
    port map (
            O => \N__18920\,
            I => \N__18909\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__18917\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__4246\ : Odrv4
    port map (
            O => \N__18912\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__18909\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__4244\ : IoInMux
    port map (
            O => \N__18902\,
            I => \N__18899\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__18899\,
            I => \N__18896\
        );

    \I__4242\ : Span4Mux_s1_v
    port map (
            O => \N__18896\,
            I => \N__18893\
        );

    \I__4241\ : Odrv4
    port map (
            O => \N__18893\,
            I => s1_phy_c
        );

    \I__4240\ : IoInMux
    port map (
            O => \N__18890\,
            I => \N__18887\
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__18887\,
            I => \N__18884\
        );

    \I__4238\ : Span4Mux_s0_v
    port map (
            O => \N__18884\,
            I => \N__18881\
        );

    \I__4237\ : Odrv4
    port map (
            O => \N__18881\,
            I => \pll_inst.red_c_i\
        );

    \I__4236\ : InMux
    port map (
            O => \N__18878\,
            I => \N__18875\
        );

    \I__4235\ : LocalMux
    port map (
            O => \N__18875\,
            I => \N__18872\
        );

    \I__4234\ : Span4Mux_h
    port map (
            O => \N__18872\,
            I => \N__18869\
        );

    \I__4233\ : Span4Mux_v
    port map (
            O => \N__18869\,
            I => \N__18866\
        );

    \I__4232\ : Odrv4
    port map (
            O => \N__18866\,
            I => delay_hc_input_c
        );

    \I__4231\ : InMux
    port map (
            O => \N__18863\,
            I => \N__18860\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__18860\,
            I => delay_hc_d1
        );

    \I__4229\ : InMux
    port map (
            O => \N__18857\,
            I => \N__18854\
        );

    \I__4228\ : LocalMux
    port map (
            O => \N__18854\,
            I => \N__18851\
        );

    \I__4227\ : Odrv12
    port map (
            O => \N__18851\,
            I => \delay_measurement_inst.tr_syncZ0Z_0\
        );

    \I__4226\ : InMux
    port map (
            O => \N__18848\,
            I => \N__18844\
        );

    \I__4225\ : InMux
    port map (
            O => \N__18847\,
            I => \N__18841\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__18844\,
            I => \N__18836\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__18841\,
            I => \N__18836\
        );

    \I__4222\ : Span4Mux_h
    port map (
            O => \N__18836\,
            I => \N__18833\
        );

    \I__4221\ : Odrv4
    port map (
            O => \N__18833\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__4220\ : InMux
    port map (
            O => \N__18830\,
            I => \N__18826\
        );

    \I__4219\ : InMux
    port map (
            O => \N__18829\,
            I => \N__18823\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__18826\,
            I => \N__18817\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__18823\,
            I => \N__18817\
        );

    \I__4216\ : InMux
    port map (
            O => \N__18822\,
            I => \N__18814\
        );

    \I__4215\ : Span4Mux_v
    port map (
            O => \N__18817\,
            I => \N__18811\
        );

    \I__4214\ : LocalMux
    port map (
            O => \N__18814\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__4213\ : Odrv4
    port map (
            O => \N__18811\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__4212\ : InMux
    port map (
            O => \N__18806\,
            I => \N__18800\
        );

    \I__4211\ : InMux
    port map (
            O => \N__18805\,
            I => \N__18795\
        );

    \I__4210\ : InMux
    port map (
            O => \N__18804\,
            I => \N__18795\
        );

    \I__4209\ : InMux
    port map (
            O => \N__18803\,
            I => \N__18792\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__18800\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__18795\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__18792\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__4205\ : IoInMux
    port map (
            O => \N__18785\,
            I => \N__18782\
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__18782\,
            I => \N__18779\
        );

    \I__4203\ : Span12Mux_s8_v
    port map (
            O => \N__18779\,
            I => \N__18776\
        );

    \I__4202\ : Odrv12
    port map (
            O => \N__18776\,
            I => \delay_measurement_inst.delay_hc_timer.N_178_i\
        );

    \I__4201\ : CEMux
    port map (
            O => \N__18773\,
            I => \N__18769\
        );

    \I__4200\ : CEMux
    port map (
            O => \N__18772\,
            I => \N__18766\
        );

    \I__4199\ : LocalMux
    port map (
            O => \N__18769\,
            I => \N__18762\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__18766\,
            I => \N__18759\
        );

    \I__4197\ : CEMux
    port map (
            O => \N__18765\,
            I => \N__18756\
        );

    \I__4196\ : Span4Mux_h
    port map (
            O => \N__18762\,
            I => \N__18753\
        );

    \I__4195\ : Span4Mux_h
    port map (
            O => \N__18759\,
            I => \N__18750\
        );

    \I__4194\ : LocalMux
    port map (
            O => \N__18756\,
            I => \N__18747\
        );

    \I__4193\ : Odrv4
    port map (
            O => \N__18753\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_RNITN7VZ0Z_1\
        );

    \I__4192\ : Odrv4
    port map (
            O => \N__18750\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_RNITN7VZ0Z_1\
        );

    \I__4191\ : Odrv12
    port map (
            O => \N__18747\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_RNITN7VZ0Z_1\
        );

    \I__4190\ : InMux
    port map (
            O => \N__18740\,
            I => \bfn_12_21_0_\
        );

    \I__4189\ : InMux
    port map (
            O => \N__18737\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_24\
        );

    \I__4188\ : InMux
    port map (
            O => \N__18734\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_25\
        );

    \I__4187\ : InMux
    port map (
            O => \N__18731\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_26\
        );

    \I__4186\ : InMux
    port map (
            O => \N__18728\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_27\
        );

    \I__4185\ : InMux
    port map (
            O => \N__18725\,
            I => \N__18687\
        );

    \I__4184\ : InMux
    port map (
            O => \N__18724\,
            I => \N__18687\
        );

    \I__4183\ : InMux
    port map (
            O => \N__18723\,
            I => \N__18687\
        );

    \I__4182\ : InMux
    port map (
            O => \N__18722\,
            I => \N__18687\
        );

    \I__4181\ : InMux
    port map (
            O => \N__18721\,
            I => \N__18678\
        );

    \I__4180\ : InMux
    port map (
            O => \N__18720\,
            I => \N__18678\
        );

    \I__4179\ : InMux
    port map (
            O => \N__18719\,
            I => \N__18678\
        );

    \I__4178\ : InMux
    port map (
            O => \N__18718\,
            I => \N__18678\
        );

    \I__4177\ : InMux
    port map (
            O => \N__18717\,
            I => \N__18669\
        );

    \I__4176\ : InMux
    port map (
            O => \N__18716\,
            I => \N__18669\
        );

    \I__4175\ : InMux
    port map (
            O => \N__18715\,
            I => \N__18669\
        );

    \I__4174\ : InMux
    port map (
            O => \N__18714\,
            I => \N__18669\
        );

    \I__4173\ : InMux
    port map (
            O => \N__18713\,
            I => \N__18664\
        );

    \I__4172\ : InMux
    port map (
            O => \N__18712\,
            I => \N__18664\
        );

    \I__4171\ : InMux
    port map (
            O => \N__18711\,
            I => \N__18655\
        );

    \I__4170\ : InMux
    port map (
            O => \N__18710\,
            I => \N__18655\
        );

    \I__4169\ : InMux
    port map (
            O => \N__18709\,
            I => \N__18655\
        );

    \I__4168\ : InMux
    port map (
            O => \N__18708\,
            I => \N__18655\
        );

    \I__4167\ : InMux
    port map (
            O => \N__18707\,
            I => \N__18646\
        );

    \I__4166\ : InMux
    port map (
            O => \N__18706\,
            I => \N__18646\
        );

    \I__4165\ : InMux
    port map (
            O => \N__18705\,
            I => \N__18646\
        );

    \I__4164\ : InMux
    port map (
            O => \N__18704\,
            I => \N__18646\
        );

    \I__4163\ : InMux
    port map (
            O => \N__18703\,
            I => \N__18637\
        );

    \I__4162\ : InMux
    port map (
            O => \N__18702\,
            I => \N__18637\
        );

    \I__4161\ : InMux
    port map (
            O => \N__18701\,
            I => \N__18637\
        );

    \I__4160\ : InMux
    port map (
            O => \N__18700\,
            I => \N__18637\
        );

    \I__4159\ : InMux
    port map (
            O => \N__18699\,
            I => \N__18628\
        );

    \I__4158\ : InMux
    port map (
            O => \N__18698\,
            I => \N__18628\
        );

    \I__4157\ : InMux
    port map (
            O => \N__18697\,
            I => \N__18628\
        );

    \I__4156\ : InMux
    port map (
            O => \N__18696\,
            I => \N__18628\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__18687\,
            I => \N__18621\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__18678\,
            I => \N__18621\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__18669\,
            I => \N__18621\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__18664\,
            I => \N__18610\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__18655\,
            I => \N__18610\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__18646\,
            I => \N__18610\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__18637\,
            I => \N__18610\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__18628\,
            I => \N__18610\
        );

    \I__4147\ : Span4Mux_v
    port map (
            O => \N__18621\,
            I => \N__18605\
        );

    \I__4146\ : Span4Mux_v
    port map (
            O => \N__18610\,
            I => \N__18605\
        );

    \I__4145\ : Span4Mux_v
    port map (
            O => \N__18605\,
            I => \N__18602\
        );

    \I__4144\ : Odrv4
    port map (
            O => \N__18602\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__4143\ : InMux
    port map (
            O => \N__18599\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_28\
        );

    \I__4142\ : CEMux
    port map (
            O => \N__18596\,
            I => \N__18584\
        );

    \I__4141\ : CEMux
    port map (
            O => \N__18595\,
            I => \N__18584\
        );

    \I__4140\ : CEMux
    port map (
            O => \N__18594\,
            I => \N__18584\
        );

    \I__4139\ : CEMux
    port map (
            O => \N__18593\,
            I => \N__18584\
        );

    \I__4138\ : GlobalMux
    port map (
            O => \N__18584\,
            I => \N__18581\
        );

    \I__4137\ : gio2CtrlBuf
    port map (
            O => \N__18581\,
            I => \delay_measurement_inst.delay_tr_timer.N_181_i_g\
        );

    \I__4136\ : InMux
    port map (
            O => \N__18578\,
            I => \N__18573\
        );

    \I__4135\ : InMux
    port map (
            O => \N__18577\,
            I => \N__18570\
        );

    \I__4134\ : InMux
    port map (
            O => \N__18576\,
            I => \N__18567\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__18573\,
            I => \N__18560\
        );

    \I__4132\ : LocalMux
    port map (
            O => \N__18570\,
            I => \N__18560\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__18567\,
            I => \N__18560\
        );

    \I__4130\ : Span12Mux_s11_v
    port map (
            O => \N__18560\,
            I => \N__18557\
        );

    \I__4129\ : Odrv12
    port map (
            O => \N__18557\,
            I => \il_max_comp1_D2\
        );

    \I__4128\ : InMux
    port map (
            O => \N__18554\,
            I => \N__18551\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__18551\,
            I => \N__18548\
        );

    \I__4126\ : Span4Mux_h
    port map (
            O => \N__18548\,
            I => \N__18544\
        );

    \I__4125\ : InMux
    port map (
            O => \N__18547\,
            I => \N__18541\
        );

    \I__4124\ : Odrv4
    port map (
            O => \N__18544\,
            I => \phase_controller_inst1.N_108\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__18541\,
            I => \phase_controller_inst1.N_108\
        );

    \I__4122\ : InMux
    port map (
            O => \N__18536\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_13\
        );

    \I__4121\ : InMux
    port map (
            O => \N__18533\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_14\
        );

    \I__4120\ : InMux
    port map (
            O => \N__18530\,
            I => \bfn_12_20_0_\
        );

    \I__4119\ : InMux
    port map (
            O => \N__18527\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_16\
        );

    \I__4118\ : InMux
    port map (
            O => \N__18524\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_17\
        );

    \I__4117\ : InMux
    port map (
            O => \N__18521\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_18\
        );

    \I__4116\ : InMux
    port map (
            O => \N__18518\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_19\
        );

    \I__4115\ : InMux
    port map (
            O => \N__18515\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_20\
        );

    \I__4114\ : InMux
    port map (
            O => \N__18512\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_21\
        );

    \I__4113\ : InMux
    port map (
            O => \N__18509\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_22\
        );

    \I__4112\ : InMux
    port map (
            O => \N__18506\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_4\
        );

    \I__4111\ : InMux
    port map (
            O => \N__18503\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_5\
        );

    \I__4110\ : InMux
    port map (
            O => \N__18500\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_6\
        );

    \I__4109\ : InMux
    port map (
            O => \N__18497\,
            I => \bfn_12_19_0_\
        );

    \I__4108\ : InMux
    port map (
            O => \N__18494\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_8\
        );

    \I__4107\ : InMux
    port map (
            O => \N__18491\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_9\
        );

    \I__4106\ : InMux
    port map (
            O => \N__18488\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_10\
        );

    \I__4105\ : InMux
    port map (
            O => \N__18485\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_11\
        );

    \I__4104\ : InMux
    port map (
            O => \N__18482\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_12\
        );

    \I__4103\ : InMux
    port map (
            O => \N__18479\,
            I => \N__18475\
        );

    \I__4102\ : InMux
    port map (
            O => \N__18478\,
            I => \N__18472\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__18475\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__18472\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__4099\ : InMux
    port map (
            O => \N__18467\,
            I => \N__18464\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__18464\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\
        );

    \I__4097\ : InMux
    port map (
            O => \N__18461\,
            I => \bfn_12_17_0_\
        );

    \I__4096\ : InMux
    port map (
            O => \N__18458\,
            I => \N__18454\
        );

    \I__4095\ : InMux
    port map (
            O => \N__18457\,
            I => \N__18451\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__18454\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__18451\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__4092\ : InMux
    port map (
            O => \N__18446\,
            I => \N__18443\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__18443\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\
        );

    \I__4090\ : InMux
    port map (
            O => \N__18440\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\
        );

    \I__4089\ : InMux
    port map (
            O => \N__18437\,
            I => \N__18433\
        );

    \I__4088\ : InMux
    port map (
            O => \N__18436\,
            I => \N__18430\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__18433\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__18430\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__4085\ : InMux
    port map (
            O => \N__18425\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\
        );

    \I__4084\ : InMux
    port map (
            O => \N__18422\,
            I => \N__18419\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__18419\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\
        );

    \I__4082\ : InMux
    port map (
            O => \N__18416\,
            I => \bfn_12_18_0_\
        );

    \I__4081\ : InMux
    port map (
            O => \N__18413\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_0\
        );

    \I__4080\ : InMux
    port map (
            O => \N__18410\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_1\
        );

    \I__4079\ : InMux
    port map (
            O => \N__18407\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_2\
        );

    \I__4078\ : InMux
    port map (
            O => \N__18404\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_3\
        );

    \I__4077\ : InMux
    port map (
            O => \N__18401\,
            I => \N__18397\
        );

    \I__4076\ : InMux
    port map (
            O => \N__18400\,
            I => \N__18394\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__18397\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__18394\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__4073\ : CascadeMux
    port map (
            O => \N__18389\,
            I => \N__18386\
        );

    \I__4072\ : InMux
    port map (
            O => \N__18386\,
            I => \N__18383\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__18383\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\
        );

    \I__4070\ : InMux
    port map (
            O => \N__18380\,
            I => \bfn_12_16_0_\
        );

    \I__4069\ : InMux
    port map (
            O => \N__18377\,
            I => \N__18373\
        );

    \I__4068\ : InMux
    port map (
            O => \N__18376\,
            I => \N__18370\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__18373\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__18370\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__4065\ : InMux
    port map (
            O => \N__18365\,
            I => \N__18362\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__18362\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\
        );

    \I__4063\ : InMux
    port map (
            O => \N__18359\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\
        );

    \I__4062\ : InMux
    port map (
            O => \N__18356\,
            I => \N__18352\
        );

    \I__4061\ : InMux
    port map (
            O => \N__18355\,
            I => \N__18349\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__18352\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__18349\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__4058\ : InMux
    port map (
            O => \N__18344\,
            I => \N__18341\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__18341\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\
        );

    \I__4056\ : InMux
    port map (
            O => \N__18338\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\
        );

    \I__4055\ : InMux
    port map (
            O => \N__18335\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\
        );

    \I__4054\ : InMux
    port map (
            O => \N__18332\,
            I => \N__18328\
        );

    \I__4053\ : InMux
    port map (
            O => \N__18331\,
            I => \N__18325\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__18328\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__18325\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__4050\ : InMux
    port map (
            O => \N__18320\,
            I => \N__18317\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__18317\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\
        );

    \I__4048\ : InMux
    port map (
            O => \N__18314\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\
        );

    \I__4047\ : InMux
    port map (
            O => \N__18311\,
            I => \N__18307\
        );

    \I__4046\ : InMux
    port map (
            O => \N__18310\,
            I => \N__18304\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__18307\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__18304\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__4043\ : InMux
    port map (
            O => \N__18299\,
            I => \N__18296\
        );

    \I__4042\ : LocalMux
    port map (
            O => \N__18296\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\
        );

    \I__4041\ : InMux
    port map (
            O => \N__18293\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\
        );

    \I__4040\ : InMux
    port map (
            O => \N__18290\,
            I => \N__18286\
        );

    \I__4039\ : InMux
    port map (
            O => \N__18289\,
            I => \N__18283\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__18286\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__18283\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__4036\ : InMux
    port map (
            O => \N__18278\,
            I => \N__18275\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__18275\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\
        );

    \I__4034\ : InMux
    port map (
            O => \N__18272\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\
        );

    \I__4033\ : InMux
    port map (
            O => \N__18269\,
            I => \N__18265\
        );

    \I__4032\ : InMux
    port map (
            O => \N__18268\,
            I => \N__18262\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__18265\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__18262\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__4029\ : InMux
    port map (
            O => \N__18257\,
            I => \N__18254\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__18254\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\
        );

    \I__4027\ : InMux
    port map (
            O => \N__18251\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\
        );

    \I__4026\ : InMux
    port map (
            O => \N__18248\,
            I => \N__18243\
        );

    \I__4025\ : InMux
    port map (
            O => \N__18247\,
            I => \N__18240\
        );

    \I__4024\ : InMux
    port map (
            O => \N__18246\,
            I => \N__18237\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__18243\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__18240\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__18237\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__4020\ : CascadeMux
    port map (
            O => \N__18230\,
            I => \N__18227\
        );

    \I__4019\ : InMux
    port map (
            O => \N__18227\,
            I => \N__18224\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__18224\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\
        );

    \I__4017\ : InMux
    port map (
            O => \N__18221\,
            I => \N__18217\
        );

    \I__4016\ : InMux
    port map (
            O => \N__18220\,
            I => \N__18214\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__18217\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__18214\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__4013\ : CascadeMux
    port map (
            O => \N__18209\,
            I => \N__18206\
        );

    \I__4012\ : InMux
    port map (
            O => \N__18206\,
            I => \N__18203\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__18203\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\
        );

    \I__4010\ : InMux
    port map (
            O => \N__18200\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\
        );

    \I__4009\ : InMux
    port map (
            O => \N__18197\,
            I => \N__18193\
        );

    \I__4008\ : InMux
    port map (
            O => \N__18196\,
            I => \N__18190\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__18193\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__18190\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__4005\ : CascadeMux
    port map (
            O => \N__18185\,
            I => \N__18182\
        );

    \I__4004\ : InMux
    port map (
            O => \N__18182\,
            I => \N__18179\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__18179\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIGEUBZ0\
        );

    \I__4002\ : CascadeMux
    port map (
            O => \N__18176\,
            I => \N__18173\
        );

    \I__4001\ : InMux
    port map (
            O => \N__18173\,
            I => \N__18170\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__18170\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\
        );

    \I__3999\ : InMux
    port map (
            O => \N__18167\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\
        );

    \I__3998\ : InMux
    port map (
            O => \N__18164\,
            I => \N__18160\
        );

    \I__3997\ : InMux
    port map (
            O => \N__18163\,
            I => \N__18157\
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__18160\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__18157\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__3994\ : InMux
    port map (
            O => \N__18152\,
            I => \N__18149\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__18149\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\
        );

    \I__3992\ : InMux
    port map (
            O => \N__18146\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\
        );

    \I__3991\ : CascadeMux
    port map (
            O => \N__18143\,
            I => \N__18140\
        );

    \I__3990\ : InMux
    port map (
            O => \N__18140\,
            I => \N__18136\
        );

    \I__3989\ : InMux
    port map (
            O => \N__18139\,
            I => \N__18133\
        );

    \I__3988\ : LocalMux
    port map (
            O => \N__18136\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__18133\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__3986\ : CascadeMux
    port map (
            O => \N__18128\,
            I => \N__18125\
        );

    \I__3985\ : InMux
    port map (
            O => \N__18125\,
            I => \N__18122\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__18122\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\
        );

    \I__3983\ : InMux
    port map (
            O => \N__18119\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\
        );

    \I__3982\ : CascadeMux
    port map (
            O => \N__18116\,
            I => \N__18113\
        );

    \I__3981\ : InMux
    port map (
            O => \N__18113\,
            I => \N__18109\
        );

    \I__3980\ : InMux
    port map (
            O => \N__18112\,
            I => \N__18106\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__18109\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__18106\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__3977\ : InMux
    port map (
            O => \N__18101\,
            I => \N__18098\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__18098\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\
        );

    \I__3975\ : InMux
    port map (
            O => \N__18095\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\
        );

    \I__3974\ : InMux
    port map (
            O => \N__18092\,
            I => \N__18088\
        );

    \I__3973\ : InMux
    port map (
            O => \N__18091\,
            I => \N__18085\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__18088\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__18085\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__3970\ : CascadeMux
    port map (
            O => \N__18080\,
            I => \N__18077\
        );

    \I__3969\ : InMux
    port map (
            O => \N__18077\,
            I => \N__18074\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__18074\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\
        );

    \I__3967\ : InMux
    port map (
            O => \N__18071\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\
        );

    \I__3966\ : CascadeMux
    port map (
            O => \N__18068\,
            I => \N__18065\
        );

    \I__3965\ : InMux
    port map (
            O => \N__18065\,
            I => \N__18061\
        );

    \I__3964\ : InMux
    port map (
            O => \N__18064\,
            I => \N__18058\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__18061\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__18058\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__3961\ : InMux
    port map (
            O => \N__18053\,
            I => \N__18050\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__18050\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\
        );

    \I__3959\ : InMux
    port map (
            O => \N__18047\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\
        );

    \I__3958\ : InMux
    port map (
            O => \N__18044\,
            I => \N__18041\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__18041\,
            I => \N__18035\
        );

    \I__3956\ : InMux
    port map (
            O => \N__18040\,
            I => \N__18032\
        );

    \I__3955\ : CascadeMux
    port map (
            O => \N__18039\,
            I => \N__18028\
        );

    \I__3954\ : CascadeMux
    port map (
            O => \N__18038\,
            I => \N__18025\
        );

    \I__3953\ : Span4Mux_h
    port map (
            O => \N__18035\,
            I => \N__18019\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__18032\,
            I => \N__18019\
        );

    \I__3951\ : InMux
    port map (
            O => \N__18031\,
            I => \N__18016\
        );

    \I__3950\ : InMux
    port map (
            O => \N__18028\,
            I => \N__18009\
        );

    \I__3949\ : InMux
    port map (
            O => \N__18025\,
            I => \N__18009\
        );

    \I__3948\ : InMux
    port map (
            O => \N__18024\,
            I => \N__18009\
        );

    \I__3947\ : Span4Mux_h
    port map (
            O => \N__18019\,
            I => \N__18006\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__18016\,
            I => \N__18001\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__18009\,
            I => \N__18001\
        );

    \I__3944\ : Odrv4
    port map (
            O => \N__18006\,
            I => \delay_measurement_inst.elapsed_time_hc_15\
        );

    \I__3943\ : Odrv4
    port map (
            O => \N__18001\,
            I => \delay_measurement_inst.elapsed_time_hc_15\
        );

    \I__3942\ : CascadeMux
    port map (
            O => \N__17996\,
            I => \N__17992\
        );

    \I__3941\ : CascadeMux
    port map (
            O => \N__17995\,
            I => \N__17989\
        );

    \I__3940\ : InMux
    port map (
            O => \N__17992\,
            I => \N__17986\
        );

    \I__3939\ : InMux
    port map (
            O => \N__17989\,
            I => \N__17983\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__17986\,
            I => \delay_measurement_inst.N_84\
        );

    \I__3937\ : LocalMux
    port map (
            O => \N__17983\,
            I => \delay_measurement_inst.N_84\
        );

    \I__3936\ : InMux
    port map (
            O => \N__17978\,
            I => \N__17975\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__17975\,
            I => \N__17969\
        );

    \I__3934\ : InMux
    port map (
            O => \N__17974\,
            I => \N__17966\
        );

    \I__3933\ : InMux
    port map (
            O => \N__17973\,
            I => \N__17955\
        );

    \I__3932\ : InMux
    port map (
            O => \N__17972\,
            I => \N__17955\
        );

    \I__3931\ : Span4Mux_v
    port map (
            O => \N__17969\,
            I => \N__17950\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__17966\,
            I => \N__17950\
        );

    \I__3929\ : InMux
    port map (
            O => \N__17965\,
            I => \N__17945\
        );

    \I__3928\ : InMux
    port map (
            O => \N__17964\,
            I => \N__17945\
        );

    \I__3927\ : InMux
    port map (
            O => \N__17963\,
            I => \N__17936\
        );

    \I__3926\ : InMux
    port map (
            O => \N__17962\,
            I => \N__17936\
        );

    \I__3925\ : InMux
    port map (
            O => \N__17961\,
            I => \N__17936\
        );

    \I__3924\ : InMux
    port map (
            O => \N__17960\,
            I => \N__17936\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__17955\,
            I => \N__17933\
        );

    \I__3922\ : Span4Mux_h
    port map (
            O => \N__17950\,
            I => \N__17926\
        );

    \I__3921\ : LocalMux
    port map (
            O => \N__17945\,
            I => \N__17926\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__17936\,
            I => \N__17926\
        );

    \I__3919\ : Odrv4
    port map (
            O => \N__17933\,
            I => \delay_measurement_inst.N_40\
        );

    \I__3918\ : Odrv4
    port map (
            O => \N__17926\,
            I => \delay_measurement_inst.N_40\
        );

    \I__3917\ : CascadeMux
    port map (
            O => \N__17921\,
            I => \N__17917\
        );

    \I__3916\ : InMux
    port map (
            O => \N__17920\,
            I => \N__17908\
        );

    \I__3915\ : InMux
    port map (
            O => \N__17917\,
            I => \N__17908\
        );

    \I__3914\ : InMux
    port map (
            O => \N__17916\,
            I => \N__17905\
        );

    \I__3913\ : InMux
    port map (
            O => \N__17915\,
            I => \N__17902\
        );

    \I__3912\ : InMux
    port map (
            O => \N__17914\,
            I => \N__17897\
        );

    \I__3911\ : InMux
    port map (
            O => \N__17913\,
            I => \N__17897\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__17908\,
            I => \N__17894\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__17905\,
            I => \N__17891\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__17902\,
            I => \N__17884\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__17897\,
            I => \N__17884\
        );

    \I__3906\ : Span4Mux_v
    port map (
            O => \N__17894\,
            I => \N__17884\
        );

    \I__3905\ : Span4Mux_h
    port map (
            O => \N__17891\,
            I => \N__17881\
        );

    \I__3904\ : Span4Mux_v
    port map (
            O => \N__17884\,
            I => \N__17875\
        );

    \I__3903\ : Span4Mux_v
    port map (
            O => \N__17881\,
            I => \N__17872\
        );

    \I__3902\ : InMux
    port map (
            O => \N__17880\,
            I => \N__17865\
        );

    \I__3901\ : InMux
    port map (
            O => \N__17879\,
            I => \N__17865\
        );

    \I__3900\ : InMux
    port map (
            O => \N__17878\,
            I => \N__17865\
        );

    \I__3899\ : Odrv4
    port map (
            O => \N__17875\,
            I => measured_delay_hc_15
        );

    \I__3898\ : Odrv4
    port map (
            O => \N__17872\,
            I => measured_delay_hc_15
        );

    \I__3897\ : LocalMux
    port map (
            O => \N__17865\,
            I => measured_delay_hc_15
        );

    \I__3896\ : InMux
    port map (
            O => \N__17858\,
            I => \N__17855\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__17855\,
            I => \N__17851\
        );

    \I__3894\ : InMux
    port map (
            O => \N__17854\,
            I => \N__17848\
        );

    \I__3893\ : Span4Mux_h
    port map (
            O => \N__17851\,
            I => \N__17845\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__17848\,
            I => \N__17842\
        );

    \I__3891\ : Odrv4
    port map (
            O => \N__17845\,
            I => \delay_measurement_inst.elapsed_time_hc_12\
        );

    \I__3890\ : Odrv4
    port map (
            O => \N__17842\,
            I => \delay_measurement_inst.elapsed_time_hc_12\
        );

    \I__3889\ : CascadeMux
    port map (
            O => \N__17837\,
            I => \N__17834\
        );

    \I__3888\ : InMux
    port map (
            O => \N__17834\,
            I => \N__17827\
        );

    \I__3887\ : InMux
    port map (
            O => \N__17833\,
            I => \N__17827\
        );

    \I__3886\ : CascadeMux
    port map (
            O => \N__17832\,
            I => \N__17822\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__17827\,
            I => \N__17815\
        );

    \I__3884\ : InMux
    port map (
            O => \N__17826\,
            I => \N__17806\
        );

    \I__3883\ : InMux
    port map (
            O => \N__17825\,
            I => \N__17806\
        );

    \I__3882\ : InMux
    port map (
            O => \N__17822\,
            I => \N__17806\
        );

    \I__3881\ : InMux
    port map (
            O => \N__17821\,
            I => \N__17806\
        );

    \I__3880\ : InMux
    port map (
            O => \N__17820\,
            I => \N__17799\
        );

    \I__3879\ : InMux
    port map (
            O => \N__17819\,
            I => \N__17799\
        );

    \I__3878\ : InMux
    port map (
            O => \N__17818\,
            I => \N__17799\
        );

    \I__3877\ : Span4Mux_v
    port map (
            O => \N__17815\,
            I => \N__17789\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__17806\,
            I => \N__17789\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__17799\,
            I => \N__17786\
        );

    \I__3874\ : InMux
    port map (
            O => \N__17798\,
            I => \N__17783\
        );

    \I__3873\ : InMux
    port map (
            O => \N__17797\,
            I => \N__17780\
        );

    \I__3872\ : InMux
    port map (
            O => \N__17796\,
            I => \N__17775\
        );

    \I__3871\ : InMux
    port map (
            O => \N__17795\,
            I => \N__17775\
        );

    \I__3870\ : InMux
    port map (
            O => \N__17794\,
            I => \N__17772\
        );

    \I__3869\ : Span4Mux_v
    port map (
            O => \N__17789\,
            I => \N__17769\
        );

    \I__3868\ : Span4Mux_h
    port map (
            O => \N__17786\,
            I => \N__17762\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__17783\,
            I => \N__17762\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__17780\,
            I => \N__17762\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__17775\,
            I => \N__17759\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__17772\,
            I => \N__17756\
        );

    \I__3863\ : Span4Mux_h
    port map (
            O => \N__17769\,
            I => \N__17753\
        );

    \I__3862\ : Span4Mux_h
    port map (
            O => \N__17762\,
            I => \N__17750\
        );

    \I__3861\ : Span4Mux_v
    port map (
            O => \N__17759\,
            I => \N__17745\
        );

    \I__3860\ : Span4Mux_v
    port map (
            O => \N__17756\,
            I => \N__17745\
        );

    \I__3859\ : Odrv4
    port map (
            O => \N__17753\,
            I => \delay_measurement_inst.elapsed_time_hc_31\
        );

    \I__3858\ : Odrv4
    port map (
            O => \N__17750\,
            I => \delay_measurement_inst.elapsed_time_hc_31\
        );

    \I__3857\ : Odrv4
    port map (
            O => \N__17745\,
            I => \delay_measurement_inst.elapsed_time_hc_31\
        );

    \I__3856\ : InMux
    port map (
            O => \N__17738\,
            I => \N__17735\
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__17735\,
            I => \N__17731\
        );

    \I__3854\ : InMux
    port map (
            O => \N__17734\,
            I => \N__17728\
        );

    \I__3853\ : Span4Mux_h
    port map (
            O => \N__17731\,
            I => \N__17725\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__17728\,
            I => \N__17722\
        );

    \I__3851\ : Odrv4
    port map (
            O => \N__17725\,
            I => \delay_measurement_inst.elapsed_time_hc_11\
        );

    \I__3850\ : Odrv4
    port map (
            O => \N__17722\,
            I => \delay_measurement_inst.elapsed_time_hc_11\
        );

    \I__3849\ : InMux
    port map (
            O => \N__17717\,
            I => \N__17711\
        );

    \I__3848\ : InMux
    port map (
            O => \N__17716\,
            I => \N__17711\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__17711\,
            I => \N__17705\
        );

    \I__3846\ : InMux
    port map (
            O => \N__17710\,
            I => \N__17702\
        );

    \I__3845\ : InMux
    port map (
            O => \N__17709\,
            I => \N__17697\
        );

    \I__3844\ : InMux
    port map (
            O => \N__17708\,
            I => \N__17697\
        );

    \I__3843\ : Odrv4
    port map (
            O => \N__17705\,
            I => \delay_measurement_inst.N_48\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__17702\,
            I => \delay_measurement_inst.N_48\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__17697\,
            I => \delay_measurement_inst.N_48\
        );

    \I__3840\ : CEMux
    port map (
            O => \N__17690\,
            I => \N__17687\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__17687\,
            I => \N__17683\
        );

    \I__3838\ : CEMux
    port map (
            O => \N__17686\,
            I => \N__17678\
        );

    \I__3837\ : Span4Mux_h
    port map (
            O => \N__17683\,
            I => \N__17675\
        );

    \I__3836\ : CEMux
    port map (
            O => \N__17682\,
            I => \N__17672\
        );

    \I__3835\ : CEMux
    port map (
            O => \N__17681\,
            I => \N__17669\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__17678\,
            I => \delay_measurement_inst.N_54_i_0\
        );

    \I__3833\ : Odrv4
    port map (
            O => \N__17675\,
            I => \delay_measurement_inst.N_54_i_0\
        );

    \I__3832\ : LocalMux
    port map (
            O => \N__17672\,
            I => \delay_measurement_inst.N_54_i_0\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__17669\,
            I => \delay_measurement_inst.N_54_i_0\
        );

    \I__3830\ : SRMux
    port map (
            O => \N__17660\,
            I => \N__17645\
        );

    \I__3829\ : SRMux
    port map (
            O => \N__17659\,
            I => \N__17645\
        );

    \I__3828\ : SRMux
    port map (
            O => \N__17658\,
            I => \N__17645\
        );

    \I__3827\ : SRMux
    port map (
            O => \N__17657\,
            I => \N__17645\
        );

    \I__3826\ : SRMux
    port map (
            O => \N__17656\,
            I => \N__17645\
        );

    \I__3825\ : GlobalMux
    port map (
            O => \N__17645\,
            I => \N__17642\
        );

    \I__3824\ : gio2CtrlBuf
    port map (
            O => \N__17642\,
            I => \delay_measurement_inst.N_32_g\
        );

    \I__3823\ : InMux
    port map (
            O => \N__17639\,
            I => \N__17627\
        );

    \I__3822\ : InMux
    port map (
            O => \N__17638\,
            I => \N__17627\
        );

    \I__3821\ : InMux
    port map (
            O => \N__17637\,
            I => \N__17627\
        );

    \I__3820\ : InMux
    port map (
            O => \N__17636\,
            I => \N__17627\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__17627\,
            I => \N__17614\
        );

    \I__3818\ : InMux
    port map (
            O => \N__17626\,
            I => \N__17609\
        );

    \I__3817\ : InMux
    port map (
            O => \N__17625\,
            I => \N__17609\
        );

    \I__3816\ : InMux
    port map (
            O => \N__17624\,
            I => \N__17600\
        );

    \I__3815\ : InMux
    port map (
            O => \N__17623\,
            I => \N__17600\
        );

    \I__3814\ : InMux
    port map (
            O => \N__17622\,
            I => \N__17600\
        );

    \I__3813\ : InMux
    port map (
            O => \N__17621\,
            I => \N__17600\
        );

    \I__3812\ : InMux
    port map (
            O => \N__17620\,
            I => \N__17591\
        );

    \I__3811\ : InMux
    port map (
            O => \N__17619\,
            I => \N__17591\
        );

    \I__3810\ : InMux
    port map (
            O => \N__17618\,
            I => \N__17591\
        );

    \I__3809\ : InMux
    port map (
            O => \N__17617\,
            I => \N__17591\
        );

    \I__3808\ : Span4Mux_v
    port map (
            O => \N__17614\,
            I => \N__17578\
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__17609\,
            I => \N__17578\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__17600\,
            I => \N__17578\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__17591\,
            I => \N__17578\
        );

    \I__3804\ : InMux
    port map (
            O => \N__17590\,
            I => \N__17561\
        );

    \I__3803\ : InMux
    port map (
            O => \N__17589\,
            I => \N__17561\
        );

    \I__3802\ : InMux
    port map (
            O => \N__17588\,
            I => \N__17561\
        );

    \I__3801\ : InMux
    port map (
            O => \N__17587\,
            I => \N__17561\
        );

    \I__3800\ : Span4Mux_v
    port map (
            O => \N__17578\,
            I => \N__17558\
        );

    \I__3799\ : InMux
    port map (
            O => \N__17577\,
            I => \N__17549\
        );

    \I__3798\ : InMux
    port map (
            O => \N__17576\,
            I => \N__17549\
        );

    \I__3797\ : InMux
    port map (
            O => \N__17575\,
            I => \N__17549\
        );

    \I__3796\ : InMux
    port map (
            O => \N__17574\,
            I => \N__17549\
        );

    \I__3795\ : InMux
    port map (
            O => \N__17573\,
            I => \N__17540\
        );

    \I__3794\ : InMux
    port map (
            O => \N__17572\,
            I => \N__17540\
        );

    \I__3793\ : InMux
    port map (
            O => \N__17571\,
            I => \N__17540\
        );

    \I__3792\ : InMux
    port map (
            O => \N__17570\,
            I => \N__17540\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__17561\,
            I => \N__17533\
        );

    \I__3790\ : Span4Mux_h
    port map (
            O => \N__17558\,
            I => \N__17526\
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__17549\,
            I => \N__17526\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__17540\,
            I => \N__17526\
        );

    \I__3787\ : InMux
    port map (
            O => \N__17539\,
            I => \N__17517\
        );

    \I__3786\ : InMux
    port map (
            O => \N__17538\,
            I => \N__17517\
        );

    \I__3785\ : InMux
    port map (
            O => \N__17537\,
            I => \N__17517\
        );

    \I__3784\ : InMux
    port map (
            O => \N__17536\,
            I => \N__17517\
        );

    \I__3783\ : Span4Mux_v
    port map (
            O => \N__17533\,
            I => \N__17512\
        );

    \I__3782\ : Span4Mux_h
    port map (
            O => \N__17526\,
            I => \N__17512\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__17517\,
            I => \N__17509\
        );

    \I__3780\ : Span4Mux_h
    port map (
            O => \N__17512\,
            I => \N__17506\
        );

    \I__3779\ : Odrv12
    port map (
            O => \N__17509\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__3778\ : Odrv4
    port map (
            O => \N__17506\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__3777\ : CEMux
    port map (
            O => \N__17501\,
            I => \N__17495\
        );

    \I__3776\ : CEMux
    port map (
            O => \N__17500\,
            I => \N__17492\
        );

    \I__3775\ : CEMux
    port map (
            O => \N__17499\,
            I => \N__17489\
        );

    \I__3774\ : CEMux
    port map (
            O => \N__17498\,
            I => \N__17486\
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__17495\,
            I => \N__17481\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__17492\,
            I => \N__17481\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__17489\,
            I => \N__17478\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__17486\,
            I => \N__17475\
        );

    \I__3769\ : Span4Mux_v
    port map (
            O => \N__17481\,
            I => \N__17472\
        );

    \I__3768\ : Span4Mux_h
    port map (
            O => \N__17478\,
            I => \N__17469\
        );

    \I__3767\ : Sp12to4
    port map (
            O => \N__17475\,
            I => \N__17466\
        );

    \I__3766\ : Span4Mux_h
    port map (
            O => \N__17472\,
            I => \N__17463\
        );

    \I__3765\ : Span4Mux_h
    port map (
            O => \N__17469\,
            I => \N__17460\
        );

    \I__3764\ : Odrv12
    port map (
            O => \N__17466\,
            I => \delay_measurement_inst.delay_hc_timer.N_179_i_g\
        );

    \I__3763\ : Odrv4
    port map (
            O => \N__17463\,
            I => \delay_measurement_inst.delay_hc_timer.N_179_i_g\
        );

    \I__3762\ : Odrv4
    port map (
            O => \N__17460\,
            I => \delay_measurement_inst.delay_hc_timer.N_179_i_g\
        );

    \I__3761\ : InMux
    port map (
            O => \N__17453\,
            I => \N__17448\
        );

    \I__3760\ : InMux
    port map (
            O => \N__17452\,
            I => \N__17445\
        );

    \I__3759\ : InMux
    port map (
            O => \N__17451\,
            I => \N__17442\
        );

    \I__3758\ : LocalMux
    port map (
            O => \N__17448\,
            I => \N__17439\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__17445\,
            I => \N__17435\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__17442\,
            I => \N__17432\
        );

    \I__3755\ : Span4Mux_v
    port map (
            O => \N__17439\,
            I => \N__17429\
        );

    \I__3754\ : InMux
    port map (
            O => \N__17438\,
            I => \N__17426\
        );

    \I__3753\ : Span4Mux_h
    port map (
            O => \N__17435\,
            I => \N__17421\
        );

    \I__3752\ : Span4Mux_v
    port map (
            O => \N__17432\,
            I => \N__17421\
        );

    \I__3751\ : Odrv4
    port map (
            O => \N__17429\,
            I => measured_delay_hc_2
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__17426\,
            I => measured_delay_hc_2
        );

    \I__3749\ : Odrv4
    port map (
            O => \N__17421\,
            I => measured_delay_hc_2
        );

    \I__3748\ : InMux
    port map (
            O => \N__17414\,
            I => \N__17411\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__17411\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto6Z0Z_0\
        );

    \I__3746\ : CascadeMux
    port map (
            O => \N__17408\,
            I => \N__17404\
        );

    \I__3745\ : CascadeMux
    port map (
            O => \N__17407\,
            I => \N__17401\
        );

    \I__3744\ : InMux
    port map (
            O => \N__17404\,
            I => \N__17396\
        );

    \I__3743\ : InMux
    port map (
            O => \N__17401\,
            I => \N__17393\
        );

    \I__3742\ : CascadeMux
    port map (
            O => \N__17400\,
            I => \N__17390\
        );

    \I__3741\ : InMux
    port map (
            O => \N__17399\,
            I => \N__17387\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__17396\,
            I => \N__17384\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__17393\,
            I => \N__17381\
        );

    \I__3738\ : InMux
    port map (
            O => \N__17390\,
            I => \N__17378\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__17387\,
            I => \N__17375\
        );

    \I__3736\ : Span4Mux_v
    port map (
            O => \N__17384\,
            I => \N__17370\
        );

    \I__3735\ : Span4Mux_h
    port map (
            O => \N__17381\,
            I => \N__17370\
        );

    \I__3734\ : LocalMux
    port map (
            O => \N__17378\,
            I => measured_delay_hc_3
        );

    \I__3733\ : Odrv4
    port map (
            O => \N__17375\,
            I => measured_delay_hc_3
        );

    \I__3732\ : Odrv4
    port map (
            O => \N__17370\,
            I => measured_delay_hc_3
        );

    \I__3731\ : CascadeMux
    port map (
            O => \N__17363\,
            I => \N__17359\
        );

    \I__3730\ : InMux
    port map (
            O => \N__17362\,
            I => \N__17356\
        );

    \I__3729\ : InMux
    port map (
            O => \N__17359\,
            I => \N__17352\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__17356\,
            I => \N__17349\
        );

    \I__3727\ : InMux
    port map (
            O => \N__17355\,
            I => \N__17346\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__17352\,
            I => \N__17342\
        );

    \I__3725\ : Span4Mux_v
    port map (
            O => \N__17349\,
            I => \N__17337\
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__17346\,
            I => \N__17337\
        );

    \I__3723\ : InMux
    port map (
            O => \N__17345\,
            I => \N__17334\
        );

    \I__3722\ : Odrv4
    port map (
            O => \N__17342\,
            I => measured_delay_hc_4
        );

    \I__3721\ : Odrv4
    port map (
            O => \N__17337\,
            I => measured_delay_hc_4
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__17334\,
            I => measured_delay_hc_4
        );

    \I__3719\ : InMux
    port map (
            O => \N__17327\,
            I => \N__17324\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__17324\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_4\
        );

    \I__3717\ : InMux
    port map (
            O => \N__17321\,
            I => \N__17317\
        );

    \I__3716\ : InMux
    port map (
            O => \N__17320\,
            I => \N__17314\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__17317\,
            I => \N__17310\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__17314\,
            I => \N__17306\
        );

    \I__3713\ : InMux
    port map (
            O => \N__17313\,
            I => \N__17303\
        );

    \I__3712\ : Span12Mux_h
    port map (
            O => \N__17310\,
            I => \N__17300\
        );

    \I__3711\ : InMux
    port map (
            O => \N__17309\,
            I => \N__17297\
        );

    \I__3710\ : Span4Mux_v
    port map (
            O => \N__17306\,
            I => \N__17292\
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__17303\,
            I => \N__17292\
        );

    \I__3708\ : Odrv12
    port map (
            O => \N__17300\,
            I => measured_delay_hc_12
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__17297\,
            I => measured_delay_hc_12
        );

    \I__3706\ : Odrv4
    port map (
            O => \N__17292\,
            I => measured_delay_hc_12
        );

    \I__3705\ : CascadeMux
    port map (
            O => \N__17285\,
            I => \phase_controller_inst1.stoper_hc.un2_startlt19_0_cascade_\
        );

    \I__3704\ : InMux
    port map (
            O => \N__17282\,
            I => \N__17279\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__17279\,
            I => \N__17275\
        );

    \I__3702\ : InMux
    port map (
            O => \N__17278\,
            I => \N__17272\
        );

    \I__3701\ : Span4Mux_h
    port map (
            O => \N__17275\,
            I => \N__17269\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__17272\,
            I => \N__17266\
        );

    \I__3699\ : Span4Mux_v
    port map (
            O => \N__17269\,
            I => \N__17261\
        );

    \I__3698\ : Span4Mux_h
    port map (
            O => \N__17266\,
            I => \N__17258\
        );

    \I__3697\ : InMux
    port map (
            O => \N__17265\,
            I => \N__17255\
        );

    \I__3696\ : InMux
    port map (
            O => \N__17264\,
            I => \N__17252\
        );

    \I__3695\ : Odrv4
    port map (
            O => \N__17261\,
            I => measured_delay_hc_11
        );

    \I__3694\ : Odrv4
    port map (
            O => \N__17258\,
            I => measured_delay_hc_11
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__17255\,
            I => measured_delay_hc_11
        );

    \I__3692\ : LocalMux
    port map (
            O => \N__17252\,
            I => measured_delay_hc_11
        );

    \I__3691\ : CascadeMux
    port map (
            O => \N__17243\,
            I => \N__17239\
        );

    \I__3690\ : CascadeMux
    port map (
            O => \N__17242\,
            I => \N__17235\
        );

    \I__3689\ : InMux
    port map (
            O => \N__17239\,
            I => \N__17229\
        );

    \I__3688\ : InMux
    port map (
            O => \N__17238\,
            I => \N__17229\
        );

    \I__3687\ : InMux
    port map (
            O => \N__17235\,
            I => \N__17224\
        );

    \I__3686\ : InMux
    port map (
            O => \N__17234\,
            I => \N__17224\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__17229\,
            I => \N__17221\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__17224\,
            I => \N__17218\
        );

    \I__3683\ : Span4Mux_h
    port map (
            O => \N__17221\,
            I => \N__17214\
        );

    \I__3682\ : Span4Mux_h
    port map (
            O => \N__17218\,
            I => \N__17211\
        );

    \I__3681\ : InMux
    port map (
            O => \N__17217\,
            I => \N__17208\
        );

    \I__3680\ : Odrv4
    port map (
            O => \N__17214\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_9\
        );

    \I__3679\ : Odrv4
    port map (
            O => \N__17211\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_9\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__17208\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_9\
        );

    \I__3677\ : InMux
    port map (
            O => \N__17201\,
            I => \N__17198\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__17198\,
            I => \N__17195\
        );

    \I__3675\ : Span4Mux_v
    port map (
            O => \N__17195\,
            I => \N__17192\
        );

    \I__3674\ : Span4Mux_h
    port map (
            O => \N__17192\,
            I => \N__17189\
        );

    \I__3673\ : Odrv4
    port map (
            O => \N__17189\,
            I => \il_max_comp1_D1\
        );

    \I__3672\ : SRMux
    port map (
            O => \N__17186\,
            I => \N__17180\
        );

    \I__3671\ : SRMux
    port map (
            O => \N__17185\,
            I => \N__17176\
        );

    \I__3670\ : SRMux
    port map (
            O => \N__17184\,
            I => \N__17173\
        );

    \I__3669\ : SRMux
    port map (
            O => \N__17183\,
            I => \N__17169\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__17180\,
            I => \N__17166\
        );

    \I__3667\ : SRMux
    port map (
            O => \N__17179\,
            I => \N__17163\
        );

    \I__3666\ : LocalMux
    port map (
            O => \N__17176\,
            I => \N__17160\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__17173\,
            I => \N__17157\
        );

    \I__3664\ : SRMux
    port map (
            O => \N__17172\,
            I => \N__17154\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__17169\,
            I => \N__17151\
        );

    \I__3662\ : Span4Mux_v
    port map (
            O => \N__17166\,
            I => \N__17146\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__17163\,
            I => \N__17146\
        );

    \I__3660\ : Span4Mux_v
    port map (
            O => \N__17160\,
            I => \N__17142\
        );

    \I__3659\ : Span4Mux_h
    port map (
            O => \N__17157\,
            I => \N__17137\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__17154\,
            I => \N__17137\
        );

    \I__3657\ : Span4Mux_h
    port map (
            O => \N__17151\,
            I => \N__17132\
        );

    \I__3656\ : Span4Mux_h
    port map (
            O => \N__17146\,
            I => \N__17132\
        );

    \I__3655\ : InMux
    port map (
            O => \N__17145\,
            I => \N__17129\
        );

    \I__3654\ : Odrv4
    port map (
            O => \N__17142\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNI6L42C_31\
        );

    \I__3653\ : Odrv4
    port map (
            O => \N__17137\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNI6L42C_31\
        );

    \I__3652\ : Odrv4
    port map (
            O => \N__17132\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNI6L42C_31\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__17129\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNI6L42C_31\
        );

    \I__3650\ : InMux
    port map (
            O => \N__17120\,
            I => \N__17117\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__17117\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_0_o2_0_7_9\
        );

    \I__3648\ : InMux
    port map (
            O => \N__17114\,
            I => \N__17111\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__17111\,
            I => \delay_measurement_inst.delay_tr_timer.un1_reset_i_a2_4\
        );

    \I__3646\ : InMux
    port map (
            O => \N__17108\,
            I => \N__17105\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__17105\,
            I => \N__17100\
        );

    \I__3644\ : InMux
    port map (
            O => \N__17104\,
            I => \N__17095\
        );

    \I__3643\ : InMux
    port map (
            O => \N__17103\,
            I => \N__17095\
        );

    \I__3642\ : Odrv4
    port map (
            O => \N__17100\,
            I => \delay_measurement_inst.delay_tr_timer.N_127\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__17095\,
            I => \delay_measurement_inst.delay_tr_timer.N_127\
        );

    \I__3640\ : InMux
    port map (
            O => \N__17090\,
            I => \N__17087\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__17087\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_0_o2_0_6_9\
        );

    \I__3638\ : InMux
    port map (
            O => \N__17084\,
            I => \N__17081\
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__17081\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_0_o2_0_0_9\
        );

    \I__3636\ : InMux
    port map (
            O => \N__17078\,
            I => \N__17075\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__17075\,
            I => \N__17072\
        );

    \I__3634\ : Glb2LocalMux
    port map (
            O => \N__17072\,
            I => \N__17069\
        );

    \I__3633\ : GlobalMux
    port map (
            O => \N__17069\,
            I => clk_12mhz
        );

    \I__3632\ : IoInMux
    port map (
            O => \N__17066\,
            I => \N__17063\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__17063\,
            I => \GB_BUFFER_clk_12mhz_THRU_CO\
        );

    \I__3630\ : InMux
    port map (
            O => \N__17060\,
            I => \N__17057\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__17057\,
            I => delay_hc_d2
        );

    \I__3628\ : InMux
    port map (
            O => \N__17054\,
            I => \N__17051\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__17051\,
            I => \delay_measurement_inst.hc_syncZ0Z_0\
        );

    \I__3626\ : InMux
    port map (
            O => \N__17048\,
            I => \N__17045\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__17045\,
            I => \N__17041\
        );

    \I__3624\ : InMux
    port map (
            O => \N__17044\,
            I => \N__17036\
        );

    \I__3623\ : Span4Mux_h
    port map (
            O => \N__17041\,
            I => \N__17033\
        );

    \I__3622\ : InMux
    port map (
            O => \N__17040\,
            I => \N__17030\
        );

    \I__3621\ : InMux
    port map (
            O => \N__17039\,
            I => \N__17027\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__17036\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__3619\ : Odrv4
    port map (
            O => \N__17033\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__17030\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__17027\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__3616\ : CascadeMux
    port map (
            O => \N__17018\,
            I => \N__17015\
        );

    \I__3615\ : InMux
    port map (
            O => \N__17015\,
            I => \N__17012\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__17012\,
            I => \N__17009\
        );

    \I__3613\ : Span4Mux_h
    port map (
            O => \N__17009\,
            I => \N__17006\
        );

    \I__3612\ : Span4Mux_h
    port map (
            O => \N__17006\,
            I => \N__17003\
        );

    \I__3611\ : Odrv4
    port map (
            O => \N__17003\,
            I => \delay_measurement_inst.elapsed_time_tr_1\
        );

    \I__3610\ : InMux
    port map (
            O => \N__17000\,
            I => \N__16996\
        );

    \I__3609\ : InMux
    port map (
            O => \N__16999\,
            I => \N__16993\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__16996\,
            I => \N__16990\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__16993\,
            I => \delay_measurement_inst.elapsed_time_tr_2\
        );

    \I__3606\ : Odrv4
    port map (
            O => \N__16990\,
            I => \delay_measurement_inst.elapsed_time_tr_2\
        );

    \I__3605\ : InMux
    port map (
            O => \N__16985\,
            I => \N__16977\
        );

    \I__3604\ : InMux
    port map (
            O => \N__16984\,
            I => \N__16971\
        );

    \I__3603\ : InMux
    port map (
            O => \N__16983\,
            I => \N__16968\
        );

    \I__3602\ : InMux
    port map (
            O => \N__16982\,
            I => \N__16961\
        );

    \I__3601\ : InMux
    port map (
            O => \N__16981\,
            I => \N__16961\
        );

    \I__3600\ : InMux
    port map (
            O => \N__16980\,
            I => \N__16961\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__16977\,
            I => \N__16958\
        );

    \I__3598\ : InMux
    port map (
            O => \N__16976\,
            I => \N__16955\
        );

    \I__3597\ : InMux
    port map (
            O => \N__16975\,
            I => \N__16952\
        );

    \I__3596\ : InMux
    port map (
            O => \N__16974\,
            I => \N__16949\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__16971\,
            I => \delay_measurement_inst.N_201\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__16968\,
            I => \delay_measurement_inst.N_201\
        );

    \I__3593\ : LocalMux
    port map (
            O => \N__16961\,
            I => \delay_measurement_inst.N_201\
        );

    \I__3592\ : Odrv4
    port map (
            O => \N__16958\,
            I => \delay_measurement_inst.N_201\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__16955\,
            I => \delay_measurement_inst.N_201\
        );

    \I__3590\ : LocalMux
    port map (
            O => \N__16952\,
            I => \delay_measurement_inst.N_201\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__16949\,
            I => \delay_measurement_inst.N_201\
        );

    \I__3588\ : InMux
    port map (
            O => \N__16934\,
            I => \N__16930\
        );

    \I__3587\ : InMux
    port map (
            O => \N__16933\,
            I => \N__16927\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__16930\,
            I => \N__16920\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__16927\,
            I => \N__16920\
        );

    \I__3584\ : InMux
    port map (
            O => \N__16926\,
            I => \N__16917\
        );

    \I__3583\ : InMux
    port map (
            O => \N__16925\,
            I => \N__16914\
        );

    \I__3582\ : Span4Mux_v
    port map (
            O => \N__16920\,
            I => \N__16911\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__16917\,
            I => \N__16908\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__16914\,
            I => \N__16905\
        );

    \I__3579\ : Span4Mux_h
    port map (
            O => \N__16911\,
            I => \N__16900\
        );

    \I__3578\ : Span4Mux_v
    port map (
            O => \N__16908\,
            I => \N__16900\
        );

    \I__3577\ : Span4Mux_h
    port map (
            O => \N__16905\,
            I => \N__16897\
        );

    \I__3576\ : Odrv4
    port map (
            O => \N__16900\,
            I => measured_delay_tr_19
        );

    \I__3575\ : Odrv4
    port map (
            O => \N__16897\,
            I => measured_delay_tr_19
        );

    \I__3574\ : CEMux
    port map (
            O => \N__16892\,
            I => \N__16888\
        );

    \I__3573\ : CEMux
    port map (
            O => \N__16891\,
            I => \N__16883\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__16888\,
            I => \N__16880\
        );

    \I__3571\ : CEMux
    port map (
            O => \N__16887\,
            I => \N__16877\
        );

    \I__3570\ : CEMux
    port map (
            O => \N__16886\,
            I => \N__16874\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__16883\,
            I => \N__16871\
        );

    \I__3568\ : Span4Mux_h
    port map (
            O => \N__16880\,
            I => \N__16866\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__16877\,
            I => \N__16866\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__16874\,
            I => \N__16863\
        );

    \I__3565\ : Span4Mux_h
    port map (
            O => \N__16871\,
            I => \N__16860\
        );

    \I__3564\ : Span4Mux_h
    port map (
            O => \N__16866\,
            I => \N__16855\
        );

    \I__3563\ : Span4Mux_h
    port map (
            O => \N__16863\,
            I => \N__16855\
        );

    \I__3562\ : Odrv4
    port map (
            O => \N__16860\,
            I => \delay_measurement_inst.N_134_i_0\
        );

    \I__3561\ : Odrv4
    port map (
            O => \N__16855\,
            I => \delay_measurement_inst.N_134_i_0\
        );

    \I__3560\ : CascadeMux
    port map (
            O => \N__16850\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0_cascade_\
        );

    \I__3559\ : InMux
    port map (
            O => \N__16847\,
            I => \N__16843\
        );

    \I__3558\ : InMux
    port map (
            O => \N__16846\,
            I => \N__16840\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__16843\,
            I => \N__16837\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__16840\,
            I => \N__16832\
        );

    \I__3555\ : Span4Mux_h
    port map (
            O => \N__16837\,
            I => \N__16829\
        );

    \I__3554\ : InMux
    port map (
            O => \N__16836\,
            I => \N__16826\
        );

    \I__3553\ : InMux
    port map (
            O => \N__16835\,
            I => \N__16823\
        );

    \I__3552\ : Odrv4
    port map (
            O => \N__16832\,
            I => measured_delay_hc_6
        );

    \I__3551\ : Odrv4
    port map (
            O => \N__16829\,
            I => measured_delay_hc_6
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__16826\,
            I => measured_delay_hc_6
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__16823\,
            I => measured_delay_hc_6
        );

    \I__3548\ : InMux
    port map (
            O => \N__16814\,
            I => \N__16811\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__16811\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ1Z_6\
        );

    \I__3546\ : InMux
    port map (
            O => \N__16808\,
            I => \N__16805\
        );

    \I__3545\ : LocalMux
    port map (
            O => \N__16805\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\
        );

    \I__3544\ : InMux
    port map (
            O => \N__16802\,
            I => \N__16798\
        );

    \I__3543\ : InMux
    port map (
            O => \N__16801\,
            I => \N__16795\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__16798\,
            I => \N__16792\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__16795\,
            I => \N__16786\
        );

    \I__3540\ : Span4Mux_v
    port map (
            O => \N__16792\,
            I => \N__16783\
        );

    \I__3539\ : InMux
    port map (
            O => \N__16791\,
            I => \N__16776\
        );

    \I__3538\ : InMux
    port map (
            O => \N__16790\,
            I => \N__16776\
        );

    \I__3537\ : InMux
    port map (
            O => \N__16789\,
            I => \N__16776\
        );

    \I__3536\ : Odrv12
    port map (
            O => \N__16786\,
            I => measured_delay_hc_9
        );

    \I__3535\ : Odrv4
    port map (
            O => \N__16783\,
            I => measured_delay_hc_9
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__16776\,
            I => measured_delay_hc_9
        );

    \I__3533\ : InMux
    port map (
            O => \N__16769\,
            I => \N__16766\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__16766\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\
        );

    \I__3531\ : InMux
    port map (
            O => \N__16763\,
            I => \N__16760\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__16760\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\
        );

    \I__3529\ : CascadeMux
    port map (
            O => \N__16757\,
            I => \N__16753\
        );

    \I__3528\ : CascadeMux
    port map (
            O => \N__16756\,
            I => \N__16750\
        );

    \I__3527\ : InMux
    port map (
            O => \N__16753\,
            I => \N__16747\
        );

    \I__3526\ : InMux
    port map (
            O => \N__16750\,
            I => \N__16744\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__16747\,
            I => \N__16740\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__16744\,
            I => \N__16737\
        );

    \I__3523\ : InMux
    port map (
            O => \N__16743\,
            I => \N__16734\
        );

    \I__3522\ : Odrv4
    port map (
            O => \N__16740\,
            I => measured_delay_hc_13
        );

    \I__3521\ : Odrv12
    port map (
            O => \N__16737\,
            I => measured_delay_hc_13
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__16734\,
            I => measured_delay_hc_13
        );

    \I__3519\ : InMux
    port map (
            O => \N__16727\,
            I => \N__16724\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__16724\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\
        );

    \I__3517\ : InMux
    port map (
            O => \N__16721\,
            I => \N__16700\
        );

    \I__3516\ : InMux
    port map (
            O => \N__16720\,
            I => \N__16700\
        );

    \I__3515\ : InMux
    port map (
            O => \N__16719\,
            I => \N__16700\
        );

    \I__3514\ : InMux
    port map (
            O => \N__16718\,
            I => \N__16700\
        );

    \I__3513\ : InMux
    port map (
            O => \N__16717\,
            I => \N__16700\
        );

    \I__3512\ : InMux
    port map (
            O => \N__16716\,
            I => \N__16697\
        );

    \I__3511\ : InMux
    port map (
            O => \N__16715\,
            I => \N__16686\
        );

    \I__3510\ : InMux
    port map (
            O => \N__16714\,
            I => \N__16686\
        );

    \I__3509\ : InMux
    port map (
            O => \N__16713\,
            I => \N__16686\
        );

    \I__3508\ : InMux
    port map (
            O => \N__16712\,
            I => \N__16686\
        );

    \I__3507\ : InMux
    port map (
            O => \N__16711\,
            I => \N__16686\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__16700\,
            I => \N__16672\
        );

    \I__3505\ : LocalMux
    port map (
            O => \N__16697\,
            I => \N__16667\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__16686\,
            I => \N__16667\
        );

    \I__3503\ : InMux
    port map (
            O => \N__16685\,
            I => \N__16656\
        );

    \I__3502\ : InMux
    port map (
            O => \N__16684\,
            I => \N__16656\
        );

    \I__3501\ : InMux
    port map (
            O => \N__16683\,
            I => \N__16656\
        );

    \I__3500\ : InMux
    port map (
            O => \N__16682\,
            I => \N__16656\
        );

    \I__3499\ : InMux
    port map (
            O => \N__16681\,
            I => \N__16656\
        );

    \I__3498\ : InMux
    port map (
            O => \N__16680\,
            I => \N__16643\
        );

    \I__3497\ : InMux
    port map (
            O => \N__16679\,
            I => \N__16643\
        );

    \I__3496\ : InMux
    port map (
            O => \N__16678\,
            I => \N__16643\
        );

    \I__3495\ : InMux
    port map (
            O => \N__16677\,
            I => \N__16643\
        );

    \I__3494\ : InMux
    port map (
            O => \N__16676\,
            I => \N__16643\
        );

    \I__3493\ : InMux
    port map (
            O => \N__16675\,
            I => \N__16643\
        );

    \I__3492\ : Span4Mux_v
    port map (
            O => \N__16672\,
            I => \N__16639\
        );

    \I__3491\ : Span4Mux_v
    port map (
            O => \N__16667\,
            I => \N__16632\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__16656\,
            I => \N__16632\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__16643\,
            I => \N__16632\
        );

    \I__3488\ : InMux
    port map (
            O => \N__16642\,
            I => \N__16629\
        );

    \I__3487\ : Odrv4
    port map (
            O => \N__16639\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt15\
        );

    \I__3486\ : Odrv4
    port map (
            O => \N__16632\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt15\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__16629\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt15\
        );

    \I__3484\ : CascadeMux
    port map (
            O => \N__16622\,
            I => \N__16617\
        );

    \I__3483\ : CascadeMux
    port map (
            O => \N__16621\,
            I => \N__16614\
        );

    \I__3482\ : CascadeMux
    port map (
            O => \N__16620\,
            I => \N__16611\
        );

    \I__3481\ : InMux
    port map (
            O => \N__16617\,
            I => \N__16590\
        );

    \I__3480\ : InMux
    port map (
            O => \N__16614\,
            I => \N__16590\
        );

    \I__3479\ : InMux
    port map (
            O => \N__16611\,
            I => \N__16590\
        );

    \I__3478\ : InMux
    port map (
            O => \N__16610\,
            I => \N__16590\
        );

    \I__3477\ : InMux
    port map (
            O => \N__16609\,
            I => \N__16590\
        );

    \I__3476\ : CascadeMux
    port map (
            O => \N__16608\,
            I => \N__16587\
        );

    \I__3475\ : CascadeMux
    port map (
            O => \N__16607\,
            I => \N__16584\
        );

    \I__3474\ : CascadeMux
    port map (
            O => \N__16606\,
            I => \N__16581\
        );

    \I__3473\ : InMux
    port map (
            O => \N__16605\,
            I => \N__16576\
        );

    \I__3472\ : InMux
    port map (
            O => \N__16604\,
            I => \N__16567\
        );

    \I__3471\ : InMux
    port map (
            O => \N__16603\,
            I => \N__16567\
        );

    \I__3470\ : InMux
    port map (
            O => \N__16602\,
            I => \N__16567\
        );

    \I__3469\ : InMux
    port map (
            O => \N__16601\,
            I => \N__16567\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__16590\,
            I => \N__16559\
        );

    \I__3467\ : InMux
    port map (
            O => \N__16587\,
            I => \N__16548\
        );

    \I__3466\ : InMux
    port map (
            O => \N__16584\,
            I => \N__16548\
        );

    \I__3465\ : InMux
    port map (
            O => \N__16581\,
            I => \N__16548\
        );

    \I__3464\ : InMux
    port map (
            O => \N__16580\,
            I => \N__16548\
        );

    \I__3463\ : InMux
    port map (
            O => \N__16579\,
            I => \N__16548\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__16576\,
            I => \N__16545\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__16567\,
            I => \N__16542\
        );

    \I__3460\ : InMux
    port map (
            O => \N__16566\,
            I => \N__16531\
        );

    \I__3459\ : InMux
    port map (
            O => \N__16565\,
            I => \N__16531\
        );

    \I__3458\ : InMux
    port map (
            O => \N__16564\,
            I => \N__16531\
        );

    \I__3457\ : InMux
    port map (
            O => \N__16563\,
            I => \N__16531\
        );

    \I__3456\ : InMux
    port map (
            O => \N__16562\,
            I => \N__16531\
        );

    \I__3455\ : Span4Mux_v
    port map (
            O => \N__16559\,
            I => \N__16528\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__16548\,
            I => \N__16521\
        );

    \I__3453\ : Span4Mux_v
    port map (
            O => \N__16545\,
            I => \N__16521\
        );

    \I__3452\ : Span4Mux_v
    port map (
            O => \N__16542\,
            I => \N__16521\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__16531\,
            I => \phase_controller_inst1.stoper_hc.un3_start\
        );

    \I__3450\ : Odrv4
    port map (
            O => \N__16528\,
            I => \phase_controller_inst1.stoper_hc.un3_start\
        );

    \I__3449\ : Odrv4
    port map (
            O => \N__16521\,
            I => \phase_controller_inst1.stoper_hc.un3_start\
        );

    \I__3448\ : InMux
    port map (
            O => \N__16514\,
            I => \N__16510\
        );

    \I__3447\ : InMux
    port map (
            O => \N__16513\,
            I => \N__16507\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__16510\,
            I => \N__16503\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__16507\,
            I => \N__16500\
        );

    \I__3444\ : InMux
    port map (
            O => \N__16506\,
            I => \N__16497\
        );

    \I__3443\ : Odrv12
    port map (
            O => \N__16503\,
            I => measured_delay_hc_10
        );

    \I__3442\ : Odrv4
    port map (
            O => \N__16500\,
            I => measured_delay_hc_10
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__16497\,
            I => measured_delay_hc_10
        );

    \I__3440\ : InMux
    port map (
            O => \N__16490\,
            I => \N__16487\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__16487\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\
        );

    \I__3438\ : InMux
    port map (
            O => \N__16484\,
            I => \N__16481\
        );

    \I__3437\ : LocalMux
    port map (
            O => \N__16481\,
            I => \N__16477\
        );

    \I__3436\ : InMux
    port map (
            O => \N__16480\,
            I => \N__16474\
        );

    \I__3435\ : Span4Mux_v
    port map (
            O => \N__16477\,
            I => \N__16469\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__16474\,
            I => \N__16469\
        );

    \I__3433\ : Span4Mux_v
    port map (
            O => \N__16469\,
            I => \N__16464\
        );

    \I__3432\ : InMux
    port map (
            O => \N__16468\,
            I => \N__16461\
        );

    \I__3431\ : InMux
    port map (
            O => \N__16467\,
            I => \N__16458\
        );

    \I__3430\ : Odrv4
    port map (
            O => \N__16464\,
            I => measured_delay_hc_14
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__16461\,
            I => measured_delay_hc_14
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__16458\,
            I => measured_delay_hc_14
        );

    \I__3427\ : InMux
    port map (
            O => \N__16451\,
            I => \N__16448\
        );

    \I__3426\ : LocalMux
    port map (
            O => \N__16448\,
            I => \N__16445\
        );

    \I__3425\ : Odrv4
    port map (
            O => \N__16445\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\
        );

    \I__3424\ : CascadeMux
    port map (
            O => \N__16442\,
            I => \N__16431\
        );

    \I__3423\ : CascadeMux
    port map (
            O => \N__16441\,
            I => \N__16425\
        );

    \I__3422\ : CascadeMux
    port map (
            O => \N__16440\,
            I => \N__16422\
        );

    \I__3421\ : CascadeMux
    port map (
            O => \N__16439\,
            I => \N__16419\
        );

    \I__3420\ : CascadeMux
    port map (
            O => \N__16438\,
            I => \N__16416\
        );

    \I__3419\ : InMux
    port map (
            O => \N__16437\,
            I => \N__16401\
        );

    \I__3418\ : InMux
    port map (
            O => \N__16436\,
            I => \N__16401\
        );

    \I__3417\ : InMux
    port map (
            O => \N__16435\,
            I => \N__16401\
        );

    \I__3416\ : InMux
    port map (
            O => \N__16434\,
            I => \N__16401\
        );

    \I__3415\ : InMux
    port map (
            O => \N__16431\,
            I => \N__16401\
        );

    \I__3414\ : InMux
    port map (
            O => \N__16430\,
            I => \N__16393\
        );

    \I__3413\ : InMux
    port map (
            O => \N__16429\,
            I => \N__16393\
        );

    \I__3412\ : InMux
    port map (
            O => \N__16428\,
            I => \N__16380\
        );

    \I__3411\ : InMux
    port map (
            O => \N__16425\,
            I => \N__16380\
        );

    \I__3410\ : InMux
    port map (
            O => \N__16422\,
            I => \N__16380\
        );

    \I__3409\ : InMux
    port map (
            O => \N__16419\,
            I => \N__16380\
        );

    \I__3408\ : InMux
    port map (
            O => \N__16416\,
            I => \N__16380\
        );

    \I__3407\ : InMux
    port map (
            O => \N__16415\,
            I => \N__16380\
        );

    \I__3406\ : CascadeMux
    port map (
            O => \N__16414\,
            I => \N__16377\
        );

    \I__3405\ : CascadeMux
    port map (
            O => \N__16413\,
            I => \N__16374\
        );

    \I__3404\ : CascadeMux
    port map (
            O => \N__16412\,
            I => \N__16367\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__16401\,
            I => \N__16363\
        );

    \I__3402\ : CascadeMux
    port map (
            O => \N__16400\,
            I => \N__16360\
        );

    \I__3401\ : CascadeMux
    port map (
            O => \N__16399\,
            I => \N__16357\
        );

    \I__3400\ : CascadeMux
    port map (
            O => \N__16398\,
            I => \N__16352\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__16393\,
            I => \N__16347\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__16380\,
            I => \N__16347\
        );

    \I__3397\ : InMux
    port map (
            O => \N__16377\,
            I => \N__16330\
        );

    \I__3396\ : InMux
    port map (
            O => \N__16374\,
            I => \N__16330\
        );

    \I__3395\ : InMux
    port map (
            O => \N__16373\,
            I => \N__16330\
        );

    \I__3394\ : InMux
    port map (
            O => \N__16372\,
            I => \N__16330\
        );

    \I__3393\ : InMux
    port map (
            O => \N__16371\,
            I => \N__16330\
        );

    \I__3392\ : InMux
    port map (
            O => \N__16370\,
            I => \N__16330\
        );

    \I__3391\ : InMux
    port map (
            O => \N__16367\,
            I => \N__16330\
        );

    \I__3390\ : InMux
    port map (
            O => \N__16366\,
            I => \N__16330\
        );

    \I__3389\ : Span4Mux_h
    port map (
            O => \N__16363\,
            I => \N__16326\
        );

    \I__3388\ : InMux
    port map (
            O => \N__16360\,
            I => \N__16315\
        );

    \I__3387\ : InMux
    port map (
            O => \N__16357\,
            I => \N__16315\
        );

    \I__3386\ : InMux
    port map (
            O => \N__16356\,
            I => \N__16315\
        );

    \I__3385\ : InMux
    port map (
            O => \N__16355\,
            I => \N__16315\
        );

    \I__3384\ : InMux
    port map (
            O => \N__16352\,
            I => \N__16315\
        );

    \I__3383\ : Span4Mux_v
    port map (
            O => \N__16347\,
            I => \N__16310\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__16330\,
            I => \N__16310\
        );

    \I__3381\ : InMux
    port map (
            O => \N__16329\,
            I => \N__16307\
        );

    \I__3380\ : Odrv4
    port map (
            O => \N__16326\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__16315\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2\
        );

    \I__3378\ : Odrv4
    port map (
            O => \N__16310\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__16307\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2\
        );

    \I__3376\ : InMux
    port map (
            O => \N__16298\,
            I => \N__16295\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__16295\,
            I => \N__16292\
        );

    \I__3374\ : Odrv4
    port map (
            O => \N__16292\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\
        );

    \I__3373\ : InMux
    port map (
            O => \N__16289\,
            I => \N__16286\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__16286\,
            I => \N__16280\
        );

    \I__3371\ : InMux
    port map (
            O => \N__16285\,
            I => \N__16277\
        );

    \I__3370\ : InMux
    port map (
            O => \N__16284\,
            I => \N__16272\
        );

    \I__3369\ : InMux
    port map (
            O => \N__16283\,
            I => \N__16272\
        );

    \I__3368\ : Odrv4
    port map (
            O => \N__16280\,
            I => measured_delay_hc_5
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__16277\,
            I => measured_delay_hc_5
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__16272\,
            I => measured_delay_hc_5
        );

    \I__3365\ : InMux
    port map (
            O => \N__16265\,
            I => \N__16262\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__16262\,
            I => \N__16256\
        );

    \I__3363\ : InMux
    port map (
            O => \N__16261\,
            I => \N__16253\
        );

    \I__3362\ : InMux
    port map (
            O => \N__16260\,
            I => \N__16248\
        );

    \I__3361\ : InMux
    port map (
            O => \N__16259\,
            I => \N__16248\
        );

    \I__3360\ : Span4Mux_v
    port map (
            O => \N__16256\,
            I => \N__16245\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__16253\,
            I => \N__16242\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__16248\,
            I => \N__16239\
        );

    \I__3357\ : Odrv4
    port map (
            O => \N__16245\,
            I => measured_delay_hc_16
        );

    \I__3356\ : Odrv4
    port map (
            O => \N__16242\,
            I => measured_delay_hc_16
        );

    \I__3355\ : Odrv4
    port map (
            O => \N__16239\,
            I => measured_delay_hc_16
        );

    \I__3354\ : InMux
    port map (
            O => \N__16232\,
            I => \N__16229\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__16229\,
            I => \N__16223\
        );

    \I__3352\ : InMux
    port map (
            O => \N__16228\,
            I => \N__16220\
        );

    \I__3351\ : InMux
    port map (
            O => \N__16227\,
            I => \N__16215\
        );

    \I__3350\ : InMux
    port map (
            O => \N__16226\,
            I => \N__16215\
        );

    \I__3349\ : Span4Mux_v
    port map (
            O => \N__16223\,
            I => \N__16212\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__16220\,
            I => \N__16209\
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__16215\,
            I => \N__16206\
        );

    \I__3346\ : Odrv4
    port map (
            O => \N__16212\,
            I => measured_delay_hc_19
        );

    \I__3345\ : Odrv4
    port map (
            O => \N__16209\,
            I => measured_delay_hc_19
        );

    \I__3344\ : Odrv4
    port map (
            O => \N__16206\,
            I => measured_delay_hc_19
        );

    \I__3343\ : InMux
    port map (
            O => \N__16199\,
            I => \N__16196\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__16196\,
            I => \N__16190\
        );

    \I__3341\ : InMux
    port map (
            O => \N__16195\,
            I => \N__16187\
        );

    \I__3340\ : CascadeMux
    port map (
            O => \N__16194\,
            I => \N__16184\
        );

    \I__3339\ : CascadeMux
    port map (
            O => \N__16193\,
            I => \N__16181\
        );

    \I__3338\ : Span4Mux_v
    port map (
            O => \N__16190\,
            I => \N__16176\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__16187\,
            I => \N__16176\
        );

    \I__3336\ : InMux
    port map (
            O => \N__16184\,
            I => \N__16171\
        );

    \I__3335\ : InMux
    port map (
            O => \N__16181\,
            I => \N__16171\
        );

    \I__3334\ : Odrv4
    port map (
            O => \N__16176\,
            I => measured_delay_hc_17
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__16171\,
            I => measured_delay_hc_17
        );

    \I__3332\ : InMux
    port map (
            O => \N__16166\,
            I => \N__16162\
        );

    \I__3331\ : InMux
    port map (
            O => \N__16165\,
            I => \N__16157\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__16162\,
            I => \N__16154\
        );

    \I__3329\ : InMux
    port map (
            O => \N__16161\,
            I => \N__16149\
        );

    \I__3328\ : InMux
    port map (
            O => \N__16160\,
            I => \N__16149\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__16157\,
            I => \N__16146\
        );

    \I__3326\ : Span4Mux_v
    port map (
            O => \N__16154\,
            I => \N__16141\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__16149\,
            I => \N__16141\
        );

    \I__3324\ : Odrv12
    port map (
            O => \N__16146\,
            I => measured_delay_hc_18
        );

    \I__3323\ : Odrv4
    port map (
            O => \N__16141\,
            I => measured_delay_hc_18
        );

    \I__3322\ : CascadeMux
    port map (
            O => \N__16136\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2_cascade_\
        );

    \I__3321\ : InMux
    port map (
            O => \N__16133\,
            I => \N__16127\
        );

    \I__3320\ : InMux
    port map (
            O => \N__16132\,
            I => \N__16127\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__16127\,
            I => \N__16124\
        );

    \I__3318\ : Span4Mux_h
    port map (
            O => \N__16124\,
            I => \N__16119\
        );

    \I__3317\ : InMux
    port map (
            O => \N__16123\,
            I => \N__16114\
        );

    \I__3316\ : InMux
    port map (
            O => \N__16122\,
            I => \N__16114\
        );

    \I__3315\ : Odrv4
    port map (
            O => \N__16119\,
            I => \phase_controller_inst1.stoper_hc.un1_start\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__16114\,
            I => \phase_controller_inst1.stoper_hc.un1_start\
        );

    \I__3313\ : CascadeMux
    port map (
            O => \N__16109\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt8_cascade_\
        );

    \I__3312\ : CascadeMux
    port map (
            O => \N__16106\,
            I => \N__16103\
        );

    \I__3311\ : InMux
    port map (
            O => \N__16103\,
            I => \N__16098\
        );

    \I__3310\ : CascadeMux
    port map (
            O => \N__16102\,
            I => \N__16094\
        );

    \I__3309\ : InMux
    port map (
            O => \N__16101\,
            I => \N__16091\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__16098\,
            I => \N__16088\
        );

    \I__3307\ : CascadeMux
    port map (
            O => \N__16097\,
            I => \N__16085\
        );

    \I__3306\ : InMux
    port map (
            O => \N__16094\,
            I => \N__16081\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__16091\,
            I => \N__16076\
        );

    \I__3304\ : Span4Mux_v
    port map (
            O => \N__16088\,
            I => \N__16076\
        );

    \I__3303\ : InMux
    port map (
            O => \N__16085\,
            I => \N__16071\
        );

    \I__3302\ : InMux
    port map (
            O => \N__16084\,
            I => \N__16071\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__16081\,
            I => measured_delay_hc_8
        );

    \I__3300\ : Odrv4
    port map (
            O => \N__16076\,
            I => measured_delay_hc_8
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__16071\,
            I => measured_delay_hc_8
        );

    \I__3298\ : CascadeMux
    port map (
            O => \N__16064\,
            I => \N__16059\
        );

    \I__3297\ : InMux
    port map (
            O => \N__16063\,
            I => \N__16056\
        );

    \I__3296\ : InMux
    port map (
            O => \N__16062\,
            I => \N__16053\
        );

    \I__3295\ : InMux
    port map (
            O => \N__16059\,
            I => \N__16048\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__16056\,
            I => \N__16043\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__16053\,
            I => \N__16043\
        );

    \I__3292\ : InMux
    port map (
            O => \N__16052\,
            I => \N__16038\
        );

    \I__3291\ : InMux
    port map (
            O => \N__16051\,
            I => \N__16038\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__16048\,
            I => measured_delay_hc_7
        );

    \I__3289\ : Odrv12
    port map (
            O => \N__16043\,
            I => measured_delay_hc_7
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__16038\,
            I => measured_delay_hc_7
        );

    \I__3287\ : CascadeMux
    port map (
            O => \N__16031\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto9_cZ0_cascade_\
        );

    \I__3286\ : InMux
    port map (
            O => \N__16028\,
            I => \N__16025\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__16025\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto13\
        );

    \I__3284\ : InMux
    port map (
            O => \N__16022\,
            I => \N__16019\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__16019\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_6\
        );

    \I__3282\ : CascadeMux
    port map (
            O => \N__16016\,
            I => \N__16012\
        );

    \I__3281\ : InMux
    port map (
            O => \N__16015\,
            I => \N__16006\
        );

    \I__3280\ : InMux
    port map (
            O => \N__16012\,
            I => \N__16006\
        );

    \I__3279\ : CascadeMux
    port map (
            O => \N__16011\,
            I => \N__16002\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__16006\,
            I => \N__15999\
        );

    \I__3277\ : InMux
    port map (
            O => \N__16005\,
            I => \N__15994\
        );

    \I__3276\ : InMux
    port map (
            O => \N__16002\,
            I => \N__15994\
        );

    \I__3275\ : Span4Mux_v
    port map (
            O => \N__15999\,
            I => \N__15991\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__15994\,
            I => \N__15988\
        );

    \I__3273\ : Odrv4
    port map (
            O => \N__15991\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_8\
        );

    \I__3272\ : Odrv4
    port map (
            O => \N__15988\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_8\
        );

    \I__3271\ : CascadeMux
    port map (
            O => \N__15983\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_8_cascade_\
        );

    \I__3270\ : InMux
    port map (
            O => \N__15980\,
            I => \N__15977\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__15977\,
            I => \N__15974\
        );

    \I__3268\ : Span4Mux_v
    port map (
            O => \N__15974\,
            I => \N__15969\
        );

    \I__3267\ : InMux
    port map (
            O => \N__15973\,
            I => \N__15966\
        );

    \I__3266\ : InMux
    port map (
            O => \N__15972\,
            I => \N__15963\
        );

    \I__3265\ : Odrv4
    port map (
            O => \N__15969\,
            I => measured_delay_hc_1
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__15966\,
            I => measured_delay_hc_1
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__15963\,
            I => measured_delay_hc_1
        );

    \I__3262\ : InMux
    port map (
            O => \N__15956\,
            I => \N__15953\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__15953\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_1\
        );

    \I__3260\ : InMux
    port map (
            O => \N__15950\,
            I => \N__15946\
        );

    \I__3259\ : InMux
    port map (
            O => \N__15949\,
            I => \N__15943\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__15946\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_2\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__15943\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_2\
        );

    \I__3256\ : InMux
    port map (
            O => \N__15938\,
            I => \N__15930\
        );

    \I__3255\ : InMux
    port map (
            O => \N__15937\,
            I => \N__15930\
        );

    \I__3254\ : InMux
    port map (
            O => \N__15936\,
            I => \N__15927\
        );

    \I__3253\ : CascadeMux
    port map (
            O => \N__15935\,
            I => \N__15923\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__15930\,
            I => \N__15919\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__15927\,
            I => \N__15916\
        );

    \I__3250\ : InMux
    port map (
            O => \N__15926\,
            I => \N__15913\
        );

    \I__3249\ : InMux
    port map (
            O => \N__15923\,
            I => \N__15908\
        );

    \I__3248\ : InMux
    port map (
            O => \N__15922\,
            I => \N__15908\
        );

    \I__3247\ : Odrv4
    port map (
            O => \N__15919\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__3246\ : Odrv4
    port map (
            O => \N__15916\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__15913\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__15908\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__3243\ : CascadeMux
    port map (
            O => \N__15899\,
            I => \N__15894\
        );

    \I__3242\ : CascadeMux
    port map (
            O => \N__15898\,
            I => \N__15891\
        );

    \I__3241\ : CascadeMux
    port map (
            O => \N__15897\,
            I => \N__15879\
        );

    \I__3240\ : InMux
    port map (
            O => \N__15894\,
            I => \N__15874\
        );

    \I__3239\ : InMux
    port map (
            O => \N__15891\,
            I => \N__15874\
        );

    \I__3238\ : InMux
    port map (
            O => \N__15890\,
            I => \N__15871\
        );

    \I__3237\ : InMux
    port map (
            O => \N__15889\,
            I => \N__15868\
        );

    \I__3236\ : InMux
    port map (
            O => \N__15888\,
            I => \N__15855\
        );

    \I__3235\ : InMux
    port map (
            O => \N__15887\,
            I => \N__15855\
        );

    \I__3234\ : InMux
    port map (
            O => \N__15886\,
            I => \N__15855\
        );

    \I__3233\ : InMux
    port map (
            O => \N__15885\,
            I => \N__15855\
        );

    \I__3232\ : InMux
    port map (
            O => \N__15884\,
            I => \N__15855\
        );

    \I__3231\ : InMux
    port map (
            O => \N__15883\,
            I => \N__15855\
        );

    \I__3230\ : InMux
    port map (
            O => \N__15882\,
            I => \N__15846\
        );

    \I__3229\ : InMux
    port map (
            O => \N__15879\,
            I => \N__15843\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__15874\,
            I => \N__15840\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__15871\,
            I => \N__15835\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__15868\,
            I => \N__15835\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__15855\,
            I => \N__15824\
        );

    \I__3224\ : InMux
    port map (
            O => \N__15854\,
            I => \N__15817\
        );

    \I__3223\ : InMux
    port map (
            O => \N__15853\,
            I => \N__15817\
        );

    \I__3222\ : InMux
    port map (
            O => \N__15852\,
            I => \N__15817\
        );

    \I__3221\ : InMux
    port map (
            O => \N__15851\,
            I => \N__15810\
        );

    \I__3220\ : InMux
    port map (
            O => \N__15850\,
            I => \N__15810\
        );

    \I__3219\ : InMux
    port map (
            O => \N__15849\,
            I => \N__15810\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__15846\,
            I => \N__15807\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__15843\,
            I => \N__15800\
        );

    \I__3216\ : Span4Mux_v
    port map (
            O => \N__15840\,
            I => \N__15800\
        );

    \I__3215\ : Span4Mux_v
    port map (
            O => \N__15835\,
            I => \N__15800\
        );

    \I__3214\ : InMux
    port map (
            O => \N__15834\,
            I => \N__15783\
        );

    \I__3213\ : InMux
    port map (
            O => \N__15833\,
            I => \N__15783\
        );

    \I__3212\ : InMux
    port map (
            O => \N__15832\,
            I => \N__15783\
        );

    \I__3211\ : InMux
    port map (
            O => \N__15831\,
            I => \N__15783\
        );

    \I__3210\ : InMux
    port map (
            O => \N__15830\,
            I => \N__15783\
        );

    \I__3209\ : InMux
    port map (
            O => \N__15829\,
            I => \N__15783\
        );

    \I__3208\ : InMux
    port map (
            O => \N__15828\,
            I => \N__15783\
        );

    \I__3207\ : InMux
    port map (
            O => \N__15827\,
            I => \N__15783\
        );

    \I__3206\ : Span4Mux_h
    port map (
            O => \N__15824\,
            I => \N__15778\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__15817\,
            I => \N__15778\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__15810\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__3203\ : Odrv4
    port map (
            O => \N__15807\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__3202\ : Odrv4
    port map (
            O => \N__15800\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__15783\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__3200\ : Odrv4
    port map (
            O => \N__15778\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__3199\ : CascadeMux
    port map (
            O => \N__15767\,
            I => \N__15764\
        );

    \I__3198\ : InMux
    port map (
            O => \N__15764\,
            I => \N__15756\
        );

    \I__3197\ : InMux
    port map (
            O => \N__15763\,
            I => \N__15756\
        );

    \I__3196\ : InMux
    port map (
            O => \N__15762\,
            I => \N__15753\
        );

    \I__3195\ : InMux
    port map (
            O => \N__15761\,
            I => \N__15750\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__15756\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__15753\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__15750\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__3191\ : CascadeMux
    port map (
            O => \N__15743\,
            I => \N__15725\
        );

    \I__3190\ : CascadeMux
    port map (
            O => \N__15742\,
            I => \N__15722\
        );

    \I__3189\ : CascadeMux
    port map (
            O => \N__15741\,
            I => \N__15719\
        );

    \I__3188\ : CascadeMux
    port map (
            O => \N__15740\,
            I => \N__15716\
        );

    \I__3187\ : CascadeMux
    port map (
            O => \N__15739\,
            I => \N__15709\
        );

    \I__3186\ : CascadeMux
    port map (
            O => \N__15738\,
            I => \N__15706\
        );

    \I__3185\ : CascadeMux
    port map (
            O => \N__15737\,
            I => \N__15703\
        );

    \I__3184\ : CascadeMux
    port map (
            O => \N__15736\,
            I => \N__15700\
        );

    \I__3183\ : CascadeMux
    port map (
            O => \N__15735\,
            I => \N__15697\
        );

    \I__3182\ : CascadeMux
    port map (
            O => \N__15734\,
            I => \N__15694\
        );

    \I__3181\ : CascadeMux
    port map (
            O => \N__15733\,
            I => \N__15691\
        );

    \I__3180\ : CascadeMux
    port map (
            O => \N__15732\,
            I => \N__15688\
        );

    \I__3179\ : InMux
    port map (
            O => \N__15731\,
            I => \N__15669\
        );

    \I__3178\ : InMux
    port map (
            O => \N__15730\,
            I => \N__15669\
        );

    \I__3177\ : InMux
    port map (
            O => \N__15729\,
            I => \N__15669\
        );

    \I__3176\ : InMux
    port map (
            O => \N__15728\,
            I => \N__15669\
        );

    \I__3175\ : InMux
    port map (
            O => \N__15725\,
            I => \N__15669\
        );

    \I__3174\ : InMux
    port map (
            O => \N__15722\,
            I => \N__15669\
        );

    \I__3173\ : InMux
    port map (
            O => \N__15719\,
            I => \N__15669\
        );

    \I__3172\ : InMux
    port map (
            O => \N__15716\,
            I => \N__15669\
        );

    \I__3171\ : CascadeMux
    port map (
            O => \N__15715\,
            I => \N__15666\
        );

    \I__3170\ : InMux
    port map (
            O => \N__15714\,
            I => \N__15657\
        );

    \I__3169\ : InMux
    port map (
            O => \N__15713\,
            I => \N__15657\
        );

    \I__3168\ : InMux
    port map (
            O => \N__15712\,
            I => \N__15657\
        );

    \I__3167\ : InMux
    port map (
            O => \N__15709\,
            I => \N__15657\
        );

    \I__3166\ : InMux
    port map (
            O => \N__15706\,
            I => \N__15648\
        );

    \I__3165\ : InMux
    port map (
            O => \N__15703\,
            I => \N__15648\
        );

    \I__3164\ : InMux
    port map (
            O => \N__15700\,
            I => \N__15648\
        );

    \I__3163\ : InMux
    port map (
            O => \N__15697\,
            I => \N__15648\
        );

    \I__3162\ : InMux
    port map (
            O => \N__15694\,
            I => \N__15639\
        );

    \I__3161\ : InMux
    port map (
            O => \N__15691\,
            I => \N__15639\
        );

    \I__3160\ : InMux
    port map (
            O => \N__15688\,
            I => \N__15639\
        );

    \I__3159\ : InMux
    port map (
            O => \N__15687\,
            I => \N__15639\
        );

    \I__3158\ : CascadeMux
    port map (
            O => \N__15686\,
            I => \N__15636\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__15669\,
            I => \N__15633\
        );

    \I__3156\ : InMux
    port map (
            O => \N__15666\,
            I => \N__15630\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__15657\,
            I => \N__15627\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__15648\,
            I => \N__15621\
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__15639\,
            I => \N__15621\
        );

    \I__3152\ : InMux
    port map (
            O => \N__15636\,
            I => \N__15618\
        );

    \I__3151\ : Span4Mux_h
    port map (
            O => \N__15633\,
            I => \N__15615\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__15630\,
            I => \N__15610\
        );

    \I__3149\ : Span4Mux_v
    port map (
            O => \N__15627\,
            I => \N__15610\
        );

    \I__3148\ : InMux
    port map (
            O => \N__15626\,
            I => \N__15607\
        );

    \I__3147\ : Span4Mux_h
    port map (
            O => \N__15621\,
            I => \N__15604\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__15618\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__3145\ : Odrv4
    port map (
            O => \N__15615\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__3144\ : Odrv4
    port map (
            O => \N__15610\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__15607\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__3142\ : Odrv4
    port map (
            O => \N__15604\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__3141\ : InMux
    port map (
            O => \N__15593\,
            I => \N__15569\
        );

    \I__3140\ : InMux
    port map (
            O => \N__15592\,
            I => \N__15569\
        );

    \I__3139\ : InMux
    port map (
            O => \N__15591\,
            I => \N__15569\
        );

    \I__3138\ : InMux
    port map (
            O => \N__15590\,
            I => \N__15569\
        );

    \I__3137\ : InMux
    port map (
            O => \N__15589\,
            I => \N__15569\
        );

    \I__3136\ : InMux
    port map (
            O => \N__15588\,
            I => \N__15569\
        );

    \I__3135\ : InMux
    port map (
            O => \N__15587\,
            I => \N__15569\
        );

    \I__3134\ : InMux
    port map (
            O => \N__15586\,
            I => \N__15569\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__15569\,
            I => \N__15563\
        );

    \I__3132\ : InMux
    port map (
            O => \N__15568\,
            I => \N__15547\
        );

    \I__3131\ : InMux
    port map (
            O => \N__15567\,
            I => \N__15544\
        );

    \I__3130\ : InMux
    port map (
            O => \N__15566\,
            I => \N__15541\
        );

    \I__3129\ : Span4Mux_h
    port map (
            O => \N__15563\,
            I => \N__15538\
        );

    \I__3128\ : InMux
    port map (
            O => \N__15562\,
            I => \N__15529\
        );

    \I__3127\ : InMux
    port map (
            O => \N__15561\,
            I => \N__15529\
        );

    \I__3126\ : InMux
    port map (
            O => \N__15560\,
            I => \N__15529\
        );

    \I__3125\ : InMux
    port map (
            O => \N__15559\,
            I => \N__15529\
        );

    \I__3124\ : InMux
    port map (
            O => \N__15558\,
            I => \N__15514\
        );

    \I__3123\ : InMux
    port map (
            O => \N__15557\,
            I => \N__15514\
        );

    \I__3122\ : InMux
    port map (
            O => \N__15556\,
            I => \N__15514\
        );

    \I__3121\ : InMux
    port map (
            O => \N__15555\,
            I => \N__15514\
        );

    \I__3120\ : InMux
    port map (
            O => \N__15554\,
            I => \N__15514\
        );

    \I__3119\ : InMux
    port map (
            O => \N__15553\,
            I => \N__15514\
        );

    \I__3118\ : InMux
    port map (
            O => \N__15552\,
            I => \N__15514\
        );

    \I__3117\ : InMux
    port map (
            O => \N__15551\,
            I => \N__15511\
        );

    \I__3116\ : InMux
    port map (
            O => \N__15550\,
            I => \N__15508\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__15547\,
            I => \N__15505\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__15544\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__15541\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__3112\ : Odrv4
    port map (
            O => \N__15538\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__15529\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__15514\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__15511\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__15508\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__3107\ : Odrv4
    port map (
            O => \N__15505\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__3106\ : InMux
    port map (
            O => \N__15488\,
            I => \N__15485\
        );

    \I__3105\ : LocalMux
    port map (
            O => \N__15485\,
            I => \phase_controller_inst1.stoper_tr.N_60\
        );

    \I__3104\ : InMux
    port map (
            O => \N__15482\,
            I => \N__15478\
        );

    \I__3103\ : InMux
    port map (
            O => \N__15481\,
            I => \N__15474\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__15478\,
            I => \N__15471\
        );

    \I__3101\ : InMux
    port map (
            O => \N__15477\,
            I => \N__15468\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__15474\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__3099\ : Odrv4
    port map (
            O => \N__15471\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__15468\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__3097\ : InMux
    port map (
            O => \N__15461\,
            I => \N__15457\
        );

    \I__3096\ : InMux
    port map (
            O => \N__15460\,
            I => \N__15454\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__15457\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__15454\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__3093\ : IoInMux
    port map (
            O => \N__15449\,
            I => \N__15446\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__15446\,
            I => \N__15443\
        );

    \I__3091\ : Span4Mux_s1_v
    port map (
            O => \N__15443\,
            I => \N__15440\
        );

    \I__3090\ : Span4Mux_v
    port map (
            O => \N__15440\,
            I => \N__15437\
        );

    \I__3089\ : Odrv4
    port map (
            O => \N__15437\,
            I => \delay_measurement_inst.delay_tr_timer.N_181_i\
        );

    \I__3088\ : InMux
    port map (
            O => \N__15434\,
            I => \N__15425\
        );

    \I__3087\ : InMux
    port map (
            O => \N__15433\,
            I => \N__15425\
        );

    \I__3086\ : InMux
    port map (
            O => \N__15432\,
            I => \N__15425\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__15425\,
            I => \delay_measurement_inst.hc_prevZ0\
        );

    \I__3084\ : InMux
    port map (
            O => \N__15422\,
            I => \N__15416\
        );

    \I__3083\ : InMux
    port map (
            O => \N__15421\,
            I => \N__15409\
        );

    \I__3082\ : InMux
    port map (
            O => \N__15420\,
            I => \N__15409\
        );

    \I__3081\ : InMux
    port map (
            O => \N__15419\,
            I => \N__15409\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__15416\,
            I => \delay_measurement_inst.hc_syncZ0Z_1\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__15409\,
            I => \delay_measurement_inst.hc_syncZ0Z_1\
        );

    \I__3078\ : InMux
    port map (
            O => \N__15404\,
            I => \N__15401\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__15401\,
            I => \N__15397\
        );

    \I__3076\ : InMux
    port map (
            O => \N__15400\,
            I => \N__15394\
        );

    \I__3075\ : Odrv12
    port map (
            O => \N__15397\,
            I => \delay_measurement_inst.delay_hc_timer.N_81\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__15394\,
            I => \delay_measurement_inst.delay_hc_timer.N_81\
        );

    \I__3073\ : InMux
    port map (
            O => \N__15389\,
            I => \N__15385\
        );

    \I__3072\ : InMux
    port map (
            O => \N__15388\,
            I => \N__15382\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__15385\,
            I => \N__15378\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__15382\,
            I => \N__15375\
        );

    \I__3069\ : InMux
    port map (
            O => \N__15381\,
            I => \N__15372\
        );

    \I__3068\ : Odrv4
    port map (
            O => \N__15378\,
            I => \delay_measurement_inst.N_54\
        );

    \I__3067\ : Odrv4
    port map (
            O => \N__15375\,
            I => \delay_measurement_inst.N_54\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__15372\,
            I => \delay_measurement_inst.N_54\
        );

    \I__3065\ : InMux
    port map (
            O => \N__15365\,
            I => \N__15356\
        );

    \I__3064\ : InMux
    port map (
            O => \N__15364\,
            I => \N__15356\
        );

    \I__3063\ : InMux
    port map (
            O => \N__15363\,
            I => \N__15349\
        );

    \I__3062\ : InMux
    port map (
            O => \N__15362\,
            I => \N__15349\
        );

    \I__3061\ : InMux
    port map (
            O => \N__15361\,
            I => \N__15349\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__15356\,
            I => \delay_measurement_inst.N_132\
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__15349\,
            I => \delay_measurement_inst.N_132\
        );

    \I__3058\ : CascadeMux
    port map (
            O => \N__15344\,
            I => \N__15340\
        );

    \I__3057\ : InMux
    port map (
            O => \N__15343\,
            I => \N__15335\
        );

    \I__3056\ : InMux
    port map (
            O => \N__15340\,
            I => \N__15335\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__15335\,
            I => \delay_measurement_inst.N_139\
        );

    \I__3054\ : CascadeMux
    port map (
            O => \N__15332\,
            I => \N__15329\
        );

    \I__3053\ : InMux
    port map (
            O => \N__15329\,
            I => \N__15326\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__15326\,
            I => \N__15322\
        );

    \I__3051\ : InMux
    port map (
            O => \N__15325\,
            I => \N__15318\
        );

    \I__3050\ : Sp12to4
    port map (
            O => \N__15322\,
            I => \N__15315\
        );

    \I__3049\ : InMux
    port map (
            O => \N__15321\,
            I => \N__15312\
        );

    \I__3048\ : LocalMux
    port map (
            O => \N__15318\,
            I => \delay_measurement_inst.N_134_i\
        );

    \I__3047\ : Odrv12
    port map (
            O => \N__15315\,
            I => \delay_measurement_inst.N_134_i\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__15312\,
            I => \delay_measurement_inst.N_134_i\
        );

    \I__3045\ : CascadeMux
    port map (
            O => \N__15305\,
            I => \delay_measurement_inst.N_201_cascade_\
        );

    \I__3044\ : CascadeMux
    port map (
            O => \N__15302\,
            I => \N__15297\
        );

    \I__3043\ : InMux
    port map (
            O => \N__15301\,
            I => \N__15294\
        );

    \I__3042\ : InMux
    port map (
            O => \N__15300\,
            I => \N__15289\
        );

    \I__3041\ : InMux
    port map (
            O => \N__15297\,
            I => \N__15289\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__15294\,
            I => \delay_measurement_inst.delay_tr_timer.N_167\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__15289\,
            I => \delay_measurement_inst.delay_tr_timer.N_167\
        );

    \I__3038\ : CascadeMux
    port map (
            O => \N__15284\,
            I => \N__15276\
        );

    \I__3037\ : CascadeMux
    port map (
            O => \N__15283\,
            I => \N__15273\
        );

    \I__3036\ : CascadeMux
    port map (
            O => \N__15282\,
            I => \N__15269\
        );

    \I__3035\ : InMux
    port map (
            O => \N__15281\,
            I => \N__15264\
        );

    \I__3034\ : InMux
    port map (
            O => \N__15280\,
            I => \N__15264\
        );

    \I__3033\ : InMux
    port map (
            O => \N__15279\,
            I => \N__15259\
        );

    \I__3032\ : InMux
    port map (
            O => \N__15276\,
            I => \N__15259\
        );

    \I__3031\ : InMux
    port map (
            O => \N__15273\,
            I => \N__15252\
        );

    \I__3030\ : InMux
    port map (
            O => \N__15272\,
            I => \N__15252\
        );

    \I__3029\ : InMux
    port map (
            O => \N__15269\,
            I => \N__15252\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__15264\,
            I => \delay_measurement_inst.N_170\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__15259\,
            I => \delay_measurement_inst.N_170\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__15252\,
            I => \delay_measurement_inst.N_170\
        );

    \I__3025\ : CascadeMux
    port map (
            O => \N__15245\,
            I => \N__15240\
        );

    \I__3024\ : InMux
    port map (
            O => \N__15244\,
            I => \N__15237\
        );

    \I__3023\ : InMux
    port map (
            O => \N__15243\,
            I => \N__15234\
        );

    \I__3022\ : InMux
    port map (
            O => \N__15240\,
            I => \N__15231\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__15237\,
            I => \N__15226\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__15234\,
            I => \N__15226\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__15231\,
            I => \N__15223\
        );

    \I__3018\ : Span4Mux_v
    port map (
            O => \N__15226\,
            I => \N__15220\
        );

    \I__3017\ : Odrv12
    port map (
            O => \N__15223\,
            I => \il_min_comp1_D2\
        );

    \I__3016\ : Odrv4
    port map (
            O => \N__15220\,
            I => \il_min_comp1_D2\
        );

    \I__3015\ : InMux
    port map (
            O => \N__15215\,
            I => \N__15211\
        );

    \I__3014\ : InMux
    port map (
            O => \N__15214\,
            I => \N__15207\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__15211\,
            I => \N__15204\
        );

    \I__3012\ : InMux
    port map (
            O => \N__15210\,
            I => \N__15201\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__15207\,
            I => \N__15196\
        );

    \I__3010\ : Span12Mux_s10_h
    port map (
            O => \N__15204\,
            I => \N__15196\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__15201\,
            I => \phase_controller_inst1.T01_0_sqmuxa\
        );

    \I__3008\ : Odrv12
    port map (
            O => \N__15196\,
            I => \phase_controller_inst1.T01_0_sqmuxa\
        );

    \I__3007\ : InMux
    port map (
            O => \N__15191\,
            I => \N__15186\
        );

    \I__3006\ : InMux
    port map (
            O => \N__15190\,
            I => \N__15181\
        );

    \I__3005\ : InMux
    port map (
            O => \N__15189\,
            I => \N__15181\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__15186\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__15181\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__3002\ : IoInMux
    port map (
            O => \N__15176\,
            I => \N__15173\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__15173\,
            I => \N__15170\
        );

    \I__3000\ : Span4Mux_s2_v
    port map (
            O => \N__15170\,
            I => \N__15167\
        );

    \I__2999\ : Span4Mux_h
    port map (
            O => \N__15167\,
            I => \N__15163\
        );

    \I__2998\ : CascadeMux
    port map (
            O => \N__15166\,
            I => \N__15160\
        );

    \I__2997\ : Span4Mux_h
    port map (
            O => \N__15163\,
            I => \N__15157\
        );

    \I__2996\ : InMux
    port map (
            O => \N__15160\,
            I => \N__15154\
        );

    \I__2995\ : Odrv4
    port map (
            O => \N__15157\,
            I => \T12_c\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__15154\,
            I => \T12_c\
        );

    \I__2993\ : InMux
    port map (
            O => \N__15149\,
            I => \N__15146\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__15146\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_13\
        );

    \I__2991\ : CEMux
    port map (
            O => \N__15143\,
            I => \N__15138\
        );

    \I__2990\ : CEMux
    port map (
            O => \N__15142\,
            I => \N__15135\
        );

    \I__2989\ : CEMux
    port map (
            O => \N__15141\,
            I => \N__15132\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__15138\,
            I => \N__15129\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__15135\,
            I => \N__15126\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__15132\,
            I => \N__15123\
        );

    \I__2985\ : Span4Mux_v
    port map (
            O => \N__15129\,
            I => \N__15116\
        );

    \I__2984\ : Span4Mux_v
    port map (
            O => \N__15126\,
            I => \N__15116\
        );

    \I__2983\ : Span4Mux_v
    port map (
            O => \N__15123\,
            I => \N__15116\
        );

    \I__2982\ : Odrv4
    port map (
            O => \N__15116\,
            I => \phase_controller_slave.stoper_hc.stoper_state_RNI10KLZ0Z_1\
        );

    \I__2981\ : InMux
    port map (
            O => \N__15113\,
            I => \N__15108\
        );

    \I__2980\ : CascadeMux
    port map (
            O => \N__15112\,
            I => \N__15104\
        );

    \I__2979\ : InMux
    port map (
            O => \N__15111\,
            I => \N__15101\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__15108\,
            I => \N__15098\
        );

    \I__2977\ : InMux
    port map (
            O => \N__15107\,
            I => \N__15095\
        );

    \I__2976\ : InMux
    port map (
            O => \N__15104\,
            I => \N__15092\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__15101\,
            I => \N__15089\
        );

    \I__2974\ : Span4Mux_v
    port map (
            O => \N__15098\,
            I => \N__15082\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__15095\,
            I => \N__15082\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__15092\,
            I => \N__15082\
        );

    \I__2971\ : Span4Mux_h
    port map (
            O => \N__15089\,
            I => \N__15079\
        );

    \I__2970\ : Span4Mux_h
    port map (
            O => \N__15082\,
            I => \N__15076\
        );

    \I__2969\ : Odrv4
    port map (
            O => \N__15079\,
            I => measured_delay_tr_3
        );

    \I__2968\ : Odrv4
    port map (
            O => \N__15076\,
            I => measured_delay_tr_3
        );

    \I__2967\ : InMux
    port map (
            O => \N__15071\,
            I => \N__15068\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__15068\,
            I => \N__15063\
        );

    \I__2965\ : InMux
    port map (
            O => \N__15067\,
            I => \N__15060\
        );

    \I__2964\ : InMux
    port map (
            O => \N__15066\,
            I => \N__15057\
        );

    \I__2963\ : Span4Mux_v
    port map (
            O => \N__15063\,
            I => \N__15051\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__15060\,
            I => \N__15051\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__15057\,
            I => \N__15048\
        );

    \I__2960\ : InMux
    port map (
            O => \N__15056\,
            I => \N__15045\
        );

    \I__2959\ : Span4Mux_h
    port map (
            O => \N__15051\,
            I => \N__15042\
        );

    \I__2958\ : Span12Mux_s5_h
    port map (
            O => \N__15048\,
            I => \N__15037\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__15045\,
            I => \N__15037\
        );

    \I__2956\ : Odrv4
    port map (
            O => \N__15042\,
            I => measured_delay_tr_18
        );

    \I__2955\ : Odrv12
    port map (
            O => \N__15037\,
            I => measured_delay_tr_18
        );

    \I__2954\ : InMux
    port map (
            O => \N__15032\,
            I => \N__15029\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__15029\,
            I => \N__15025\
        );

    \I__2952\ : InMux
    port map (
            O => \N__15028\,
            I => \N__15022\
        );

    \I__2951\ : Span4Mux_v
    port map (
            O => \N__15025\,
            I => \N__15017\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__15022\,
            I => \N__15014\
        );

    \I__2949\ : InMux
    port map (
            O => \N__15021\,
            I => \N__15009\
        );

    \I__2948\ : InMux
    port map (
            O => \N__15020\,
            I => \N__15009\
        );

    \I__2947\ : Span4Mux_h
    port map (
            O => \N__15017\,
            I => \N__15004\
        );

    \I__2946\ : Span4Mux_v
    port map (
            O => \N__15014\,
            I => \N__15004\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__15009\,
            I => \N__15001\
        );

    \I__2944\ : Odrv4
    port map (
            O => \N__15004\,
            I => measured_delay_tr_4
        );

    \I__2943\ : Odrv4
    port map (
            O => \N__15001\,
            I => measured_delay_tr_4
        );

    \I__2942\ : InMux
    port map (
            O => \N__14996\,
            I => \N__14992\
        );

    \I__2941\ : CascadeMux
    port map (
            O => \N__14995\,
            I => \N__14984\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__14992\,
            I => \N__14980\
        );

    \I__2939\ : InMux
    port map (
            O => \N__14991\,
            I => \N__14977\
        );

    \I__2938\ : InMux
    port map (
            O => \N__14990\,
            I => \N__14970\
        );

    \I__2937\ : InMux
    port map (
            O => \N__14989\,
            I => \N__14970\
        );

    \I__2936\ : InMux
    port map (
            O => \N__14988\,
            I => \N__14970\
        );

    \I__2935\ : InMux
    port map (
            O => \N__14987\,
            I => \N__14963\
        );

    \I__2934\ : InMux
    port map (
            O => \N__14984\,
            I => \N__14963\
        );

    \I__2933\ : InMux
    port map (
            O => \N__14983\,
            I => \N__14963\
        );

    \I__2932\ : Span4Mux_v
    port map (
            O => \N__14980\,
            I => \N__14960\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__14977\,
            I => \delay_measurement_inst.N_129\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__14970\,
            I => \delay_measurement_inst.N_129\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__14963\,
            I => \delay_measurement_inst.N_129\
        );

    \I__2928\ : Odrv4
    port map (
            O => \N__14960\,
            I => \delay_measurement_inst.N_129\
        );

    \I__2927\ : InMux
    port map (
            O => \N__14951\,
            I => \N__14942\
        );

    \I__2926\ : InMux
    port map (
            O => \N__14950\,
            I => \N__14935\
        );

    \I__2925\ : InMux
    port map (
            O => \N__14949\,
            I => \N__14935\
        );

    \I__2924\ : InMux
    port map (
            O => \N__14948\,
            I => \N__14935\
        );

    \I__2923\ : InMux
    port map (
            O => \N__14947\,
            I => \N__14928\
        );

    \I__2922\ : InMux
    port map (
            O => \N__14946\,
            I => \N__14928\
        );

    \I__2921\ : InMux
    port map (
            O => \N__14945\,
            I => \N__14928\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__14942\,
            I => \N__14925\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__14935\,
            I => \delay_measurement_inst.N_172\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__14928\,
            I => \delay_measurement_inst.N_172\
        );

    \I__2917\ : Odrv4
    port map (
            O => \N__14925\,
            I => \delay_measurement_inst.N_172\
        );

    \I__2916\ : InMux
    port map (
            O => \N__14918\,
            I => \N__14915\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__14915\,
            I => \N__14911\
        );

    \I__2914\ : InMux
    port map (
            O => \N__14914\,
            I => \N__14908\
        );

    \I__2913\ : Span4Mux_h
    port map (
            O => \N__14911\,
            I => \N__14903\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__14908\,
            I => \N__14900\
        );

    \I__2911\ : InMux
    port map (
            O => \N__14907\,
            I => \N__14895\
        );

    \I__2910\ : InMux
    port map (
            O => \N__14906\,
            I => \N__14895\
        );

    \I__2909\ : Span4Mux_h
    port map (
            O => \N__14903\,
            I => \N__14892\
        );

    \I__2908\ : Span4Mux_v
    port map (
            O => \N__14900\,
            I => \N__14887\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__14895\,
            I => \N__14887\
        );

    \I__2906\ : Odrv4
    port map (
            O => \N__14892\,
            I => measured_delay_tr_2
        );

    \I__2905\ : Odrv4
    port map (
            O => \N__14887\,
            I => measured_delay_tr_2
        );

    \I__2904\ : CascadeMux
    port map (
            O => \N__14882\,
            I => \N__14878\
        );

    \I__2903\ : InMux
    port map (
            O => \N__14881\,
            I => \N__14875\
        );

    \I__2902\ : InMux
    port map (
            O => \N__14878\,
            I => \N__14872\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__14875\,
            I => \N__14869\
        );

    \I__2900\ : LocalMux
    port map (
            O => \N__14872\,
            I => \N__14866\
        );

    \I__2899\ : Span4Mux_h
    port map (
            O => \N__14869\,
            I => \N__14863\
        );

    \I__2898\ : Span4Mux_h
    port map (
            O => \N__14866\,
            I => \N__14857\
        );

    \I__2897\ : Span4Mux_v
    port map (
            O => \N__14863\,
            I => \N__14857\
        );

    \I__2896\ : InMux
    port map (
            O => \N__14862\,
            I => \N__14854\
        );

    \I__2895\ : Odrv4
    port map (
            O => \N__14857\,
            I => measured_delay_tr_10
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__14854\,
            I => measured_delay_tr_10
        );

    \I__2893\ : CascadeMux
    port map (
            O => \N__14849\,
            I => \N__14846\
        );

    \I__2892\ : InMux
    port map (
            O => \N__14846\,
            I => \N__14843\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__14843\,
            I => \N__14838\
        );

    \I__2890\ : InMux
    port map (
            O => \N__14842\,
            I => \N__14834\
        );

    \I__2889\ : InMux
    port map (
            O => \N__14841\,
            I => \N__14831\
        );

    \I__2888\ : Span4Mux_h
    port map (
            O => \N__14838\,
            I => \N__14828\
        );

    \I__2887\ : InMux
    port map (
            O => \N__14837\,
            I => \N__14825\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__14834\,
            I => \N__14822\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__14831\,
            I => \N__14819\
        );

    \I__2884\ : Span4Mux_v
    port map (
            O => \N__14828\,
            I => \N__14814\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__14825\,
            I => \N__14814\
        );

    \I__2882\ : Odrv12
    port map (
            O => \N__14822\,
            I => measured_delay_tr_11
        );

    \I__2881\ : Odrv4
    port map (
            O => \N__14819\,
            I => measured_delay_tr_11
        );

    \I__2880\ : Odrv4
    port map (
            O => \N__14814\,
            I => measured_delay_tr_11
        );

    \I__2879\ : CascadeMux
    port map (
            O => \N__14807\,
            I => \N__14803\
        );

    \I__2878\ : InMux
    port map (
            O => \N__14806\,
            I => \N__14800\
        );

    \I__2877\ : InMux
    port map (
            O => \N__14803\,
            I => \N__14797\
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__14800\,
            I => \N__14794\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__14797\,
            I => \N__14791\
        );

    \I__2874\ : Span4Mux_h
    port map (
            O => \N__14794\,
            I => \N__14788\
        );

    \I__2873\ : Span4Mux_h
    port map (
            O => \N__14791\,
            I => \N__14784\
        );

    \I__2872\ : Span4Mux_h
    port map (
            O => \N__14788\,
            I => \N__14781\
        );

    \I__2871\ : InMux
    port map (
            O => \N__14787\,
            I => \N__14778\
        );

    \I__2870\ : Odrv4
    port map (
            O => \N__14784\,
            I => measured_delay_tr_13
        );

    \I__2869\ : Odrv4
    port map (
            O => \N__14781\,
            I => measured_delay_tr_13
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__14778\,
            I => measured_delay_tr_13
        );

    \I__2867\ : InMux
    port map (
            O => \N__14771\,
            I => \N__14768\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__14768\,
            I => \delay_measurement_inst.delay_tr_timer.un1_reset_i_a2_6\
        );

    \I__2865\ : InMux
    port map (
            O => \N__14765\,
            I => \N__14762\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__14762\,
            I => \N__14759\
        );

    \I__2863\ : Odrv4
    port map (
            O => \N__14759\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_11\
        );

    \I__2862\ : InMux
    port map (
            O => \N__14756\,
            I => \N__14753\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__14753\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_7\
        );

    \I__2860\ : InMux
    port map (
            O => \N__14750\,
            I => \N__14747\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__14747\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_9\
        );

    \I__2858\ : InMux
    port map (
            O => \N__14744\,
            I => \N__14741\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__14741\,
            I => \N__14738\
        );

    \I__2856\ : Odrv4
    port map (
            O => \N__14738\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_10\
        );

    \I__2855\ : InMux
    port map (
            O => \N__14735\,
            I => \N__14732\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__14732\,
            I => \N__14729\
        );

    \I__2853\ : Odrv4
    port map (
            O => \N__14729\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_15\
        );

    \I__2852\ : InMux
    port map (
            O => \N__14726\,
            I => \N__14723\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__14723\,
            I => \N__14720\
        );

    \I__2850\ : Odrv4
    port map (
            O => \N__14720\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_14\
        );

    \I__2849\ : InMux
    port map (
            O => \N__14717\,
            I => \N__14714\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__14714\,
            I => \N__14711\
        );

    \I__2847\ : Odrv4
    port map (
            O => \N__14711\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_16\
        );

    \I__2846\ : InMux
    port map (
            O => \N__14708\,
            I => \N__14705\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__14705\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_17\
        );

    \I__2844\ : InMux
    port map (
            O => \N__14702\,
            I => \N__14699\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__14699\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_18\
        );

    \I__2842\ : CascadeMux
    port map (
            O => \N__14696\,
            I => \N__14693\
        );

    \I__2841\ : InMux
    port map (
            O => \N__14693\,
            I => \N__14690\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__14690\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\
        );

    \I__2839\ : InMux
    port map (
            O => \N__14687\,
            I => \N__14684\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__14684\,
            I => \N__14681\
        );

    \I__2837\ : Span4Mux_h
    port map (
            O => \N__14681\,
            I => \N__14678\
        );

    \I__2836\ : Odrv4
    port map (
            O => \N__14678\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\
        );

    \I__2835\ : CascadeMux
    port map (
            O => \N__14675\,
            I => \N__14672\
        );

    \I__2834\ : InMux
    port map (
            O => \N__14672\,
            I => \N__14669\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__14669\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_16\
        );

    \I__2832\ : InMux
    port map (
            O => \N__14666\,
            I => \N__14663\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__14663\,
            I => \N__14660\
        );

    \I__2830\ : Odrv4
    port map (
            O => \N__14660\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\
        );

    \I__2829\ : CascadeMux
    port map (
            O => \N__14657\,
            I => \N__14654\
        );

    \I__2828\ : InMux
    port map (
            O => \N__14654\,
            I => \N__14651\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__14651\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_17\
        );

    \I__2826\ : InMux
    port map (
            O => \N__14648\,
            I => \N__14645\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__14645\,
            I => \N__14642\
        );

    \I__2824\ : Odrv4
    port map (
            O => \N__14642\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\
        );

    \I__2823\ : CascadeMux
    port map (
            O => \N__14639\,
            I => \N__14636\
        );

    \I__2822\ : InMux
    port map (
            O => \N__14636\,
            I => \N__14633\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__14633\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_18\
        );

    \I__2820\ : InMux
    port map (
            O => \N__14630\,
            I => \N__14627\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__14627\,
            I => \N__14624\
        );

    \I__2818\ : Odrv4
    port map (
            O => \N__14624\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\
        );

    \I__2817\ : CascadeMux
    port map (
            O => \N__14621\,
            I => \N__14618\
        );

    \I__2816\ : InMux
    port map (
            O => \N__14618\,
            I => \N__14615\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__14615\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_19\
        );

    \I__2814\ : InMux
    port map (
            O => \N__14612\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__2813\ : InMux
    port map (
            O => \N__14609\,
            I => \N__14606\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__14606\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_12\
        );

    \I__2811\ : InMux
    port map (
            O => \N__14603\,
            I => \N__14600\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__14600\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_19\
        );

    \I__2809\ : CascadeMux
    port map (
            O => \N__14597\,
            I => \N__14594\
        );

    \I__2808\ : InMux
    port map (
            O => \N__14594\,
            I => \N__14591\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__14591\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\
        );

    \I__2806\ : InMux
    port map (
            O => \N__14588\,
            I => \N__14585\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__14585\,
            I => \N__14582\
        );

    \I__2804\ : Odrv4
    port map (
            O => \N__14582\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\
        );

    \I__2803\ : CascadeMux
    port map (
            O => \N__14579\,
            I => \N__14576\
        );

    \I__2802\ : InMux
    port map (
            O => \N__14576\,
            I => \N__14573\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__14573\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\
        );

    \I__2800\ : InMux
    port map (
            O => \N__14570\,
            I => \N__14567\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__14567\,
            I => \N__14564\
        );

    \I__2798\ : Odrv4
    port map (
            O => \N__14564\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\
        );

    \I__2797\ : CascadeMux
    port map (
            O => \N__14561\,
            I => \N__14558\
        );

    \I__2796\ : InMux
    port map (
            O => \N__14558\,
            I => \N__14555\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__14555\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\
        );

    \I__2794\ : CascadeMux
    port map (
            O => \N__14552\,
            I => \N__14549\
        );

    \I__2793\ : InMux
    port map (
            O => \N__14549\,
            I => \N__14546\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__14546\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\
        );

    \I__2791\ : CascadeMux
    port map (
            O => \N__14543\,
            I => \N__14540\
        );

    \I__2790\ : InMux
    port map (
            O => \N__14540\,
            I => \N__14537\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__14537\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\
        );

    \I__2788\ : CascadeMux
    port map (
            O => \N__14534\,
            I => \N__14531\
        );

    \I__2787\ : InMux
    port map (
            O => \N__14531\,
            I => \N__14528\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__14528\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\
        );

    \I__2785\ : CascadeMux
    port map (
            O => \N__14525\,
            I => \N__14522\
        );

    \I__2784\ : InMux
    port map (
            O => \N__14522\,
            I => \N__14519\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__14519\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\
        );

    \I__2782\ : CascadeMux
    port map (
            O => \N__14516\,
            I => \N__14513\
        );

    \I__2781\ : InMux
    port map (
            O => \N__14513\,
            I => \N__14510\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__14510\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\
        );

    \I__2779\ : CascadeMux
    port map (
            O => \N__14507\,
            I => \N__14504\
        );

    \I__2778\ : InMux
    port map (
            O => \N__14504\,
            I => \N__14501\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__14501\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\
        );

    \I__2776\ : InMux
    port map (
            O => \N__14498\,
            I => \N__14495\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__14495\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\
        );

    \I__2774\ : CascadeMux
    port map (
            O => \N__14492\,
            I => \N__14489\
        );

    \I__2773\ : InMux
    port map (
            O => \N__14489\,
            I => \N__14486\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__14486\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\
        );

    \I__2771\ : InMux
    port map (
            O => \N__14483\,
            I => \N__14480\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__14480\,
            I => \N__14477\
        );

    \I__2769\ : Odrv4
    port map (
            O => \N__14477\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\
        );

    \I__2768\ : CascadeMux
    port map (
            O => \N__14474\,
            I => \N__14471\
        );

    \I__2767\ : InMux
    port map (
            O => \N__14471\,
            I => \N__14468\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__14468\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\
        );

    \I__2765\ : InMux
    port map (
            O => \N__14465\,
            I => \N__14462\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__14462\,
            I => \N__14459\
        );

    \I__2763\ : Odrv4
    port map (
            O => \N__14459\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\
        );

    \I__2762\ : CascadeMux
    port map (
            O => \N__14456\,
            I => \N__14453\
        );

    \I__2761\ : InMux
    port map (
            O => \N__14453\,
            I => \N__14450\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__14450\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\
        );

    \I__2759\ : InMux
    port map (
            O => \N__14447\,
            I => \N__14444\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__14444\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\
        );

    \I__2757\ : CascadeMux
    port map (
            O => \N__14441\,
            I => \N__14438\
        );

    \I__2756\ : InMux
    port map (
            O => \N__14438\,
            I => \N__14435\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__14435\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\
        );

    \I__2754\ : InMux
    port map (
            O => \N__14432\,
            I => \N__14429\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__14429\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\
        );

    \I__2752\ : CascadeMux
    port map (
            O => \N__14426\,
            I => \N__14423\
        );

    \I__2751\ : InMux
    port map (
            O => \N__14423\,
            I => \N__14420\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__14420\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\
        );

    \I__2749\ : CascadeMux
    port map (
            O => \N__14417\,
            I => \N__14414\
        );

    \I__2748\ : InMux
    port map (
            O => \N__14414\,
            I => \N__14411\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__14411\,
            I => \N__14407\
        );

    \I__2746\ : InMux
    port map (
            O => \N__14410\,
            I => \N__14404\
        );

    \I__2745\ : Odrv12
    port map (
            O => \N__14407\,
            I => \delay_measurement_inst.elapsed_time_hc_4\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__14404\,
            I => \delay_measurement_inst.elapsed_time_hc_4\
        );

    \I__2743\ : CascadeMux
    port map (
            O => \N__14399\,
            I => \N__14394\
        );

    \I__2742\ : InMux
    port map (
            O => \N__14398\,
            I => \N__14391\
        );

    \I__2741\ : InMux
    port map (
            O => \N__14397\,
            I => \N__14386\
        );

    \I__2740\ : InMux
    port map (
            O => \N__14394\,
            I => \N__14386\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__14391\,
            I => \N__14383\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__14386\,
            I => \N__14380\
        );

    \I__2737\ : Span4Mux_h
    port map (
            O => \N__14383\,
            I => \N__14377\
        );

    \I__2736\ : Span4Mux_h
    port map (
            O => \N__14380\,
            I => \N__14374\
        );

    \I__2735\ : Odrv4
    port map (
            O => \N__14377\,
            I => \delay_measurement_inst.elapsed_time_hc_18\
        );

    \I__2734\ : Odrv4
    port map (
            O => \N__14374\,
            I => \delay_measurement_inst.elapsed_time_hc_18\
        );

    \I__2733\ : InMux
    port map (
            O => \N__14369\,
            I => \N__14366\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__14366\,
            I => \N__14361\
        );

    \I__2731\ : InMux
    port map (
            O => \N__14365\,
            I => \N__14356\
        );

    \I__2730\ : InMux
    port map (
            O => \N__14364\,
            I => \N__14356\
        );

    \I__2729\ : Span4Mux_h
    port map (
            O => \N__14361\,
            I => \N__14353\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__14356\,
            I => \N__14350\
        );

    \I__2727\ : Odrv4
    port map (
            O => \N__14353\,
            I => \delay_measurement_inst.elapsed_time_hc_17\
        );

    \I__2726\ : Odrv4
    port map (
            O => \N__14350\,
            I => \delay_measurement_inst.elapsed_time_hc_17\
        );

    \I__2725\ : InMux
    port map (
            O => \N__14345\,
            I => \N__14342\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__14342\,
            I => \N__14338\
        );

    \I__2723\ : InMux
    port map (
            O => \N__14341\,
            I => \N__14335\
        );

    \I__2722\ : Odrv4
    port map (
            O => \N__14338\,
            I => \delay_measurement_inst.elapsed_time_hc_6\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__14335\,
            I => \delay_measurement_inst.elapsed_time_hc_6\
        );

    \I__2720\ : InMux
    port map (
            O => \N__14330\,
            I => \N__14327\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__14327\,
            I => \N__14323\
        );

    \I__2718\ : CascadeMux
    port map (
            O => \N__14326\,
            I => \N__14320\
        );

    \I__2717\ : Span4Mux_h
    port map (
            O => \N__14323\,
            I => \N__14317\
        );

    \I__2716\ : InMux
    port map (
            O => \N__14320\,
            I => \N__14314\
        );

    \I__2715\ : Span4Mux_h
    port map (
            O => \N__14317\,
            I => \N__14311\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__14314\,
            I => \N__14308\
        );

    \I__2713\ : Odrv4
    port map (
            O => \N__14311\,
            I => \delay_measurement_inst.elapsed_time_hc_13\
        );

    \I__2712\ : Odrv4
    port map (
            O => \N__14308\,
            I => \delay_measurement_inst.elapsed_time_hc_13\
        );

    \I__2711\ : CascadeMux
    port map (
            O => \N__14303\,
            I => \N__14296\
        );

    \I__2710\ : InMux
    port map (
            O => \N__14302\,
            I => \N__14287\
        );

    \I__2709\ : InMux
    port map (
            O => \N__14301\,
            I => \N__14287\
        );

    \I__2708\ : InMux
    port map (
            O => \N__14300\,
            I => \N__14287\
        );

    \I__2707\ : InMux
    port map (
            O => \N__14299\,
            I => \N__14287\
        );

    \I__2706\ : InMux
    port map (
            O => \N__14296\,
            I => \N__14284\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__14287\,
            I => \N__14280\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__14284\,
            I => \N__14276\
        );

    \I__2703\ : InMux
    port map (
            O => \N__14283\,
            I => \N__14273\
        );

    \I__2702\ : Span4Mux_h
    port map (
            O => \N__14280\,
            I => \N__14270\
        );

    \I__2701\ : InMux
    port map (
            O => \N__14279\,
            I => \N__14267\
        );

    \I__2700\ : Odrv4
    port map (
            O => \N__14276\,
            I => \delay_measurement_inst.N_109\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__14273\,
            I => \delay_measurement_inst.N_109\
        );

    \I__2698\ : Odrv4
    port map (
            O => \N__14270\,
            I => \delay_measurement_inst.N_109\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__14267\,
            I => \delay_measurement_inst.N_109\
        );

    \I__2696\ : InMux
    port map (
            O => \N__14258\,
            I => \N__14242\
        );

    \I__2695\ : InMux
    port map (
            O => \N__14257\,
            I => \N__14242\
        );

    \I__2694\ : InMux
    port map (
            O => \N__14256\,
            I => \N__14242\
        );

    \I__2693\ : InMux
    port map (
            O => \N__14255\,
            I => \N__14242\
        );

    \I__2692\ : InMux
    port map (
            O => \N__14254\,
            I => \N__14237\
        );

    \I__2691\ : InMux
    port map (
            O => \N__14253\,
            I => \N__14237\
        );

    \I__2690\ : InMux
    port map (
            O => \N__14252\,
            I => \N__14232\
        );

    \I__2689\ : InMux
    port map (
            O => \N__14251\,
            I => \N__14232\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__14242\,
            I => \delay_measurement_inst.N_45\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__14237\,
            I => \delay_measurement_inst.N_45\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__14232\,
            I => \delay_measurement_inst.N_45\
        );

    \I__2685\ : CascadeMux
    port map (
            O => \N__14225\,
            I => \N__14219\
        );

    \I__2684\ : CascadeMux
    port map (
            O => \N__14224\,
            I => \N__14216\
        );

    \I__2683\ : CascadeMux
    port map (
            O => \N__14223\,
            I => \N__14212\
        );

    \I__2682\ : InMux
    port map (
            O => \N__14222\,
            I => \N__14201\
        );

    \I__2681\ : InMux
    port map (
            O => \N__14219\,
            I => \N__14201\
        );

    \I__2680\ : InMux
    port map (
            O => \N__14216\,
            I => \N__14201\
        );

    \I__2679\ : InMux
    port map (
            O => \N__14215\,
            I => \N__14201\
        );

    \I__2678\ : InMux
    port map (
            O => \N__14212\,
            I => \N__14196\
        );

    \I__2677\ : InMux
    port map (
            O => \N__14211\,
            I => \N__14196\
        );

    \I__2676\ : InMux
    port map (
            O => \N__14210\,
            I => \N__14193\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__14201\,
            I => \delay_measurement_inst.N_107\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__14196\,
            I => \delay_measurement_inst.N_107\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__14193\,
            I => \delay_measurement_inst.N_107\
        );

    \I__2672\ : InMux
    port map (
            O => \N__14186\,
            I => \N__14183\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__14183\,
            I => \N__14179\
        );

    \I__2670\ : InMux
    port map (
            O => \N__14182\,
            I => \N__14176\
        );

    \I__2669\ : Odrv4
    port map (
            O => \N__14179\,
            I => \delay_measurement_inst.elapsed_time_hc_5\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__14176\,
            I => \delay_measurement_inst.elapsed_time_hc_5\
        );

    \I__2667\ : CascadeMux
    port map (
            O => \N__14171\,
            I => \N__14168\
        );

    \I__2666\ : InMux
    port map (
            O => \N__14168\,
            I => \N__14163\
        );

    \I__2665\ : InMux
    port map (
            O => \N__14167\,
            I => \N__14158\
        );

    \I__2664\ : InMux
    port map (
            O => \N__14166\,
            I => \N__14158\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__14163\,
            I => \delay_measurement_inst.tr_stateZ0Z_0\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__14158\,
            I => \delay_measurement_inst.tr_stateZ0Z_0\
        );

    \I__2661\ : InMux
    port map (
            O => \N__14153\,
            I => \N__14148\
        );

    \I__2660\ : InMux
    port map (
            O => \N__14152\,
            I => \N__14143\
        );

    \I__2659\ : InMux
    port map (
            O => \N__14151\,
            I => \N__14143\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__14148\,
            I => \delay_measurement_inst.tr_prevZ0\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__14143\,
            I => \delay_measurement_inst.tr_prevZ0\
        );

    \I__2656\ : CascadeMux
    port map (
            O => \N__14138\,
            I => \N__14134\
        );

    \I__2655\ : CascadeMux
    port map (
            O => \N__14137\,
            I => \N__14131\
        );

    \I__2654\ : InMux
    port map (
            O => \N__14134\,
            I => \N__14123\
        );

    \I__2653\ : InMux
    port map (
            O => \N__14131\,
            I => \N__14123\
        );

    \I__2652\ : InMux
    port map (
            O => \N__14130\,
            I => \N__14123\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__14123\,
            I => \delay_measurement_inst.hc_stateZ0Z_0\
        );

    \I__2650\ : InMux
    port map (
            O => \N__14120\,
            I => \N__14117\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__14117\,
            I => \N__14111\
        );

    \I__2648\ : InMux
    port map (
            O => \N__14116\,
            I => \N__14108\
        );

    \I__2647\ : InMux
    port map (
            O => \N__14115\,
            I => \N__14103\
        );

    \I__2646\ : InMux
    port map (
            O => \N__14114\,
            I => \N__14103\
        );

    \I__2645\ : Span4Mux_h
    port map (
            O => \N__14111\,
            I => \N__14100\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__14108\,
            I => \N__14095\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__14103\,
            I => \N__14095\
        );

    \I__2642\ : Odrv4
    port map (
            O => \N__14100\,
            I => \delay_measurement_inst.elapsed_time_hc_14\
        );

    \I__2641\ : Odrv4
    port map (
            O => \N__14095\,
            I => \delay_measurement_inst.elapsed_time_hc_14\
        );

    \I__2640\ : InMux
    port map (
            O => \N__14090\,
            I => \N__14087\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__14087\,
            I => \N__14083\
        );

    \I__2638\ : CascadeMux
    port map (
            O => \N__14086\,
            I => \N__14079\
        );

    \I__2637\ : Span4Mux_h
    port map (
            O => \N__14083\,
            I => \N__14076\
        );

    \I__2636\ : InMux
    port map (
            O => \N__14082\,
            I => \N__14073\
        );

    \I__2635\ : InMux
    port map (
            O => \N__14079\,
            I => \N__14070\
        );

    \I__2634\ : Odrv4
    port map (
            O => \N__14076\,
            I => \delay_measurement_inst.elapsed_time_hc_9\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__14073\,
            I => \delay_measurement_inst.elapsed_time_hc_9\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__14070\,
            I => \delay_measurement_inst.elapsed_time_hc_9\
        );

    \I__2631\ : InMux
    port map (
            O => \N__14063\,
            I => \N__14060\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__14060\,
            I => \N__14057\
        );

    \I__2629\ : Span4Mux_h
    port map (
            O => \N__14057\,
            I => \N__14053\
        );

    \I__2628\ : InMux
    port map (
            O => \N__14056\,
            I => \N__14050\
        );

    \I__2627\ : Odrv4
    port map (
            O => \N__14053\,
            I => \delay_measurement_inst.elapsed_time_hc_7\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__14050\,
            I => \delay_measurement_inst.elapsed_time_hc_7\
        );

    \I__2625\ : IoInMux
    port map (
            O => \N__14045\,
            I => \N__14042\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__14042\,
            I => \N__14038\
        );

    \I__2623\ : InMux
    port map (
            O => \N__14041\,
            I => \N__14035\
        );

    \I__2622\ : Span12Mux_s11_v
    port map (
            O => \N__14038\,
            I => \N__14032\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__14035\,
            I => \delay_measurement_inst.delay_hc_timer.N_32\
        );

    \I__2620\ : Odrv12
    port map (
            O => \N__14032\,
            I => \delay_measurement_inst.delay_hc_timer.N_32\
        );

    \I__2619\ : InMux
    port map (
            O => \N__14027\,
            I => \N__14018\
        );

    \I__2618\ : InMux
    port map (
            O => \N__14026\,
            I => \N__14018\
        );

    \I__2617\ : InMux
    port map (
            O => \N__14025\,
            I => \N__14018\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__14018\,
            I => \N__14015\
        );

    \I__2615\ : Odrv4
    port map (
            O => \N__14015\,
            I => \delay_measurement_inst.N_54_i\
        );

    \I__2614\ : InMux
    port map (
            O => \N__14012\,
            I => \N__14009\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__14009\,
            I => \N__14006\
        );

    \I__2612\ : Span4Mux_h
    port map (
            O => \N__14006\,
            I => \N__14002\
        );

    \I__2611\ : InMux
    port map (
            O => \N__14005\,
            I => \N__13999\
        );

    \I__2610\ : Odrv4
    port map (
            O => \N__14002\,
            I => \delay_measurement_inst.elapsed_time_hc_8\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__13999\,
            I => \delay_measurement_inst.elapsed_time_hc_8\
        );

    \I__2608\ : CascadeMux
    port map (
            O => \N__13994\,
            I => \N__13991\
        );

    \I__2607\ : InMux
    port map (
            O => \N__13991\,
            I => \N__13988\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__13988\,
            I => \N__13985\
        );

    \I__2605\ : Span4Mux_h
    port map (
            O => \N__13985\,
            I => \N__13982\
        );

    \I__2604\ : Span4Mux_h
    port map (
            O => \N__13982\,
            I => \N__13979\
        );

    \I__2603\ : Odrv4
    port map (
            O => \N__13979\,
            I => \delay_measurement_inst.elapsed_time_hc_1\
        );

    \I__2602\ : InMux
    port map (
            O => \N__13976\,
            I => \N__13973\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__13973\,
            I => \N__13969\
        );

    \I__2600\ : InMux
    port map (
            O => \N__13972\,
            I => \N__13966\
        );

    \I__2599\ : Odrv4
    port map (
            O => \N__13969\,
            I => \delay_measurement_inst.elapsed_time_hc_10\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__13966\,
            I => \delay_measurement_inst.elapsed_time_hc_10\
        );

    \I__2597\ : InMux
    port map (
            O => \N__13961\,
            I => \N__13958\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__13958\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\
        );

    \I__2595\ : InMux
    port map (
            O => \N__13955\,
            I => \N__13952\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__13952\,
            I => \N__13948\
        );

    \I__2593\ : InMux
    port map (
            O => \N__13951\,
            I => \N__13945\
        );

    \I__2592\ : Span4Mux_h
    port map (
            O => \N__13948\,
            I => \N__13942\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__13945\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__2590\ : Odrv4
    port map (
            O => \N__13942\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__2589\ : InMux
    port map (
            O => \N__13937\,
            I => \N__13934\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__13934\,
            I => \N__13931\
        );

    \I__2587\ : Span4Mux_s3_v
    port map (
            O => \N__13931\,
            I => \N__13927\
        );

    \I__2586\ : CascadeMux
    port map (
            O => \N__13930\,
            I => \N__13924\
        );

    \I__2585\ : Span4Mux_v
    port map (
            O => \N__13927\,
            I => \N__13920\
        );

    \I__2584\ : InMux
    port map (
            O => \N__13924\,
            I => \N__13917\
        );

    \I__2583\ : InMux
    port map (
            O => \N__13923\,
            I => \N__13913\
        );

    \I__2582\ : Span4Mux_v
    port map (
            O => \N__13920\,
            I => \N__13910\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__13917\,
            I => \N__13907\
        );

    \I__2580\ : InMux
    port map (
            O => \N__13916\,
            I => \N__13904\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__13913\,
            I => \N__13901\
        );

    \I__2578\ : Odrv4
    port map (
            O => \N__13910\,
            I => \phase_controller_slave.stateZ0Z_3\
        );

    \I__2577\ : Odrv4
    port map (
            O => \N__13907\,
            I => \phase_controller_slave.stateZ0Z_3\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__13904\,
            I => \phase_controller_slave.stateZ0Z_3\
        );

    \I__2575\ : Odrv12
    port map (
            O => \N__13901\,
            I => \phase_controller_slave.stateZ0Z_3\
        );

    \I__2574\ : IoInMux
    port map (
            O => \N__13892\,
            I => \N__13889\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__13889\,
            I => s3_phy_c
        );

    \I__2572\ : CascadeMux
    port map (
            O => \N__13886\,
            I => \delay_measurement_inst.N_54_cascade_\
        );

    \I__2571\ : InMux
    port map (
            O => \N__13883\,
            I => \N__13877\
        );

    \I__2570\ : InMux
    port map (
            O => \N__13882\,
            I => \N__13874\
        );

    \I__2569\ : InMux
    port map (
            O => \N__13881\,
            I => \N__13869\
        );

    \I__2568\ : InMux
    port map (
            O => \N__13880\,
            I => \N__13869\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__13877\,
            I => \delay_measurement_inst.tr_syncZ0Z_1\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__13874\,
            I => \delay_measurement_inst.tr_syncZ0Z_1\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__13869\,
            I => \delay_measurement_inst.tr_syncZ0Z_1\
        );

    \I__2564\ : CascadeMux
    port map (
            O => \N__13862\,
            I => \delay_measurement_inst.delay_tr_timer.un1_reset_i_a2_5_cascade_\
        );

    \I__2563\ : CascadeMux
    port map (
            O => \N__13859\,
            I => \delay_measurement_inst.delay_tr_timer.un1_reset_i_a2_9_cascade_\
        );

    \I__2562\ : CascadeMux
    port map (
            O => \N__13856\,
            I => \delay_measurement_inst.delay_tr_timer.N_160_cascade_\
        );

    \I__2561\ : InMux
    port map (
            O => \N__13853\,
            I => \N__13845\
        );

    \I__2560\ : InMux
    port map (
            O => \N__13852\,
            I => \N__13845\
        );

    \I__2559\ : InMux
    port map (
            O => \N__13851\,
            I => \N__13842\
        );

    \I__2558\ : InMux
    port map (
            O => \N__13850\,
            I => \N__13839\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__13845\,
            I => \N__13834\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__13842\,
            I => \N__13834\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__13839\,
            I => \N__13831\
        );

    \I__2554\ : Span12Mux_v
    port map (
            O => \N__13834\,
            I => \N__13828\
        );

    \I__2553\ : Odrv4
    port map (
            O => \N__13831\,
            I => \delay_measurement_inst.tr_state_RNIVV8GZ0Z_0\
        );

    \I__2552\ : Odrv12
    port map (
            O => \N__13828\,
            I => \delay_measurement_inst.tr_state_RNIVV8GZ0Z_0\
        );

    \I__2551\ : InMux
    port map (
            O => \N__13823\,
            I => \N__13820\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__13820\,
            I => \delay_measurement_inst.delay_tr_timer.un1_reset_i_0\
        );

    \I__2549\ : InMux
    port map (
            O => \N__13817\,
            I => \N__13813\
        );

    \I__2548\ : InMux
    port map (
            O => \N__13816\,
            I => \N__13810\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__13813\,
            I => \phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_2\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__13810\,
            I => \phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_2\
        );

    \I__2545\ : CascadeMux
    port map (
            O => \N__13805\,
            I => \N__13802\
        );

    \I__2544\ : InMux
    port map (
            O => \N__13802\,
            I => \N__13799\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__13799\,
            I => \N__13795\
        );

    \I__2542\ : CascadeMux
    port map (
            O => \N__13798\,
            I => \N__13789\
        );

    \I__2541\ : Span4Mux_h
    port map (
            O => \N__13795\,
            I => \N__13786\
        );

    \I__2540\ : InMux
    port map (
            O => \N__13794\,
            I => \N__13783\
        );

    \I__2539\ : InMux
    port map (
            O => \N__13793\,
            I => \N__13780\
        );

    \I__2538\ : InMux
    port map (
            O => \N__13792\,
            I => \N__13777\
        );

    \I__2537\ : InMux
    port map (
            O => \N__13789\,
            I => \N__13774\
        );

    \I__2536\ : Span4Mux_h
    port map (
            O => \N__13786\,
            I => \N__13769\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__13783\,
            I => \N__13769\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__13780\,
            I => measured_delay_tr_7
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__13777\,
            I => measured_delay_tr_7
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__13774\,
            I => measured_delay_tr_7
        );

    \I__2531\ : Odrv4
    port map (
            O => \N__13769\,
            I => measured_delay_tr_7
        );

    \I__2530\ : InMux
    port map (
            O => \N__13760\,
            I => \N__13757\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__13757\,
            I => \N__13754\
        );

    \I__2528\ : Span4Mux_h
    port map (
            O => \N__13754\,
            I => \N__13749\
        );

    \I__2527\ : InMux
    port map (
            O => \N__13753\,
            I => \N__13743\
        );

    \I__2526\ : InMux
    port map (
            O => \N__13752\,
            I => \N__13743\
        );

    \I__2525\ : Span4Mux_h
    port map (
            O => \N__13749\,
            I => \N__13740\
        );

    \I__2524\ : InMux
    port map (
            O => \N__13748\,
            I => \N__13737\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__13743\,
            I => \N__13734\
        );

    \I__2522\ : Odrv4
    port map (
            O => \N__13740\,
            I => measured_delay_tr_16
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__13737\,
            I => measured_delay_tr_16
        );

    \I__2520\ : Odrv4
    port map (
            O => \N__13734\,
            I => measured_delay_tr_16
        );

    \I__2519\ : InMux
    port map (
            O => \N__13727\,
            I => \N__13722\
        );

    \I__2518\ : CascadeMux
    port map (
            O => \N__13726\,
            I => \N__13719\
        );

    \I__2517\ : InMux
    port map (
            O => \N__13725\,
            I => \N__13715\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__13722\,
            I => \N__13709\
        );

    \I__2515\ : InMux
    port map (
            O => \N__13719\,
            I => \N__13704\
        );

    \I__2514\ : InMux
    port map (
            O => \N__13718\,
            I => \N__13704\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__13715\,
            I => \N__13701\
        );

    \I__2512\ : InMux
    port map (
            O => \N__13714\,
            I => \N__13698\
        );

    \I__2511\ : InMux
    port map (
            O => \N__13713\,
            I => \N__13695\
        );

    \I__2510\ : InMux
    port map (
            O => \N__13712\,
            I => \N__13692\
        );

    \I__2509\ : Span4Mux_v
    port map (
            O => \N__13709\,
            I => \N__13688\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__13704\,
            I => \N__13684\
        );

    \I__2507\ : Span4Mux_h
    port map (
            O => \N__13701\,
            I => \N__13677\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__13698\,
            I => \N__13677\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__13695\,
            I => \N__13677\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__13692\,
            I => \N__13674\
        );

    \I__2503\ : InMux
    port map (
            O => \N__13691\,
            I => \N__13671\
        );

    \I__2502\ : Span4Mux_h
    port map (
            O => \N__13688\,
            I => \N__13668\
        );

    \I__2501\ : InMux
    port map (
            O => \N__13687\,
            I => \N__13665\
        );

    \I__2500\ : Span4Mux_h
    port map (
            O => \N__13684\,
            I => \N__13656\
        );

    \I__2499\ : Span4Mux_v
    port map (
            O => \N__13677\,
            I => \N__13656\
        );

    \I__2498\ : Span4Mux_v
    port map (
            O => \N__13674\,
            I => \N__13656\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__13671\,
            I => \N__13656\
        );

    \I__2496\ : Odrv4
    port map (
            O => \N__13668\,
            I => measured_delay_tr_15
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__13665\,
            I => measured_delay_tr_15
        );

    \I__2494\ : Odrv4
    port map (
            O => \N__13656\,
            I => measured_delay_tr_15
        );

    \I__2493\ : InMux
    port map (
            O => \N__13649\,
            I => \N__13645\
        );

    \I__2492\ : InMux
    port map (
            O => \N__13648\,
            I => \N__13642\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__13645\,
            I => \N__13637\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__13642\,
            I => \N__13634\
        );

    \I__2489\ : InMux
    port map (
            O => \N__13641\,
            I => \N__13629\
        );

    \I__2488\ : InMux
    port map (
            O => \N__13640\,
            I => \N__13629\
        );

    \I__2487\ : Span12Mux_v
    port map (
            O => \N__13637\,
            I => \N__13626\
        );

    \I__2486\ : Span4Mux_h
    port map (
            O => \N__13634\,
            I => \N__13623\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__13629\,
            I => \N__13620\
        );

    \I__2484\ : Odrv12
    port map (
            O => \N__13626\,
            I => measured_delay_tr_6
        );

    \I__2483\ : Odrv4
    port map (
            O => \N__13623\,
            I => measured_delay_tr_6
        );

    \I__2482\ : Odrv4
    port map (
            O => \N__13620\,
            I => measured_delay_tr_6
        );

    \I__2481\ : InMux
    port map (
            O => \N__13613\,
            I => \N__13608\
        );

    \I__2480\ : InMux
    port map (
            O => \N__13612\,
            I => \N__13605\
        );

    \I__2479\ : InMux
    port map (
            O => \N__13611\,
            I => \N__13602\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__13608\,
            I => \N__13598\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__13605\,
            I => \N__13593\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__13602\,
            I => \N__13593\
        );

    \I__2475\ : InMux
    port map (
            O => \N__13601\,
            I => \N__13590\
        );

    \I__2474\ : Span4Mux_v
    port map (
            O => \N__13598\,
            I => \N__13583\
        );

    \I__2473\ : Span4Mux_h
    port map (
            O => \N__13593\,
            I => \N__13583\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__13590\,
            I => \N__13583\
        );

    \I__2471\ : Odrv4
    port map (
            O => \N__13583\,
            I => measured_delay_tr_12
        );

    \I__2470\ : InMux
    port map (
            O => \N__13580\,
            I => \N__13576\
        );

    \I__2469\ : InMux
    port map (
            O => \N__13579\,
            I => \N__13572\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__13576\,
            I => \N__13569\
        );

    \I__2467\ : InMux
    port map (
            O => \N__13575\,
            I => \N__13566\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__13572\,
            I => \N__13563\
        );

    \I__2465\ : Span4Mux_v
    port map (
            O => \N__13569\,
            I => \N__13558\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__13566\,
            I => \N__13558\
        );

    \I__2463\ : Span4Mux_v
    port map (
            O => \N__13563\,
            I => \N__13552\
        );

    \I__2462\ : Span4Mux_h
    port map (
            O => \N__13558\,
            I => \N__13552\
        );

    \I__2461\ : InMux
    port map (
            O => \N__13557\,
            I => \N__13549\
        );

    \I__2460\ : Odrv4
    port map (
            O => \N__13552\,
            I => measured_delay_tr_14
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__13549\,
            I => measured_delay_tr_14
        );

    \I__2458\ : CascadeMux
    port map (
            O => \N__13544\,
            I => \N__13541\
        );

    \I__2457\ : InMux
    port map (
            O => \N__13541\,
            I => \N__13538\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__13538\,
            I => \N__13534\
        );

    \I__2455\ : InMux
    port map (
            O => \N__13537\,
            I => \N__13531\
        );

    \I__2454\ : Span4Mux_h
    port map (
            O => \N__13534\,
            I => \N__13527\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__13531\,
            I => \N__13524\
        );

    \I__2452\ : InMux
    port map (
            O => \N__13530\,
            I => \N__13521\
        );

    \I__2451\ : Span4Mux_h
    port map (
            O => \N__13527\,
            I => \N__13518\
        );

    \I__2450\ : Span4Mux_v
    port map (
            O => \N__13524\,
            I => \N__13513\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__13521\,
            I => \N__13513\
        );

    \I__2448\ : Odrv4
    port map (
            O => \N__13518\,
            I => measured_delay_tr_1
        );

    \I__2447\ : Odrv4
    port map (
            O => \N__13513\,
            I => measured_delay_tr_1
        );

    \I__2446\ : InMux
    port map (
            O => \N__13508\,
            I => \N__13505\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__13505\,
            I => \N__13500\
        );

    \I__2444\ : InMux
    port map (
            O => \N__13504\,
            I => \N__13497\
        );

    \I__2443\ : CascadeMux
    port map (
            O => \N__13503\,
            I => \N__13493\
        );

    \I__2442\ : Span4Mux_h
    port map (
            O => \N__13500\,
            I => \N__13490\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__13497\,
            I => \N__13487\
        );

    \I__2440\ : InMux
    port map (
            O => \N__13496\,
            I => \N__13484\
        );

    \I__2439\ : InMux
    port map (
            O => \N__13493\,
            I => \N__13481\
        );

    \I__2438\ : Odrv4
    port map (
            O => \N__13490\,
            I => measured_delay_tr_17
        );

    \I__2437\ : Odrv4
    port map (
            O => \N__13487\,
            I => measured_delay_tr_17
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__13484\,
            I => measured_delay_tr_17
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__13481\,
            I => measured_delay_tr_17
        );

    \I__2434\ : InMux
    port map (
            O => \N__13472\,
            I => \N__13469\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__13469\,
            I => \N__13464\
        );

    \I__2432\ : InMux
    port map (
            O => \N__13468\,
            I => \N__13461\
        );

    \I__2431\ : InMux
    port map (
            O => \N__13467\,
            I => \N__13458\
        );

    \I__2430\ : Span4Mux_v
    port map (
            O => \N__13464\,
            I => \N__13453\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__13461\,
            I => \N__13450\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__13458\,
            I => \N__13447\
        );

    \I__2427\ : InMux
    port map (
            O => \N__13457\,
            I => \N__13444\
        );

    \I__2426\ : InMux
    port map (
            O => \N__13456\,
            I => \N__13441\
        );

    \I__2425\ : Odrv4
    port map (
            O => \N__13453\,
            I => measured_delay_tr_9
        );

    \I__2424\ : Odrv12
    port map (
            O => \N__13450\,
            I => measured_delay_tr_9
        );

    \I__2423\ : Odrv4
    port map (
            O => \N__13447\,
            I => measured_delay_tr_9
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__13444\,
            I => measured_delay_tr_9
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__13441\,
            I => measured_delay_tr_9
        );

    \I__2420\ : InMux
    port map (
            O => \N__13430\,
            I => \N__13427\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__13427\,
            I => \N__13423\
        );

    \I__2418\ : InMux
    port map (
            O => \N__13426\,
            I => \N__13420\
        );

    \I__2417\ : Span4Mux_v
    port map (
            O => \N__13423\,
            I => \N__13413\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__13420\,
            I => \N__13413\
        );

    \I__2415\ : InMux
    port map (
            O => \N__13419\,
            I => \N__13408\
        );

    \I__2414\ : InMux
    port map (
            O => \N__13418\,
            I => \N__13408\
        );

    \I__2413\ : Span4Mux_h
    port map (
            O => \N__13413\,
            I => \N__13405\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__13408\,
            I => \N__13402\
        );

    \I__2411\ : Odrv4
    port map (
            O => \N__13405\,
            I => measured_delay_tr_5
        );

    \I__2410\ : Odrv4
    port map (
            O => \N__13402\,
            I => measured_delay_tr_5
        );

    \I__2409\ : InMux
    port map (
            O => \N__13397\,
            I => \N__13393\
        );

    \I__2408\ : InMux
    port map (
            O => \N__13396\,
            I => \N__13390\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__13393\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__13390\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__2405\ : CascadeMux
    port map (
            O => \N__13385\,
            I => \N__13382\
        );

    \I__2404\ : InMux
    port map (
            O => \N__13382\,
            I => \N__13379\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__13379\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_15\
        );

    \I__2402\ : InMux
    port map (
            O => \N__13376\,
            I => \N__13372\
        );

    \I__2401\ : InMux
    port map (
            O => \N__13375\,
            I => \N__13369\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__13372\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__13369\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__2398\ : CascadeMux
    port map (
            O => \N__13364\,
            I => \N__13361\
        );

    \I__2397\ : InMux
    port map (
            O => \N__13361\,
            I => \N__13358\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__13358\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_16\
        );

    \I__2395\ : InMux
    port map (
            O => \N__13355\,
            I => \N__13351\
        );

    \I__2394\ : InMux
    port map (
            O => \N__13354\,
            I => \N__13348\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__13351\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__13348\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__2391\ : CascadeMux
    port map (
            O => \N__13343\,
            I => \N__13340\
        );

    \I__2390\ : InMux
    port map (
            O => \N__13340\,
            I => \N__13337\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__13337\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_17\
        );

    \I__2388\ : InMux
    port map (
            O => \N__13334\,
            I => \N__13330\
        );

    \I__2387\ : InMux
    port map (
            O => \N__13333\,
            I => \N__13327\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__13330\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__13327\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__2384\ : CascadeMux
    port map (
            O => \N__13322\,
            I => \N__13319\
        );

    \I__2383\ : InMux
    port map (
            O => \N__13319\,
            I => \N__13316\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__13316\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_18\
        );

    \I__2381\ : InMux
    port map (
            O => \N__13313\,
            I => \N__13309\
        );

    \I__2380\ : InMux
    port map (
            O => \N__13312\,
            I => \N__13306\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__13309\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__13306\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__2377\ : CascadeMux
    port map (
            O => \N__13301\,
            I => \N__13298\
        );

    \I__2376\ : InMux
    port map (
            O => \N__13298\,
            I => \N__13295\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__13295\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_19\
        );

    \I__2374\ : InMux
    port map (
            O => \N__13292\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__2373\ : CascadeMux
    port map (
            O => \N__13289\,
            I => \N__13278\
        );

    \I__2372\ : InMux
    port map (
            O => \N__13288\,
            I => \N__13275\
        );

    \I__2371\ : InMux
    port map (
            O => \N__13287\,
            I => \N__13256\
        );

    \I__2370\ : InMux
    port map (
            O => \N__13286\,
            I => \N__13256\
        );

    \I__2369\ : InMux
    port map (
            O => \N__13285\,
            I => \N__13256\
        );

    \I__2368\ : InMux
    port map (
            O => \N__13284\,
            I => \N__13256\
        );

    \I__2367\ : InMux
    port map (
            O => \N__13283\,
            I => \N__13256\
        );

    \I__2366\ : InMux
    port map (
            O => \N__13282\,
            I => \N__13256\
        );

    \I__2365\ : InMux
    port map (
            O => \N__13281\,
            I => \N__13256\
        );

    \I__2364\ : InMux
    port map (
            O => \N__13278\,
            I => \N__13245\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__13275\,
            I => \N__13242\
        );

    \I__2362\ : CascadeMux
    port map (
            O => \N__13274\,
            I => \N__13239\
        );

    \I__2361\ : InMux
    port map (
            O => \N__13273\,
            I => \N__13236\
        );

    \I__2360\ : CascadeMux
    port map (
            O => \N__13272\,
            I => \N__13233\
        );

    \I__2359\ : CascadeMux
    port map (
            O => \N__13271\,
            I => \N__13230\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__13256\,
            I => \N__13222\
        );

    \I__2357\ : InMux
    port map (
            O => \N__13255\,
            I => \N__13205\
        );

    \I__2356\ : InMux
    port map (
            O => \N__13254\,
            I => \N__13205\
        );

    \I__2355\ : InMux
    port map (
            O => \N__13253\,
            I => \N__13205\
        );

    \I__2354\ : InMux
    port map (
            O => \N__13252\,
            I => \N__13205\
        );

    \I__2353\ : InMux
    port map (
            O => \N__13251\,
            I => \N__13205\
        );

    \I__2352\ : InMux
    port map (
            O => \N__13250\,
            I => \N__13205\
        );

    \I__2351\ : InMux
    port map (
            O => \N__13249\,
            I => \N__13205\
        );

    \I__2350\ : InMux
    port map (
            O => \N__13248\,
            I => \N__13205\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__13245\,
            I => \N__13202\
        );

    \I__2348\ : Span4Mux_h
    port map (
            O => \N__13242\,
            I => \N__13199\
        );

    \I__2347\ : InMux
    port map (
            O => \N__13239\,
            I => \N__13196\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__13236\,
            I => \N__13193\
        );

    \I__2345\ : InMux
    port map (
            O => \N__13233\,
            I => \N__13178\
        );

    \I__2344\ : InMux
    port map (
            O => \N__13230\,
            I => \N__13178\
        );

    \I__2343\ : InMux
    port map (
            O => \N__13229\,
            I => \N__13178\
        );

    \I__2342\ : InMux
    port map (
            O => \N__13228\,
            I => \N__13178\
        );

    \I__2341\ : InMux
    port map (
            O => \N__13227\,
            I => \N__13178\
        );

    \I__2340\ : InMux
    port map (
            O => \N__13226\,
            I => \N__13178\
        );

    \I__2339\ : InMux
    port map (
            O => \N__13225\,
            I => \N__13178\
        );

    \I__2338\ : Odrv4
    port map (
            O => \N__13222\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__13205\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__2336\ : Odrv4
    port map (
            O => \N__13202\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__2335\ : Odrv4
    port map (
            O => \N__13199\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__13196\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__2333\ : Odrv4
    port map (
            O => \N__13193\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__13178\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__2331\ : InMux
    port map (
            O => \N__13163\,
            I => \N__13158\
        );

    \I__2330\ : InMux
    port map (
            O => \N__13162\,
            I => \N__13155\
        );

    \I__2329\ : InMux
    port map (
            O => \N__13161\,
            I => \N__13152\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__13158\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__13155\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__13152\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__2325\ : InMux
    port map (
            O => \N__13145\,
            I => \N__13142\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__13142\,
            I => \N__13134\
        );

    \I__2323\ : InMux
    port map (
            O => \N__13141\,
            I => \N__13131\
        );

    \I__2322\ : InMux
    port map (
            O => \N__13140\,
            I => \N__13122\
        );

    \I__2321\ : InMux
    port map (
            O => \N__13139\,
            I => \N__13122\
        );

    \I__2320\ : InMux
    port map (
            O => \N__13138\,
            I => \N__13122\
        );

    \I__2319\ : InMux
    port map (
            O => \N__13137\,
            I => \N__13122\
        );

    \I__2318\ : Odrv12
    port map (
            O => \N__13134\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__13131\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__13122\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__2315\ : CascadeMux
    port map (
            O => \N__13115\,
            I => \N__13112\
        );

    \I__2314\ : InMux
    port map (
            O => \N__13112\,
            I => \N__13109\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__13109\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0\
        );

    \I__2312\ : InMux
    port map (
            O => \N__13106\,
            I => \N__13103\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__13103\,
            I => \N__13100\
        );

    \I__2310\ : Span12Mux_v
    port map (
            O => \N__13100\,
            I => \N__13097\
        );

    \I__2309\ : Odrv12
    port map (
            O => \N__13097\,
            I => \il_min_comp1_D1\
        );

    \I__2308\ : InMux
    port map (
            O => \N__13094\,
            I => \N__13091\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__13091\,
            I => \N__13088\
        );

    \I__2306\ : Odrv4
    port map (
            O => \N__13088\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_8\
        );

    \I__2305\ : CascadeMux
    port map (
            O => \N__13085\,
            I => \N__13082\
        );

    \I__2304\ : InMux
    port map (
            O => \N__13082\,
            I => \N__13078\
        );

    \I__2303\ : InMux
    port map (
            O => \N__13081\,
            I => \N__13075\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__13078\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__13075\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__2300\ : CascadeMux
    port map (
            O => \N__13070\,
            I => \N__13067\
        );

    \I__2299\ : InMux
    port map (
            O => \N__13067\,
            I => \N__13064\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__13064\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_8\
        );

    \I__2297\ : InMux
    port map (
            O => \N__13061\,
            I => \N__13057\
        );

    \I__2296\ : InMux
    port map (
            O => \N__13060\,
            I => \N__13054\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__13057\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__13054\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__2293\ : CascadeMux
    port map (
            O => \N__13049\,
            I => \N__13046\
        );

    \I__2292\ : InMux
    port map (
            O => \N__13046\,
            I => \N__13043\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__13043\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_9\
        );

    \I__2290\ : InMux
    port map (
            O => \N__13040\,
            I => \N__13036\
        );

    \I__2289\ : InMux
    port map (
            O => \N__13039\,
            I => \N__13033\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__13036\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__13033\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__2286\ : CascadeMux
    port map (
            O => \N__13028\,
            I => \N__13025\
        );

    \I__2285\ : InMux
    port map (
            O => \N__13025\,
            I => \N__13022\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__13022\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_10\
        );

    \I__2283\ : InMux
    port map (
            O => \N__13019\,
            I => \N__13015\
        );

    \I__2282\ : InMux
    port map (
            O => \N__13018\,
            I => \N__13012\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__13015\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__13012\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__2279\ : CascadeMux
    port map (
            O => \N__13007\,
            I => \N__13004\
        );

    \I__2278\ : InMux
    port map (
            O => \N__13004\,
            I => \N__13001\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__13001\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_11\
        );

    \I__2276\ : InMux
    port map (
            O => \N__12998\,
            I => \N__12994\
        );

    \I__2275\ : InMux
    port map (
            O => \N__12997\,
            I => \N__12991\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__12994\,
            I => \N__12986\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__12991\,
            I => \N__12986\
        );

    \I__2272\ : Span4Mux_h
    port map (
            O => \N__12986\,
            I => \N__12983\
        );

    \I__2271\ : Odrv4
    port map (
            O => \N__12983\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__2270\ : CascadeMux
    port map (
            O => \N__12980\,
            I => \N__12977\
        );

    \I__2269\ : InMux
    port map (
            O => \N__12977\,
            I => \N__12974\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__12974\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_12\
        );

    \I__2267\ : InMux
    port map (
            O => \N__12971\,
            I => \N__12967\
        );

    \I__2266\ : InMux
    port map (
            O => \N__12970\,
            I => \N__12964\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__12967\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__12964\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__2263\ : CascadeMux
    port map (
            O => \N__12959\,
            I => \N__12956\
        );

    \I__2262\ : InMux
    port map (
            O => \N__12956\,
            I => \N__12953\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__12953\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_13\
        );

    \I__2260\ : InMux
    port map (
            O => \N__12950\,
            I => \N__12946\
        );

    \I__2259\ : InMux
    port map (
            O => \N__12949\,
            I => \N__12943\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__12946\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__12943\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__2256\ : CascadeMux
    port map (
            O => \N__12938\,
            I => \N__12935\
        );

    \I__2255\ : InMux
    port map (
            O => \N__12935\,
            I => \N__12932\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__12932\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_14\
        );

    \I__2253\ : InMux
    port map (
            O => \N__12929\,
            I => \N__12926\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__12926\,
            I => \N__12923\
        );

    \I__2251\ : Odrv4
    port map (
            O => \N__12923\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_1\
        );

    \I__2250\ : CascadeMux
    port map (
            O => \N__12920\,
            I => \N__12917\
        );

    \I__2249\ : InMux
    port map (
            O => \N__12917\,
            I => \N__12914\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__12914\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_1\
        );

    \I__2247\ : InMux
    port map (
            O => \N__12911\,
            I => \N__12908\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__12908\,
            I => \N__12905\
        );

    \I__2245\ : Odrv4
    port map (
            O => \N__12905\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_2\
        );

    \I__2244\ : InMux
    port map (
            O => \N__12902\,
            I => \N__12898\
        );

    \I__2243\ : InMux
    port map (
            O => \N__12901\,
            I => \N__12895\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__12898\,
            I => \N__12892\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__12895\,
            I => \N__12889\
        );

    \I__2240\ : Odrv4
    port map (
            O => \N__12892\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__2239\ : Odrv4
    port map (
            O => \N__12889\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__2238\ : CascadeMux
    port map (
            O => \N__12884\,
            I => \N__12881\
        );

    \I__2237\ : InMux
    port map (
            O => \N__12881\,
            I => \N__12878\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__12878\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_2\
        );

    \I__2235\ : InMux
    port map (
            O => \N__12875\,
            I => \N__12872\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__12872\,
            I => \N__12869\
        );

    \I__2233\ : Odrv4
    port map (
            O => \N__12869\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_3\
        );

    \I__2232\ : InMux
    port map (
            O => \N__12866\,
            I => \N__12863\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__12863\,
            I => \N__12859\
        );

    \I__2230\ : InMux
    port map (
            O => \N__12862\,
            I => \N__12856\
        );

    \I__2229\ : Odrv4
    port map (
            O => \N__12859\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__12856\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__2227\ : CascadeMux
    port map (
            O => \N__12851\,
            I => \N__12848\
        );

    \I__2226\ : InMux
    port map (
            O => \N__12848\,
            I => \N__12845\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__12845\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_3\
        );

    \I__2224\ : InMux
    port map (
            O => \N__12842\,
            I => \N__12839\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__12839\,
            I => \N__12836\
        );

    \I__2222\ : Odrv4
    port map (
            O => \N__12836\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_4\
        );

    \I__2221\ : InMux
    port map (
            O => \N__12833\,
            I => \N__12829\
        );

    \I__2220\ : InMux
    port map (
            O => \N__12832\,
            I => \N__12826\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__12829\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__12826\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__2217\ : CascadeMux
    port map (
            O => \N__12821\,
            I => \N__12818\
        );

    \I__2216\ : InMux
    port map (
            O => \N__12818\,
            I => \N__12815\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__12815\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_4\
        );

    \I__2214\ : InMux
    port map (
            O => \N__12812\,
            I => \N__12809\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__12809\,
            I => \N__12806\
        );

    \I__2212\ : Odrv4
    port map (
            O => \N__12806\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_5\
        );

    \I__2211\ : InMux
    port map (
            O => \N__12803\,
            I => \N__12799\
        );

    \I__2210\ : InMux
    port map (
            O => \N__12802\,
            I => \N__12796\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__12799\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__12796\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__2207\ : CascadeMux
    port map (
            O => \N__12791\,
            I => \N__12788\
        );

    \I__2206\ : InMux
    port map (
            O => \N__12788\,
            I => \N__12785\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__12785\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_5\
        );

    \I__2204\ : InMux
    port map (
            O => \N__12782\,
            I => \N__12779\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__12779\,
            I => \phase_controller_slave.stoper_hc.target_timeZ1Z_6\
        );

    \I__2202\ : CascadeMux
    port map (
            O => \N__12776\,
            I => \N__12773\
        );

    \I__2201\ : InMux
    port map (
            O => \N__12773\,
            I => \N__12769\
        );

    \I__2200\ : InMux
    port map (
            O => \N__12772\,
            I => \N__12766\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__12769\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__12766\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__2197\ : CascadeMux
    port map (
            O => \N__12761\,
            I => \N__12758\
        );

    \I__2196\ : InMux
    port map (
            O => \N__12758\,
            I => \N__12755\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__12755\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_6\
        );

    \I__2194\ : InMux
    port map (
            O => \N__12752\,
            I => \N__12748\
        );

    \I__2193\ : InMux
    port map (
            O => \N__12751\,
            I => \N__12745\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__12748\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__12745\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__2190\ : CascadeMux
    port map (
            O => \N__12740\,
            I => \N__12737\
        );

    \I__2189\ : InMux
    port map (
            O => \N__12737\,
            I => \N__12734\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__12734\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_7\
        );

    \I__2187\ : InMux
    port map (
            O => \N__12731\,
            I => \N__12728\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__12728\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__2185\ : InMux
    port map (
            O => \N__12725\,
            I => \N__12722\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__12722\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg_5_0_o2_0_7_9\
        );

    \I__2183\ : CascadeMux
    port map (
            O => \N__12719\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg_5_0_o2_0_6_9_cascade_\
        );

    \I__2182\ : InMux
    port map (
            O => \N__12716\,
            I => \N__12713\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__12713\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_30\
        );

    \I__2180\ : InMux
    port map (
            O => \N__12710\,
            I => \N__12707\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__12707\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__2178\ : InMux
    port map (
            O => \N__12704\,
            I => \N__12701\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__12701\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg_5_0_o2_0_0_9\
        );

    \I__2176\ : CascadeMux
    port map (
            O => \N__12698\,
            I => \N__12693\
        );

    \I__2175\ : InMux
    port map (
            O => \N__12697\,
            I => \N__12690\
        );

    \I__2174\ : InMux
    port map (
            O => \N__12696\,
            I => \N__12687\
        );

    \I__2173\ : InMux
    port map (
            O => \N__12693\,
            I => \N__12684\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__12690\,
            I => \N__12679\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__12687\,
            I => \N__12679\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__12684\,
            I => \N__12676\
        );

    \I__2169\ : Odrv4
    port map (
            O => \N__12679\,
            I => \delay_measurement_inst.elapsed_time_hc_19\
        );

    \I__2168\ : Odrv4
    port map (
            O => \N__12676\,
            I => \delay_measurement_inst.elapsed_time_hc_19\
        );

    \I__2167\ : CascadeMux
    port map (
            O => \N__12671\,
            I => \N__12668\
        );

    \I__2166\ : InMux
    port map (
            O => \N__12668\,
            I => \N__12663\
        );

    \I__2165\ : InMux
    port map (
            O => \N__12667\,
            I => \N__12660\
        );

    \I__2164\ : InMux
    port map (
            O => \N__12666\,
            I => \N__12657\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__12663\,
            I => \N__12654\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__12660\,
            I => \N__12651\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__12657\,
            I => \delay_measurement_inst.elapsed_time_hc_16\
        );

    \I__2160\ : Odrv4
    port map (
            O => \N__12654\,
            I => \delay_measurement_inst.elapsed_time_hc_16\
        );

    \I__2159\ : Odrv4
    port map (
            O => \N__12651\,
            I => \delay_measurement_inst.elapsed_time_hc_16\
        );

    \I__2158\ : InMux
    port map (
            O => \N__12644\,
            I => \N__12640\
        );

    \I__2157\ : InMux
    port map (
            O => \N__12643\,
            I => \N__12637\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__12640\,
            I => \delay_measurement_inst.elapsed_time_hc_3\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__12637\,
            I => \delay_measurement_inst.elapsed_time_hc_3\
        );

    \I__2154\ : InMux
    port map (
            O => \N__12632\,
            I => \N__12627\
        );

    \I__2153\ : InMux
    port map (
            O => \N__12631\,
            I => \N__12624\
        );

    \I__2152\ : InMux
    port map (
            O => \N__12630\,
            I => \N__12620\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__12627\,
            I => \N__12615\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__12624\,
            I => \N__12615\
        );

    \I__2149\ : InMux
    port map (
            O => \N__12623\,
            I => \N__12612\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__12620\,
            I => \N__12608\
        );

    \I__2147\ : Span4Mux_v
    port map (
            O => \N__12615\,
            I => \N__12603\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__12612\,
            I => \N__12603\
        );

    \I__2145\ : InMux
    port map (
            O => \N__12611\,
            I => \N__12600\
        );

    \I__2144\ : Span12Mux_v
    port map (
            O => \N__12608\,
            I => \N__12597\
        );

    \I__2143\ : Span4Mux_v
    port map (
            O => \N__12603\,
            I => \N__12594\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__12600\,
            I => measured_delay_tr_8
        );

    \I__2141\ : Odrv12
    port map (
            O => \N__12597\,
            I => measured_delay_tr_8
        );

    \I__2140\ : Odrv4
    port map (
            O => \N__12594\,
            I => measured_delay_tr_8
        );

    \I__2139\ : InMux
    port map (
            O => \N__12587\,
            I => \N__12584\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__12584\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__2137\ : InMux
    port map (
            O => \N__12581\,
            I => \N__12578\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__12578\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__2135\ : CascadeMux
    port map (
            O => \N__12575\,
            I => \N__12572\
        );

    \I__2134\ : InMux
    port map (
            O => \N__12572\,
            I => \N__12569\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__12569\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__2132\ : InMux
    port map (
            O => \N__12566\,
            I => \N__12563\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__12563\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__2130\ : InMux
    port map (
            O => \N__12560\,
            I => \N__12557\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__12557\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__2128\ : InMux
    port map (
            O => \N__12554\,
            I => \N__12551\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__12551\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__2126\ : CascadeMux
    port map (
            O => \N__12548\,
            I => \N__12545\
        );

    \I__2125\ : InMux
    port map (
            O => \N__12545\,
            I => \N__12542\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__12542\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__2123\ : InMux
    port map (
            O => \N__12539\,
            I => \N__12536\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__12536\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__2121\ : InMux
    port map (
            O => \N__12533\,
            I => \N__12530\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__12530\,
            I => \delay_measurement_inst.delay_hc_timer.N_101\
        );

    \I__2119\ : CascadeMux
    port map (
            O => \N__12527\,
            I => \delay_measurement_inst.delay_hc_timer.N_81_cascade_\
        );

    \I__2118\ : InMux
    port map (
            O => \N__12524\,
            I => \N__12521\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__12521\,
            I => \delay_measurement_inst.delay_hc_timer.un1_reset_1_i_a2_4\
        );

    \I__2116\ : CascadeMux
    port map (
            O => \N__12518\,
            I => \delay_measurement_inst.delay_hc_timer.un1_reset_1_i_a2_6_cascade_\
        );

    \I__2115\ : InMux
    port map (
            O => \N__12515\,
            I => \N__12512\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__12512\,
            I => \delay_measurement_inst.delay_hc_timer.un1_reset_1_i_a2_5\
        );

    \I__2113\ : InMux
    port map (
            O => \N__12509\,
            I => \N__12503\
        );

    \I__2112\ : InMux
    port map (
            O => \N__12508\,
            I => \N__12503\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__12503\,
            I => \delay_measurement_inst.delay_hc_timer.N_105\
        );

    \I__2110\ : InMux
    port map (
            O => \N__12500\,
            I => \N__12497\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__12497\,
            I => \delay_measurement_inst.delay_hc_timer.un1_reset_1_i_0\
        );

    \I__2108\ : CascadeMux
    port map (
            O => \N__12494\,
            I => \delay_measurement_inst.delay_hc_timer.un1_reset_1_i_a2_9_cascade_\
        );

    \I__2107\ : InMux
    port map (
            O => \N__12491\,
            I => \N__12488\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__12488\,
            I => \N__12484\
        );

    \I__2105\ : InMux
    port map (
            O => \N__12487\,
            I => \N__12481\
        );

    \I__2104\ : Span4Mux_v
    port map (
            O => \N__12484\,
            I => \N__12476\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__12481\,
            I => \N__12476\
        );

    \I__2102\ : Odrv4
    port map (
            O => \N__12476\,
            I => \delay_measurement_inst.elapsed_time_hc_2\
        );

    \I__2101\ : InMux
    port map (
            O => \N__12473\,
            I => \N__12469\
        );

    \I__2100\ : InMux
    port map (
            O => \N__12472\,
            I => \N__12466\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__12469\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__12466\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__2097\ : InMux
    port map (
            O => \N__12461\,
            I => \N__12458\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__12458\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\
        );

    \I__2095\ : InMux
    port map (
            O => \N__12455\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\
        );

    \I__2094\ : InMux
    port map (
            O => \N__12452\,
            I => \N__12448\
        );

    \I__2093\ : InMux
    port map (
            O => \N__12451\,
            I => \N__12445\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__12448\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__12445\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__2090\ : InMux
    port map (
            O => \N__12440\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\
        );

    \I__2089\ : InMux
    port map (
            O => \N__12437\,
            I => \N__12434\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__12434\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\
        );

    \I__2087\ : IoInMux
    port map (
            O => \N__12431\,
            I => \N__12428\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__12428\,
            I => \N__12425\
        );

    \I__2085\ : Span4Mux_s3_v
    port map (
            O => \N__12425\,
            I => \N__12422\
        );

    \I__2084\ : Sp12to4
    port map (
            O => \N__12422\,
            I => \N__12419\
        );

    \I__2083\ : Span12Mux_s9_h
    port map (
            O => \N__12419\,
            I => \N__12416\
        );

    \I__2082\ : Span12Mux_v
    port map (
            O => \N__12416\,
            I => \N__12413\
        );

    \I__2081\ : Odrv12
    port map (
            O => \N__12413\,
            I => \delay_measurement_inst.delay_tr_timer.N_180_i\
        );

    \I__2080\ : InMux
    port map (
            O => \N__12410\,
            I => \N__12407\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__12407\,
            I => \N__12404\
        );

    \I__2078\ : Odrv12
    port map (
            O => \N__12404\,
            I => il_min_comp1_c
        );

    \I__2077\ : InMux
    port map (
            O => \N__12401\,
            I => \N__12398\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__12398\,
            I => \N__12394\
        );

    \I__2075\ : InMux
    port map (
            O => \N__12397\,
            I => \N__12391\
        );

    \I__2074\ : Odrv4
    port map (
            O => \N__12394\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__12391\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__2072\ : CascadeMux
    port map (
            O => \N__12386\,
            I => \N__12383\
        );

    \I__2071\ : InMux
    port map (
            O => \N__12383\,
            I => \N__12380\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__12380\,
            I => \N__12377\
        );

    \I__2069\ : Odrv4
    port map (
            O => \N__12377\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\
        );

    \I__2068\ : InMux
    port map (
            O => \N__12374\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\
        );

    \I__2067\ : InMux
    port map (
            O => \N__12371\,
            I => \N__12367\
        );

    \I__2066\ : InMux
    port map (
            O => \N__12370\,
            I => \N__12364\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__12367\,
            I => \N__12361\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__12364\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__2063\ : Odrv4
    port map (
            O => \N__12361\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__2062\ : InMux
    port map (
            O => \N__12356\,
            I => \N__12353\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__12353\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\
        );

    \I__2060\ : InMux
    port map (
            O => \N__12350\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\
        );

    \I__2059\ : InMux
    port map (
            O => \N__12347\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\
        );

    \I__2058\ : InMux
    port map (
            O => \N__12344\,
            I => \N__12340\
        );

    \I__2057\ : InMux
    port map (
            O => \N__12343\,
            I => \N__12337\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__12340\,
            I => \N__12334\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__12337\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__2054\ : Odrv4
    port map (
            O => \N__12334\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__2053\ : InMux
    port map (
            O => \N__12329\,
            I => \N__12326\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__12326\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\
        );

    \I__2051\ : InMux
    port map (
            O => \N__12323\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__12320\,
            I => \N__12316\
        );

    \I__2049\ : InMux
    port map (
            O => \N__12319\,
            I => \N__12313\
        );

    \I__2048\ : InMux
    port map (
            O => \N__12316\,
            I => \N__12310\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__12313\,
            I => \N__12307\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__12310\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__2045\ : Odrv4
    port map (
            O => \N__12307\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__2044\ : CascadeMux
    port map (
            O => \N__12302\,
            I => \N__12299\
        );

    \I__2043\ : InMux
    port map (
            O => \N__12299\,
            I => \N__12296\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__12296\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\
        );

    \I__2041\ : InMux
    port map (
            O => \N__12293\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\
        );

    \I__2040\ : InMux
    port map (
            O => \N__12290\,
            I => \N__12286\
        );

    \I__2039\ : InMux
    port map (
            O => \N__12289\,
            I => \N__12283\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__12286\,
            I => \N__12280\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__12283\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__2036\ : Odrv4
    port map (
            O => \N__12280\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__2035\ : InMux
    port map (
            O => \N__12275\,
            I => \N__12272\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__12272\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\
        );

    \I__2033\ : InMux
    port map (
            O => \N__12269\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\
        );

    \I__2032\ : InMux
    port map (
            O => \N__12266\,
            I => \N__12262\
        );

    \I__2031\ : InMux
    port map (
            O => \N__12265\,
            I => \N__12259\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__12262\,
            I => \N__12256\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__12259\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__2028\ : Odrv4
    port map (
            O => \N__12256\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__2027\ : CascadeMux
    port map (
            O => \N__12251\,
            I => \N__12248\
        );

    \I__2026\ : InMux
    port map (
            O => \N__12248\,
            I => \N__12245\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__12245\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\
        );

    \I__2024\ : InMux
    port map (
            O => \N__12242\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\
        );

    \I__2023\ : InMux
    port map (
            O => \N__12239\,
            I => \N__12235\
        );

    \I__2022\ : InMux
    port map (
            O => \N__12238\,
            I => \N__12232\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__12235\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__12232\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__2019\ : InMux
    port map (
            O => \N__12227\,
            I => \N__12224\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__12224\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\
        );

    \I__2017\ : InMux
    port map (
            O => \N__12221\,
            I => \bfn_8_27_0_\
        );

    \I__2016\ : InMux
    port map (
            O => \N__12218\,
            I => \N__12215\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__12215\,
            I => \N__12212\
        );

    \I__2014\ : Odrv4
    port map (
            O => \N__12212\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\
        );

    \I__2013\ : InMux
    port map (
            O => \N__12209\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\
        );

    \I__2012\ : InMux
    port map (
            O => \N__12206\,
            I => \N__12202\
        );

    \I__2011\ : InMux
    port map (
            O => \N__12205\,
            I => \N__12199\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__12202\,
            I => \N__12196\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__12199\,
            I => \N__12193\
        );

    \I__2008\ : Odrv4
    port map (
            O => \N__12196\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__2007\ : Odrv4
    port map (
            O => \N__12193\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__2006\ : CascadeMux
    port map (
            O => \N__12188\,
            I => \N__12185\
        );

    \I__2005\ : InMux
    port map (
            O => \N__12185\,
            I => \N__12182\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__12182\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNI62NAZ0\
        );

    \I__2003\ : InMux
    port map (
            O => \N__12179\,
            I => \N__12176\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__12176\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\
        );

    \I__2001\ : InMux
    port map (
            O => \N__12173\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\
        );

    \I__2000\ : InMux
    port map (
            O => \N__12170\,
            I => \N__12166\
        );

    \I__1999\ : InMux
    port map (
            O => \N__12169\,
            I => \N__12163\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__12166\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__12163\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__1996\ : InMux
    port map (
            O => \N__12158\,
            I => \N__12155\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__12155\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\
        );

    \I__1994\ : InMux
    port map (
            O => \N__12152\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\
        );

    \I__1993\ : InMux
    port map (
            O => \N__12149\,
            I => \N__12145\
        );

    \I__1992\ : InMux
    port map (
            O => \N__12148\,
            I => \N__12142\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__12145\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__12142\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__1989\ : InMux
    port map (
            O => \N__12137\,
            I => \N__12134\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__12134\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\
        );

    \I__1987\ : InMux
    port map (
            O => \N__12131\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\
        );

    \I__1986\ : InMux
    port map (
            O => \N__12128\,
            I => \N__12124\
        );

    \I__1985\ : InMux
    port map (
            O => \N__12127\,
            I => \N__12121\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__12124\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__12121\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__1982\ : InMux
    port map (
            O => \N__12116\,
            I => \N__12113\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__12113\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\
        );

    \I__1980\ : InMux
    port map (
            O => \N__12110\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\
        );

    \I__1979\ : InMux
    port map (
            O => \N__12107\,
            I => \N__12103\
        );

    \I__1978\ : InMux
    port map (
            O => \N__12106\,
            I => \N__12100\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__12103\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__12100\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__1975\ : InMux
    port map (
            O => \N__12095\,
            I => \N__12092\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__12092\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\
        );

    \I__1973\ : InMux
    port map (
            O => \N__12089\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\
        );

    \I__1972\ : InMux
    port map (
            O => \N__12086\,
            I => \N__12083\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__12083\,
            I => \N__12079\
        );

    \I__1970\ : InMux
    port map (
            O => \N__12082\,
            I => \N__12076\
        );

    \I__1969\ : Odrv4
    port map (
            O => \N__12079\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__12076\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__1967\ : InMux
    port map (
            O => \N__12071\,
            I => \N__12068\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__12068\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\
        );

    \I__1965\ : InMux
    port map (
            O => \N__12065\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\
        );

    \I__1964\ : InMux
    port map (
            O => \N__12062\,
            I => \N__12059\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__12059\,
            I => \N__12055\
        );

    \I__1962\ : InMux
    port map (
            O => \N__12058\,
            I => \N__12052\
        );

    \I__1961\ : Odrv4
    port map (
            O => \N__12055\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__12052\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__1959\ : InMux
    port map (
            O => \N__12047\,
            I => \N__12044\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__12044\,
            I => \N__12041\
        );

    \I__1957\ : Odrv4
    port map (
            O => \N__12041\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\
        );

    \I__1956\ : InMux
    port map (
            O => \N__12038\,
            I => \bfn_8_26_0_\
        );

    \I__1955\ : CEMux
    port map (
            O => \N__12035\,
            I => \N__12032\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__12032\,
            I => \N__12026\
        );

    \I__1953\ : CEMux
    port map (
            O => \N__12031\,
            I => \N__12023\
        );

    \I__1952\ : CEMux
    port map (
            O => \N__12030\,
            I => \N__12020\
        );

    \I__1951\ : CEMux
    port map (
            O => \N__12029\,
            I => \N__12017\
        );

    \I__1950\ : Span4Mux_v
    port map (
            O => \N__12026\,
            I => \N__12011\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__12023\,
            I => \N__12011\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__12020\,
            I => \N__12008\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__12017\,
            I => \N__12005\
        );

    \I__1946\ : CEMux
    port map (
            O => \N__12016\,
            I => \N__12002\
        );

    \I__1945\ : Span4Mux_h
    port map (
            O => \N__12011\,
            I => \N__11999\
        );

    \I__1944\ : Span4Mux_v
    port map (
            O => \N__12008\,
            I => \N__11994\
        );

    \I__1943\ : Span4Mux_h
    port map (
            O => \N__12005\,
            I => \N__11994\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__12002\,
            I => \N__11991\
        );

    \I__1941\ : Odrv4
    port map (
            O => \N__11999\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJMZ0Z_1\
        );

    \I__1940\ : Odrv4
    port map (
            O => \N__11994\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJMZ0Z_1\
        );

    \I__1939\ : Odrv12
    port map (
            O => \N__11991\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJMZ0Z_1\
        );

    \I__1938\ : CascadeMux
    port map (
            O => \N__11984\,
            I => \N__11981\
        );

    \I__1937\ : InMux
    port map (
            O => \N__11981\,
            I => \N__11977\
        );

    \I__1936\ : InMux
    port map (
            O => \N__11980\,
            I => \N__11974\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__11977\,
            I => \N__11968\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__11974\,
            I => \N__11968\
        );

    \I__1933\ : InMux
    port map (
            O => \N__11973\,
            I => \N__11965\
        );

    \I__1932\ : Odrv4
    port map (
            O => \N__11968\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__11965\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__1930\ : CascadeMux
    port map (
            O => \N__11960\,
            I => \N__11957\
        );

    \I__1929\ : InMux
    port map (
            O => \N__11957\,
            I => \N__11954\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__11954\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\
        );

    \I__1927\ : InMux
    port map (
            O => \N__11951\,
            I => \N__11948\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__11948\,
            I => \N__11944\
        );

    \I__1925\ : InMux
    port map (
            O => \N__11947\,
            I => \N__11941\
        );

    \I__1924\ : Odrv4
    port map (
            O => \N__11944\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__11941\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__1922\ : InMux
    port map (
            O => \N__11936\,
            I => \N__11933\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__11933\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\
        );

    \I__1920\ : InMux
    port map (
            O => \N__11930\,
            I => \N__11927\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__11927\,
            I => \N__11924\
        );

    \I__1918\ : Span4Mux_h
    port map (
            O => \N__11924\,
            I => \N__11921\
        );

    \I__1917\ : Odrv4
    port map (
            O => \N__11921\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\
        );

    \I__1916\ : InMux
    port map (
            O => \N__11918\,
            I => \N__11915\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__11915\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\
        );

    \I__1914\ : InMux
    port map (
            O => \N__11912\,
            I => \N__11909\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__11909\,
            I => \N__11906\
        );

    \I__1912\ : Sp12to4
    port map (
            O => \N__11906\,
            I => \N__11903\
        );

    \I__1911\ : Odrv12
    port map (
            O => \N__11903\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\
        );

    \I__1910\ : CascadeMux
    port map (
            O => \N__11900\,
            I => \N__11894\
        );

    \I__1909\ : InMux
    port map (
            O => \N__11899\,
            I => \N__11883\
        );

    \I__1908\ : InMux
    port map (
            O => \N__11898\,
            I => \N__11883\
        );

    \I__1907\ : InMux
    port map (
            O => \N__11897\,
            I => \N__11883\
        );

    \I__1906\ : InMux
    port map (
            O => \N__11894\,
            I => \N__11878\
        );

    \I__1905\ : InMux
    port map (
            O => \N__11893\,
            I => \N__11878\
        );

    \I__1904\ : CascadeMux
    port map (
            O => \N__11892\,
            I => \N__11869\
        );

    \I__1903\ : InMux
    port map (
            O => \N__11891\,
            I => \N__11864\
        );

    \I__1902\ : InMux
    port map (
            O => \N__11890\,
            I => \N__11864\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__11883\,
            I => \N__11861\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__11878\,
            I => \N__11858\
        );

    \I__1899\ : InMux
    port map (
            O => \N__11877\,
            I => \N__11847\
        );

    \I__1898\ : InMux
    port map (
            O => \N__11876\,
            I => \N__11847\
        );

    \I__1897\ : InMux
    port map (
            O => \N__11875\,
            I => \N__11847\
        );

    \I__1896\ : InMux
    port map (
            O => \N__11874\,
            I => \N__11847\
        );

    \I__1895\ : InMux
    port map (
            O => \N__11873\,
            I => \N__11847\
        );

    \I__1894\ : CascadeMux
    port map (
            O => \N__11872\,
            I => \N__11844\
        );

    \I__1893\ : InMux
    port map (
            O => \N__11869\,
            I => \N__11835\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__11864\,
            I => \N__11832\
        );

    \I__1891\ : Span4Mux_v
    port map (
            O => \N__11861\,
            I => \N__11825\
        );

    \I__1890\ : Span4Mux_v
    port map (
            O => \N__11858\,
            I => \N__11825\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__11847\,
            I => \N__11825\
        );

    \I__1888\ : InMux
    port map (
            O => \N__11844\,
            I => \N__11818\
        );

    \I__1887\ : InMux
    port map (
            O => \N__11843\,
            I => \N__11818\
        );

    \I__1886\ : InMux
    port map (
            O => \N__11842\,
            I => \N__11818\
        );

    \I__1885\ : InMux
    port map (
            O => \N__11841\,
            I => \N__11811\
        );

    \I__1884\ : InMux
    port map (
            O => \N__11840\,
            I => \N__11811\
        );

    \I__1883\ : InMux
    port map (
            O => \N__11839\,
            I => \N__11811\
        );

    \I__1882\ : InMux
    port map (
            O => \N__11838\,
            I => \N__11808\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__11835\,
            I => \N__11803\
        );

    \I__1880\ : Span4Mux_h
    port map (
            O => \N__11832\,
            I => \N__11803\
        );

    \I__1879\ : Span4Mux_h
    port map (
            O => \N__11825\,
            I => \N__11800\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__11818\,
            I => \phase_controller_inst1.stoper_tr.un3_start\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__11811\,
            I => \phase_controller_inst1.stoper_tr.un3_start\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__11808\,
            I => \phase_controller_inst1.stoper_tr.un3_start\
        );

    \I__1875\ : Odrv4
    port map (
            O => \N__11803\,
            I => \phase_controller_inst1.stoper_tr.un3_start\
        );

    \I__1874\ : Odrv4
    port map (
            O => \N__11800\,
            I => \phase_controller_inst1.stoper_tr.un3_start\
        );

    \I__1873\ : CascadeMux
    port map (
            O => \N__11789\,
            I => \N__11778\
        );

    \I__1872\ : CascadeMux
    port map (
            O => \N__11788\,
            I => \N__11774\
        );

    \I__1871\ : CascadeMux
    port map (
            O => \N__11787\,
            I => \N__11771\
        );

    \I__1870\ : CascadeMux
    port map (
            O => \N__11786\,
            I => \N__11767\
        );

    \I__1869\ : CascadeMux
    port map (
            O => \N__11785\,
            I => \N__11764\
        );

    \I__1868\ : CascadeMux
    port map (
            O => \N__11784\,
            I => \N__11758\
        );

    \I__1867\ : CascadeMux
    port map (
            O => \N__11783\,
            I => \N__11755\
        );

    \I__1866\ : CascadeMux
    port map (
            O => \N__11782\,
            I => \N__11752\
        );

    \I__1865\ : InMux
    port map (
            O => \N__11781\,
            I => \N__11742\
        );

    \I__1864\ : InMux
    port map (
            O => \N__11778\,
            I => \N__11735\
        );

    \I__1863\ : InMux
    port map (
            O => \N__11777\,
            I => \N__11735\
        );

    \I__1862\ : InMux
    port map (
            O => \N__11774\,
            I => \N__11735\
        );

    \I__1861\ : InMux
    port map (
            O => \N__11771\,
            I => \N__11724\
        );

    \I__1860\ : InMux
    port map (
            O => \N__11770\,
            I => \N__11724\
        );

    \I__1859\ : InMux
    port map (
            O => \N__11767\,
            I => \N__11724\
        );

    \I__1858\ : InMux
    port map (
            O => \N__11764\,
            I => \N__11724\
        );

    \I__1857\ : InMux
    port map (
            O => \N__11763\,
            I => \N__11724\
        );

    \I__1856\ : InMux
    port map (
            O => \N__11762\,
            I => \N__11717\
        );

    \I__1855\ : InMux
    port map (
            O => \N__11761\,
            I => \N__11717\
        );

    \I__1854\ : InMux
    port map (
            O => \N__11758\,
            I => \N__11717\
        );

    \I__1853\ : InMux
    port map (
            O => \N__11755\,
            I => \N__11708\
        );

    \I__1852\ : InMux
    port map (
            O => \N__11752\,
            I => \N__11708\
        );

    \I__1851\ : InMux
    port map (
            O => \N__11751\,
            I => \N__11708\
        );

    \I__1850\ : InMux
    port map (
            O => \N__11750\,
            I => \N__11708\
        );

    \I__1849\ : CascadeMux
    port map (
            O => \N__11749\,
            I => \N__11703\
        );

    \I__1848\ : CascadeMux
    port map (
            O => \N__11748\,
            I => \N__11698\
        );

    \I__1847\ : CascadeMux
    port map (
            O => \N__11747\,
            I => \N__11695\
        );

    \I__1846\ : CascadeMux
    port map (
            O => \N__11746\,
            I => \N__11692\
        );

    \I__1845\ : CascadeMux
    port map (
            O => \N__11745\,
            I => \N__11689\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__11742\,
            I => \N__11686\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__11735\,
            I => \N__11683\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__11724\,
            I => \N__11676\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__11717\,
            I => \N__11676\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__11708\,
            I => \N__11676\
        );

    \I__1839\ : InMux
    port map (
            O => \N__11707\,
            I => \N__11670\
        );

    \I__1838\ : InMux
    port map (
            O => \N__11706\,
            I => \N__11667\
        );

    \I__1837\ : InMux
    port map (
            O => \N__11703\,
            I => \N__11658\
        );

    \I__1836\ : InMux
    port map (
            O => \N__11702\,
            I => \N__11658\
        );

    \I__1835\ : InMux
    port map (
            O => \N__11701\,
            I => \N__11658\
        );

    \I__1834\ : InMux
    port map (
            O => \N__11698\,
            I => \N__11658\
        );

    \I__1833\ : InMux
    port map (
            O => \N__11695\,
            I => \N__11651\
        );

    \I__1832\ : InMux
    port map (
            O => \N__11692\,
            I => \N__11651\
        );

    \I__1831\ : InMux
    port map (
            O => \N__11689\,
            I => \N__11651\
        );

    \I__1830\ : Span4Mux_v
    port map (
            O => \N__11686\,
            I => \N__11644\
        );

    \I__1829\ : Span4Mux_v
    port map (
            O => \N__11683\,
            I => \N__11644\
        );

    \I__1828\ : Span4Mux_v
    port map (
            O => \N__11676\,
            I => \N__11644\
        );

    \I__1827\ : InMux
    port map (
            O => \N__11675\,
            I => \N__11639\
        );

    \I__1826\ : InMux
    port map (
            O => \N__11674\,
            I => \N__11639\
        );

    \I__1825\ : InMux
    port map (
            O => \N__11673\,
            I => \N__11636\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__11670\,
            I => \N__11633\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__11667\,
            I => \phase_controller_inst1.stoper_tr.un1_startlto19Z0Z_2\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__11658\,
            I => \phase_controller_inst1.stoper_tr.un1_startlto19Z0Z_2\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__11651\,
            I => \phase_controller_inst1.stoper_tr.un1_startlto19Z0Z_2\
        );

    \I__1820\ : Odrv4
    port map (
            O => \N__11644\,
            I => \phase_controller_inst1.stoper_tr.un1_startlto19Z0Z_2\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__11639\,
            I => \phase_controller_inst1.stoper_tr.un1_startlto19Z0Z_2\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__11636\,
            I => \phase_controller_inst1.stoper_tr.un1_startlto19Z0Z_2\
        );

    \I__1817\ : Odrv4
    port map (
            O => \N__11633\,
            I => \phase_controller_inst1.stoper_tr.un1_startlto19Z0Z_2\
        );

    \I__1816\ : InMux
    port map (
            O => \N__11618\,
            I => \N__11602\
        );

    \I__1815\ : InMux
    port map (
            O => \N__11617\,
            I => \N__11602\
        );

    \I__1814\ : InMux
    port map (
            O => \N__11616\,
            I => \N__11602\
        );

    \I__1813\ : InMux
    port map (
            O => \N__11615\,
            I => \N__11591\
        );

    \I__1812\ : InMux
    port map (
            O => \N__11614\,
            I => \N__11591\
        );

    \I__1811\ : InMux
    port map (
            O => \N__11613\,
            I => \N__11591\
        );

    \I__1810\ : InMux
    port map (
            O => \N__11612\,
            I => \N__11591\
        );

    \I__1809\ : InMux
    port map (
            O => \N__11611\,
            I => \N__11591\
        );

    \I__1808\ : InMux
    port map (
            O => \N__11610\,
            I => \N__11586\
        );

    \I__1807\ : InMux
    port map (
            O => \N__11609\,
            I => \N__11586\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__11602\,
            I => \N__11572\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__11591\,
            I => \N__11567\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__11586\,
            I => \N__11567\
        );

    \I__1803\ : InMux
    port map (
            O => \N__11585\,
            I => \N__11560\
        );

    \I__1802\ : InMux
    port map (
            O => \N__11584\,
            I => \N__11560\
        );

    \I__1801\ : InMux
    port map (
            O => \N__11583\,
            I => \N__11560\
        );

    \I__1800\ : InMux
    port map (
            O => \N__11582\,
            I => \N__11551\
        );

    \I__1799\ : InMux
    port map (
            O => \N__11581\,
            I => \N__11551\
        );

    \I__1798\ : InMux
    port map (
            O => \N__11580\,
            I => \N__11551\
        );

    \I__1797\ : InMux
    port map (
            O => \N__11579\,
            I => \N__11551\
        );

    \I__1796\ : InMux
    port map (
            O => \N__11578\,
            I => \N__11542\
        );

    \I__1795\ : InMux
    port map (
            O => \N__11577\,
            I => \N__11542\
        );

    \I__1794\ : InMux
    port map (
            O => \N__11576\,
            I => \N__11542\
        );

    \I__1793\ : InMux
    port map (
            O => \N__11575\,
            I => \N__11542\
        );

    \I__1792\ : Span4Mux_v
    port map (
            O => \N__11572\,
            I => \N__11535\
        );

    \I__1791\ : Span4Mux_v
    port map (
            O => \N__11567\,
            I => \N__11535\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__11560\,
            I => \N__11532\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__11551\,
            I => \N__11529\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__11542\,
            I => \N__11526\
        );

    \I__1787\ : InMux
    port map (
            O => \N__11541\,
            I => \N__11523\
        );

    \I__1786\ : InMux
    port map (
            O => \N__11540\,
            I => \N__11520\
        );

    \I__1785\ : Odrv4
    port map (
            O => \N__11535\,
            I => \phase_controller_inst1.stoper_tr.un1_startlt15\
        );

    \I__1784\ : Odrv4
    port map (
            O => \N__11532\,
            I => \phase_controller_inst1.stoper_tr.un1_startlt15\
        );

    \I__1783\ : Odrv12
    port map (
            O => \N__11529\,
            I => \phase_controller_inst1.stoper_tr.un1_startlt15\
        );

    \I__1782\ : Odrv4
    port map (
            O => \N__11526\,
            I => \phase_controller_inst1.stoper_tr.un1_startlt15\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__11523\,
            I => \phase_controller_inst1.stoper_tr.un1_startlt15\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__11520\,
            I => \phase_controller_inst1.stoper_tr.un1_startlt15\
        );

    \I__1779\ : InMux
    port map (
            O => \N__11507\,
            I => \N__11504\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__11504\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\
        );

    \I__1777\ : CascadeMux
    port map (
            O => \N__11501\,
            I => \N__11498\
        );

    \I__1776\ : InMux
    port map (
            O => \N__11498\,
            I => \N__11495\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__11495\,
            I => \N__11492\
        );

    \I__1774\ : Odrv4
    port map (
            O => \N__11492\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0\
        );

    \I__1773\ : InMux
    port map (
            O => \N__11489\,
            I => \N__11486\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__11486\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18\
        );

    \I__1771\ : InMux
    port map (
            O => \N__11483\,
            I => \N__11480\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__11480\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19\
        );

    \I__1769\ : InMux
    port map (
            O => \N__11477\,
            I => \N__11441\
        );

    \I__1768\ : InMux
    port map (
            O => \N__11476\,
            I => \N__11441\
        );

    \I__1767\ : InMux
    port map (
            O => \N__11475\,
            I => \N__11441\
        );

    \I__1766\ : InMux
    port map (
            O => \N__11474\,
            I => \N__11441\
        );

    \I__1765\ : InMux
    port map (
            O => \N__11473\,
            I => \N__11441\
        );

    \I__1764\ : InMux
    port map (
            O => \N__11472\,
            I => \N__11441\
        );

    \I__1763\ : InMux
    port map (
            O => \N__11471\,
            I => \N__11441\
        );

    \I__1762\ : InMux
    port map (
            O => \N__11470\,
            I => \N__11441\
        );

    \I__1761\ : InMux
    port map (
            O => \N__11469\,
            I => \N__11430\
        );

    \I__1760\ : InMux
    port map (
            O => \N__11468\,
            I => \N__11430\
        );

    \I__1759\ : InMux
    port map (
            O => \N__11467\,
            I => \N__11430\
        );

    \I__1758\ : InMux
    port map (
            O => \N__11466\,
            I => \N__11430\
        );

    \I__1757\ : InMux
    port map (
            O => \N__11465\,
            I => \N__11430\
        );

    \I__1756\ : InMux
    port map (
            O => \N__11464\,
            I => \N__11411\
        );

    \I__1755\ : InMux
    port map (
            O => \N__11463\,
            I => \N__11411\
        );

    \I__1754\ : InMux
    port map (
            O => \N__11462\,
            I => \N__11411\
        );

    \I__1753\ : InMux
    port map (
            O => \N__11461\,
            I => \N__11411\
        );

    \I__1752\ : InMux
    port map (
            O => \N__11460\,
            I => \N__11411\
        );

    \I__1751\ : InMux
    port map (
            O => \N__11459\,
            I => \N__11411\
        );

    \I__1750\ : InMux
    port map (
            O => \N__11458\,
            I => \N__11411\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__11441\,
            I => \N__11406\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__11430\,
            I => \N__11406\
        );

    \I__1747\ : InMux
    port map (
            O => \N__11429\,
            I => \N__11403\
        );

    \I__1746\ : InMux
    port map (
            O => \N__11428\,
            I => \N__11400\
        );

    \I__1745\ : InMux
    port map (
            O => \N__11427\,
            I => \N__11397\
        );

    \I__1744\ : InMux
    port map (
            O => \N__11426\,
            I => \N__11394\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__11411\,
            I => \N__11387\
        );

    \I__1742\ : Span4Mux_v
    port map (
            O => \N__11406\,
            I => \N__11387\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__11403\,
            I => \N__11387\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__11400\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__11397\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__11394\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__1737\ : Odrv4
    port map (
            O => \N__11387\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__1736\ : CascadeMux
    port map (
            O => \N__11378\,
            I => \N__11375\
        );

    \I__1735\ : InMux
    port map (
            O => \N__11375\,
            I => \N__11372\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__11372\,
            I => \N__11369\
        );

    \I__1733\ : Odrv4
    port map (
            O => \N__11369\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2\
        );

    \I__1732\ : CascadeMux
    port map (
            O => \N__11366\,
            I => \N__11353\
        );

    \I__1731\ : CascadeMux
    port map (
            O => \N__11365\,
            I => \N__11347\
        );

    \I__1730\ : CascadeMux
    port map (
            O => \N__11364\,
            I => \N__11344\
        );

    \I__1729\ : CascadeMux
    port map (
            O => \N__11363\,
            I => \N__11341\
        );

    \I__1728\ : CascadeMux
    port map (
            O => \N__11362\,
            I => \N__11338\
        );

    \I__1727\ : CascadeMux
    port map (
            O => \N__11361\,
            I => \N__11334\
        );

    \I__1726\ : InMux
    port map (
            O => \N__11360\,
            I => \N__11326\
        );

    \I__1725\ : InMux
    port map (
            O => \N__11359\,
            I => \N__11326\
        );

    \I__1724\ : CascadeMux
    port map (
            O => \N__11358\,
            I => \N__11319\
        );

    \I__1723\ : CascadeMux
    port map (
            O => \N__11357\,
            I => \N__11316\
        );

    \I__1722\ : CascadeMux
    port map (
            O => \N__11356\,
            I => \N__11313\
        );

    \I__1721\ : InMux
    port map (
            O => \N__11353\,
            I => \N__11309\
        );

    \I__1720\ : InMux
    port map (
            O => \N__11352\,
            I => \N__11294\
        );

    \I__1719\ : InMux
    port map (
            O => \N__11351\,
            I => \N__11294\
        );

    \I__1718\ : InMux
    port map (
            O => \N__11350\,
            I => \N__11294\
        );

    \I__1717\ : InMux
    port map (
            O => \N__11347\,
            I => \N__11294\
        );

    \I__1716\ : InMux
    port map (
            O => \N__11344\,
            I => \N__11294\
        );

    \I__1715\ : InMux
    port map (
            O => \N__11341\,
            I => \N__11294\
        );

    \I__1714\ : InMux
    port map (
            O => \N__11338\,
            I => \N__11294\
        );

    \I__1713\ : InMux
    port map (
            O => \N__11337\,
            I => \N__11283\
        );

    \I__1712\ : InMux
    port map (
            O => \N__11334\,
            I => \N__11283\
        );

    \I__1711\ : InMux
    port map (
            O => \N__11333\,
            I => \N__11283\
        );

    \I__1710\ : InMux
    port map (
            O => \N__11332\,
            I => \N__11283\
        );

    \I__1709\ : InMux
    port map (
            O => \N__11331\,
            I => \N__11283\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__11326\,
            I => \N__11280\
        );

    \I__1707\ : InMux
    port map (
            O => \N__11325\,
            I => \N__11263\
        );

    \I__1706\ : InMux
    port map (
            O => \N__11324\,
            I => \N__11263\
        );

    \I__1705\ : InMux
    port map (
            O => \N__11323\,
            I => \N__11263\
        );

    \I__1704\ : InMux
    port map (
            O => \N__11322\,
            I => \N__11263\
        );

    \I__1703\ : InMux
    port map (
            O => \N__11319\,
            I => \N__11263\
        );

    \I__1702\ : InMux
    port map (
            O => \N__11316\,
            I => \N__11263\
        );

    \I__1701\ : InMux
    port map (
            O => \N__11313\,
            I => \N__11263\
        );

    \I__1700\ : InMux
    port map (
            O => \N__11312\,
            I => \N__11263\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__11309\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__11294\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__11283\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__1696\ : Odrv4
    port map (
            O => \N__11280\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__11263\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__1694\ : CascadeMux
    port map (
            O => \N__11252\,
            I => \phase_controller_inst1.stoper_tr.un1_startlto9_cZ0_cascade_\
        );

    \I__1693\ : InMux
    port map (
            O => \N__11249\,
            I => \N__11246\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__11246\,
            I => \phase_controller_inst1.stoper_tr.un1_startlto13\
        );

    \I__1691\ : CascadeMux
    port map (
            O => \N__11243\,
            I => \phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_6_cascade_\
        );

    \I__1690\ : CascadeMux
    port map (
            O => \N__11240\,
            I => \N__11236\
        );

    \I__1689\ : InMux
    port map (
            O => \N__11239\,
            I => \N__11231\
        );

    \I__1688\ : InMux
    port map (
            O => \N__11236\,
            I => \N__11231\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__11231\,
            I => \N__11227\
        );

    \I__1686\ : CascadeMux
    port map (
            O => \N__11230\,
            I => \N__11223\
        );

    \I__1685\ : Span4Mux_h
    port map (
            O => \N__11227\,
            I => \N__11220\
        );

    \I__1684\ : InMux
    port map (
            O => \N__11226\,
            I => \N__11215\
        );

    \I__1683\ : InMux
    port map (
            O => \N__11223\,
            I => \N__11215\
        );

    \I__1682\ : Odrv4
    port map (
            O => \N__11220\,
            I => \phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_8\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__11215\,
            I => \phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_8\
        );

    \I__1680\ : CascadeMux
    port map (
            O => \N__11210\,
            I => \phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_8_cascade_\
        );

    \I__1679\ : CascadeMux
    port map (
            O => \N__11207\,
            I => \N__11203\
        );

    \I__1678\ : CascadeMux
    port map (
            O => \N__11206\,
            I => \N__11199\
        );

    \I__1677\ : InMux
    port map (
            O => \N__11203\,
            I => \N__11195\
        );

    \I__1676\ : InMux
    port map (
            O => \N__11202\,
            I => \N__11192\
        );

    \I__1675\ : InMux
    port map (
            O => \N__11199\,
            I => \N__11187\
        );

    \I__1674\ : InMux
    port map (
            O => \N__11198\,
            I => \N__11187\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__11195\,
            I => \N__11182\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__11192\,
            I => \N__11182\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__11187\,
            I => \N__11176\
        );

    \I__1670\ : Span4Mux_h
    port map (
            O => \N__11182\,
            I => \N__11176\
        );

    \I__1669\ : InMux
    port map (
            O => \N__11181\,
            I => \N__11173\
        );

    \I__1668\ : Odrv4
    port map (
            O => \N__11176\,
            I => \phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_9\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__11173\,
            I => \phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_9\
        );

    \I__1666\ : CascadeMux
    port map (
            O => \N__11168\,
            I => \N__11165\
        );

    \I__1665\ : InMux
    port map (
            O => \N__11165\,
            I => \N__11162\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__11162\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNI89DKZ0\
        );

    \I__1663\ : CascadeMux
    port map (
            O => \N__11159\,
            I => \N__11156\
        );

    \I__1662\ : InMux
    port map (
            O => \N__11156\,
            I => \N__11153\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__11153\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10\
        );

    \I__1660\ : InMux
    port map (
            O => \N__11150\,
            I => \N__11147\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__11147\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11\
        );

    \I__1658\ : InMux
    port map (
            O => \N__11144\,
            I => \N__11141\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__11141\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13\
        );

    \I__1656\ : CascadeMux
    port map (
            O => \N__11138\,
            I => \N__11135\
        );

    \I__1655\ : InMux
    port map (
            O => \N__11135\,
            I => \N__11132\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__11132\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14\
        );

    \I__1653\ : InMux
    port map (
            O => \N__11129\,
            I => \N__11126\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__11126\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15\
        );

    \I__1651\ : CascadeMux
    port map (
            O => \N__11123\,
            I => \N__11120\
        );

    \I__1650\ : InMux
    port map (
            O => \N__11120\,
            I => \N__11117\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__11117\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16\
        );

    \I__1648\ : InMux
    port map (
            O => \N__11114\,
            I => \N__11111\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__11111\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17\
        );

    \I__1646\ : InMux
    port map (
            O => \N__11108\,
            I => \N__11105\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__11105\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4\
        );

    \I__1644\ : CascadeMux
    port map (
            O => \N__11102\,
            I => \N__11099\
        );

    \I__1643\ : InMux
    port map (
            O => \N__11099\,
            I => \N__11096\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__11096\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5\
        );

    \I__1641\ : InMux
    port map (
            O => \N__11093\,
            I => \N__11090\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__11090\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6\
        );

    \I__1639\ : CascadeMux
    port map (
            O => \N__11087\,
            I => \N__11084\
        );

    \I__1638\ : InMux
    port map (
            O => \N__11084\,
            I => \N__11081\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__11081\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7\
        );

    \I__1636\ : InMux
    port map (
            O => \N__11078\,
            I => \N__11075\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__11075\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8\
        );

    \I__1634\ : CascadeMux
    port map (
            O => \N__11072\,
            I => \N__11069\
        );

    \I__1633\ : InMux
    port map (
            O => \N__11069\,
            I => \N__11066\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__11066\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9\
        );

    \I__1631\ : CascadeMux
    port map (
            O => \N__11063\,
            I => \N__11060\
        );

    \I__1630\ : InMux
    port map (
            O => \N__11060\,
            I => \N__11057\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__11057\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\
        );

    \I__1628\ : CascadeMux
    port map (
            O => \N__11054\,
            I => \N__11049\
        );

    \I__1627\ : CascadeMux
    port map (
            O => \N__11053\,
            I => \N__11046\
        );

    \I__1626\ : InMux
    port map (
            O => \N__11052\,
            I => \N__11043\
        );

    \I__1625\ : InMux
    port map (
            O => \N__11049\,
            I => \N__11038\
        );

    \I__1624\ : InMux
    port map (
            O => \N__11046\,
            I => \N__11038\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__11043\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__11038\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__1621\ : InMux
    port map (
            O => \N__11033\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__1620\ : CascadeMux
    port map (
            O => \N__11030\,
            I => \N__11025\
        );

    \I__1619\ : CascadeMux
    port map (
            O => \N__11029\,
            I => \N__11022\
        );

    \I__1618\ : InMux
    port map (
            O => \N__11028\,
            I => \N__11019\
        );

    \I__1617\ : InMux
    port map (
            O => \N__11025\,
            I => \N__11014\
        );

    \I__1616\ : InMux
    port map (
            O => \N__11022\,
            I => \N__11014\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__11019\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__11014\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__1613\ : InMux
    port map (
            O => \N__11009\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__1612\ : InMux
    port map (
            O => \N__11006\,
            I => \N__11001\
        );

    \I__1611\ : InMux
    port map (
            O => \N__11005\,
            I => \N__10998\
        );

    \I__1610\ : InMux
    port map (
            O => \N__11004\,
            I => \N__10995\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__11001\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__10998\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__10995\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__1606\ : InMux
    port map (
            O => \N__10988\,
            I => \bfn_8_16_0_\
        );

    \I__1605\ : InMux
    port map (
            O => \N__10985\,
            I => \N__10980\
        );

    \I__1604\ : InMux
    port map (
            O => \N__10984\,
            I => \N__10977\
        );

    \I__1603\ : InMux
    port map (
            O => \N__10983\,
            I => \N__10974\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__10980\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__10977\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__10974\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__1599\ : InMux
    port map (
            O => \N__10967\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__1598\ : InMux
    port map (
            O => \N__10964\,
            I => \N__10960\
        );

    \I__1597\ : InMux
    port map (
            O => \N__10963\,
            I => \N__10957\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__10960\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__10957\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__1594\ : CascadeMux
    port map (
            O => \N__10952\,
            I => \N__10947\
        );

    \I__1593\ : CascadeMux
    port map (
            O => \N__10951\,
            I => \N__10944\
        );

    \I__1592\ : InMux
    port map (
            O => \N__10950\,
            I => \N__10941\
        );

    \I__1591\ : InMux
    port map (
            O => \N__10947\,
            I => \N__10936\
        );

    \I__1590\ : InMux
    port map (
            O => \N__10944\,
            I => \N__10936\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__10941\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__10936\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__1587\ : InMux
    port map (
            O => \N__10931\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__1586\ : InMux
    port map (
            O => \N__10928\,
            I => \N__10924\
        );

    \I__1585\ : InMux
    port map (
            O => \N__10927\,
            I => \N__10921\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__10924\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__10921\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__1582\ : CascadeMux
    port map (
            O => \N__10916\,
            I => \N__10911\
        );

    \I__1581\ : CascadeMux
    port map (
            O => \N__10915\,
            I => \N__10908\
        );

    \I__1580\ : InMux
    port map (
            O => \N__10914\,
            I => \N__10905\
        );

    \I__1579\ : InMux
    port map (
            O => \N__10911\,
            I => \N__10900\
        );

    \I__1578\ : InMux
    port map (
            O => \N__10908\,
            I => \N__10900\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__10905\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__10900\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__1575\ : InMux
    port map (
            O => \N__10895\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__1574\ : InMux
    port map (
            O => \N__10892\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__1573\ : CEMux
    port map (
            O => \N__10889\,
            I => \N__10874\
        );

    \I__1572\ : CEMux
    port map (
            O => \N__10888\,
            I => \N__10874\
        );

    \I__1571\ : CEMux
    port map (
            O => \N__10887\,
            I => \N__10874\
        );

    \I__1570\ : CEMux
    port map (
            O => \N__10886\,
            I => \N__10874\
        );

    \I__1569\ : CEMux
    port map (
            O => \N__10885\,
            I => \N__10874\
        );

    \I__1568\ : GlobalMux
    port map (
            O => \N__10874\,
            I => \N__10871\
        );

    \I__1567\ : gio2CtrlBuf
    port map (
            O => \N__10871\,
            I => \delay_measurement_inst.delay_hc_timer.N_178_i_g\
        );

    \I__1566\ : CascadeMux
    port map (
            O => \N__10868\,
            I => \N__10865\
        );

    \I__1565\ : InMux
    port map (
            O => \N__10865\,
            I => \N__10862\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__10862\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3\
        );

    \I__1563\ : InMux
    port map (
            O => \N__10859\,
            I => \N__10854\
        );

    \I__1562\ : InMux
    port map (
            O => \N__10858\,
            I => \N__10849\
        );

    \I__1561\ : InMux
    port map (
            O => \N__10857\,
            I => \N__10849\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__10854\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__10849\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__1558\ : InMux
    port map (
            O => \N__10844\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__1557\ : CascadeMux
    port map (
            O => \N__10841\,
            I => \N__10836\
        );

    \I__1556\ : CascadeMux
    port map (
            O => \N__10840\,
            I => \N__10833\
        );

    \I__1555\ : InMux
    port map (
            O => \N__10839\,
            I => \N__10830\
        );

    \I__1554\ : InMux
    port map (
            O => \N__10836\,
            I => \N__10825\
        );

    \I__1553\ : InMux
    port map (
            O => \N__10833\,
            I => \N__10825\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__10830\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__10825\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__1550\ : InMux
    port map (
            O => \N__10820\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__1549\ : CascadeMux
    port map (
            O => \N__10817\,
            I => \N__10812\
        );

    \I__1548\ : CascadeMux
    port map (
            O => \N__10816\,
            I => \N__10809\
        );

    \I__1547\ : InMux
    port map (
            O => \N__10815\,
            I => \N__10806\
        );

    \I__1546\ : InMux
    port map (
            O => \N__10812\,
            I => \N__10801\
        );

    \I__1545\ : InMux
    port map (
            O => \N__10809\,
            I => \N__10801\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__10806\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__10801\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__1542\ : InMux
    port map (
            O => \N__10796\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__1541\ : InMux
    port map (
            O => \N__10793\,
            I => \N__10788\
        );

    \I__1540\ : InMux
    port map (
            O => \N__10792\,
            I => \N__10785\
        );

    \I__1539\ : InMux
    port map (
            O => \N__10791\,
            I => \N__10782\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__10788\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__10785\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__10782\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__1535\ : InMux
    port map (
            O => \N__10775\,
            I => \bfn_8_15_0_\
        );

    \I__1534\ : InMux
    port map (
            O => \N__10772\,
            I => \N__10767\
        );

    \I__1533\ : InMux
    port map (
            O => \N__10771\,
            I => \N__10764\
        );

    \I__1532\ : InMux
    port map (
            O => \N__10770\,
            I => \N__10761\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__10767\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__10764\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__10761\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__1528\ : InMux
    port map (
            O => \N__10754\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__1527\ : CascadeMux
    port map (
            O => \N__10751\,
            I => \N__10746\
        );

    \I__1526\ : CascadeMux
    port map (
            O => \N__10750\,
            I => \N__10743\
        );

    \I__1525\ : InMux
    port map (
            O => \N__10749\,
            I => \N__10740\
        );

    \I__1524\ : InMux
    port map (
            O => \N__10746\,
            I => \N__10735\
        );

    \I__1523\ : InMux
    port map (
            O => \N__10743\,
            I => \N__10735\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__10740\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__10735\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__1520\ : InMux
    port map (
            O => \N__10730\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__1519\ : CascadeMux
    port map (
            O => \N__10727\,
            I => \N__10722\
        );

    \I__1518\ : CascadeMux
    port map (
            O => \N__10726\,
            I => \N__10719\
        );

    \I__1517\ : InMux
    port map (
            O => \N__10725\,
            I => \N__10716\
        );

    \I__1516\ : InMux
    port map (
            O => \N__10722\,
            I => \N__10711\
        );

    \I__1515\ : InMux
    port map (
            O => \N__10719\,
            I => \N__10711\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__10716\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__10711\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__1512\ : InMux
    port map (
            O => \N__10706\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__1511\ : InMux
    port map (
            O => \N__10703\,
            I => \N__10698\
        );

    \I__1510\ : InMux
    port map (
            O => \N__10702\,
            I => \N__10693\
        );

    \I__1509\ : InMux
    port map (
            O => \N__10701\,
            I => \N__10693\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__10698\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__10693\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__1506\ : InMux
    port map (
            O => \N__10688\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__1505\ : InMux
    port map (
            O => \N__10685\,
            I => \N__10680\
        );

    \I__1504\ : InMux
    port map (
            O => \N__10684\,
            I => \N__10675\
        );

    \I__1503\ : InMux
    port map (
            O => \N__10683\,
            I => \N__10675\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__10680\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__10675\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__1500\ : InMux
    port map (
            O => \N__10670\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__1499\ : InMux
    port map (
            O => \N__10667\,
            I => \N__10662\
        );

    \I__1498\ : InMux
    port map (
            O => \N__10666\,
            I => \N__10657\
        );

    \I__1497\ : InMux
    port map (
            O => \N__10665\,
            I => \N__10657\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__10662\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__10657\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__1494\ : InMux
    port map (
            O => \N__10652\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__1493\ : CascadeMux
    port map (
            O => \N__10649\,
            I => \N__10644\
        );

    \I__1492\ : CascadeMux
    port map (
            O => \N__10648\,
            I => \N__10641\
        );

    \I__1491\ : InMux
    port map (
            O => \N__10647\,
            I => \N__10638\
        );

    \I__1490\ : InMux
    port map (
            O => \N__10644\,
            I => \N__10633\
        );

    \I__1489\ : InMux
    port map (
            O => \N__10641\,
            I => \N__10633\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__10638\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__10633\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__1486\ : InMux
    port map (
            O => \N__10628\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__1485\ : CascadeMux
    port map (
            O => \N__10625\,
            I => \N__10620\
        );

    \I__1484\ : CascadeMux
    port map (
            O => \N__10624\,
            I => \N__10617\
        );

    \I__1483\ : InMux
    port map (
            O => \N__10623\,
            I => \N__10614\
        );

    \I__1482\ : InMux
    port map (
            O => \N__10620\,
            I => \N__10609\
        );

    \I__1481\ : InMux
    port map (
            O => \N__10617\,
            I => \N__10609\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__10614\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__10609\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__1478\ : InMux
    port map (
            O => \N__10604\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__1477\ : InMux
    port map (
            O => \N__10601\,
            I => \N__10596\
        );

    \I__1476\ : InMux
    port map (
            O => \N__10600\,
            I => \N__10593\
        );

    \I__1475\ : InMux
    port map (
            O => \N__10599\,
            I => \N__10590\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__10596\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__10593\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__10590\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__1471\ : InMux
    port map (
            O => \N__10583\,
            I => \bfn_8_14_0_\
        );

    \I__1470\ : InMux
    port map (
            O => \N__10580\,
            I => \N__10575\
        );

    \I__1469\ : InMux
    port map (
            O => \N__10579\,
            I => \N__10572\
        );

    \I__1468\ : InMux
    port map (
            O => \N__10578\,
            I => \N__10569\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__10575\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__10572\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__10569\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__1464\ : InMux
    port map (
            O => \N__10562\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__1463\ : CascadeMux
    port map (
            O => \N__10559\,
            I => \N__10554\
        );

    \I__1462\ : CascadeMux
    port map (
            O => \N__10558\,
            I => \N__10551\
        );

    \I__1461\ : InMux
    port map (
            O => \N__10557\,
            I => \N__10548\
        );

    \I__1460\ : InMux
    port map (
            O => \N__10554\,
            I => \N__10543\
        );

    \I__1459\ : InMux
    port map (
            O => \N__10551\,
            I => \N__10543\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__10548\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__10543\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__1456\ : InMux
    port map (
            O => \N__10538\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__1455\ : CascadeMux
    port map (
            O => \N__10535\,
            I => \N__10530\
        );

    \I__1454\ : CascadeMux
    port map (
            O => \N__10534\,
            I => \N__10527\
        );

    \I__1453\ : InMux
    port map (
            O => \N__10533\,
            I => \N__10524\
        );

    \I__1452\ : InMux
    port map (
            O => \N__10530\,
            I => \N__10519\
        );

    \I__1451\ : InMux
    port map (
            O => \N__10527\,
            I => \N__10519\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__10524\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__10519\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__1448\ : InMux
    port map (
            O => \N__10514\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__1447\ : InMux
    port map (
            O => \N__10511\,
            I => \N__10506\
        );

    \I__1446\ : InMux
    port map (
            O => \N__10510\,
            I => \N__10501\
        );

    \I__1445\ : InMux
    port map (
            O => \N__10509\,
            I => \N__10501\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__10506\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__10501\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__1442\ : InMux
    port map (
            O => \N__10496\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__1441\ : CascadeMux
    port map (
            O => \N__10493\,
            I => \delay_measurement_inst.delay_hc_timer.N_105_cascade_\
        );

    \I__1440\ : InMux
    port map (
            O => \N__10490\,
            I => \N__10485\
        );

    \I__1439\ : InMux
    port map (
            O => \N__10489\,
            I => \N__10482\
        );

    \I__1438\ : InMux
    port map (
            O => \N__10488\,
            I => \N__10479\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__10485\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__10482\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__10479\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__1434\ : InMux
    port map (
            O => \N__10472\,
            I => \N__10467\
        );

    \I__1433\ : InMux
    port map (
            O => \N__10471\,
            I => \N__10464\
        );

    \I__1432\ : InMux
    port map (
            O => \N__10470\,
            I => \N__10461\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__10467\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__10464\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__10461\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__1428\ : InMux
    port map (
            O => \N__10454\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__1427\ : CascadeMux
    port map (
            O => \N__10451\,
            I => \N__10446\
        );

    \I__1426\ : CascadeMux
    port map (
            O => \N__10450\,
            I => \N__10443\
        );

    \I__1425\ : InMux
    port map (
            O => \N__10449\,
            I => \N__10440\
        );

    \I__1424\ : InMux
    port map (
            O => \N__10446\,
            I => \N__10435\
        );

    \I__1423\ : InMux
    port map (
            O => \N__10443\,
            I => \N__10435\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__10440\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__10435\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__1420\ : InMux
    port map (
            O => \N__10430\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__1419\ : CascadeMux
    port map (
            O => \N__10427\,
            I => \N__10422\
        );

    \I__1418\ : CascadeMux
    port map (
            O => \N__10426\,
            I => \N__10419\
        );

    \I__1417\ : InMux
    port map (
            O => \N__10425\,
            I => \N__10416\
        );

    \I__1416\ : InMux
    port map (
            O => \N__10422\,
            I => \N__10411\
        );

    \I__1415\ : InMux
    port map (
            O => \N__10419\,
            I => \N__10411\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__10416\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__10411\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__1412\ : InMux
    port map (
            O => \N__10406\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__1411\ : InMux
    port map (
            O => \N__10403\,
            I => \N__10398\
        );

    \I__1410\ : InMux
    port map (
            O => \N__10402\,
            I => \N__10393\
        );

    \I__1409\ : InMux
    port map (
            O => \N__10401\,
            I => \N__10393\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__10398\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__10393\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__1406\ : InMux
    port map (
            O => \N__10388\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__1405\ : InMux
    port map (
            O => \N__10385\,
            I => \N__10382\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__10382\,
            I => \N__10379\
        );

    \I__1403\ : Odrv12
    port map (
            O => \N__10379\,
            I => il_max_comp1_c
        );

    \I__1402\ : InMux
    port map (
            O => \N__10376\,
            I => \N__10373\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__10373\,
            I => \N__10370\
        );

    \I__1400\ : Span4Mux_h
    port map (
            O => \N__10370\,
            I => \N__10367\
        );

    \I__1399\ : Odrv4
    port map (
            O => \N__10367\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\
        );

    \I__1398\ : CascadeMux
    port map (
            O => \N__10364\,
            I => \N__10361\
        );

    \I__1397\ : InMux
    port map (
            O => \N__10361\,
            I => \N__10358\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__10358\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\
        );

    \I__1395\ : CascadeMux
    port map (
            O => \N__10355\,
            I => \N__10352\
        );

    \I__1394\ : InMux
    port map (
            O => \N__10352\,
            I => \N__10349\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__10349\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_16\
        );

    \I__1392\ : CascadeMux
    port map (
            O => \N__10346\,
            I => \N__10343\
        );

    \I__1391\ : InMux
    port map (
            O => \N__10343\,
            I => \N__10340\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__10340\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_17\
        );

    \I__1389\ : InMux
    port map (
            O => \N__10337\,
            I => \N__10334\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__10334\,
            I => \N__10331\
        );

    \I__1387\ : Odrv4
    port map (
            O => \N__10331\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\
        );

    \I__1386\ : CascadeMux
    port map (
            O => \N__10328\,
            I => \N__10325\
        );

    \I__1385\ : InMux
    port map (
            O => \N__10325\,
            I => \N__10322\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__10322\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_18\
        );

    \I__1383\ : InMux
    port map (
            O => \N__10319\,
            I => \N__10316\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__10316\,
            I => \N__10313\
        );

    \I__1381\ : Span4Mux_h
    port map (
            O => \N__10313\,
            I => \N__10310\
        );

    \I__1380\ : Odrv4
    port map (
            O => \N__10310\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\
        );

    \I__1379\ : CascadeMux
    port map (
            O => \N__10307\,
            I => \N__10304\
        );

    \I__1378\ : InMux
    port map (
            O => \N__10304\,
            I => \N__10301\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__10301\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_19\
        );

    \I__1376\ : InMux
    port map (
            O => \N__10298\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__1375\ : CascadeMux
    port map (
            O => \N__10295\,
            I => \N__10292\
        );

    \I__1374\ : InMux
    port map (
            O => \N__10292\,
            I => \N__10289\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__10289\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\
        );

    \I__1372\ : CascadeMux
    port map (
            O => \N__10286\,
            I => \N__10283\
        );

    \I__1371\ : InMux
    port map (
            O => \N__10283\,
            I => \N__10280\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__10280\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\
        );

    \I__1369\ : InMux
    port map (
            O => \N__10277\,
            I => \N__10274\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__10274\,
            I => \N__10271\
        );

    \I__1367\ : Odrv12
    port map (
            O => \N__10271\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\
        );

    \I__1366\ : CascadeMux
    port map (
            O => \N__10268\,
            I => \N__10265\
        );

    \I__1365\ : InMux
    port map (
            O => \N__10265\,
            I => \N__10262\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__10262\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\
        );

    \I__1363\ : InMux
    port map (
            O => \N__10259\,
            I => \N__10256\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__10256\,
            I => \N__10253\
        );

    \I__1361\ : Span4Mux_h
    port map (
            O => \N__10253\,
            I => \N__10250\
        );

    \I__1360\ : Odrv4
    port map (
            O => \N__10250\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\
        );

    \I__1359\ : CascadeMux
    port map (
            O => \N__10247\,
            I => \N__10244\
        );

    \I__1358\ : InMux
    port map (
            O => \N__10244\,
            I => \N__10241\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__10241\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\
        );

    \I__1356\ : InMux
    port map (
            O => \N__10238\,
            I => \N__10235\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__10235\,
            I => \N__10232\
        );

    \I__1354\ : Odrv12
    port map (
            O => \N__10232\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\
        );

    \I__1353\ : CascadeMux
    port map (
            O => \N__10229\,
            I => \N__10226\
        );

    \I__1352\ : InMux
    port map (
            O => \N__10226\,
            I => \N__10223\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__10223\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\
        );

    \I__1350\ : InMux
    port map (
            O => \N__10220\,
            I => \N__10217\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__10217\,
            I => \N__10214\
        );

    \I__1348\ : Span4Mux_h
    port map (
            O => \N__10214\,
            I => \N__10211\
        );

    \I__1347\ : Odrv4
    port map (
            O => \N__10211\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\
        );

    \I__1346\ : CascadeMux
    port map (
            O => \N__10208\,
            I => \N__10205\
        );

    \I__1345\ : InMux
    port map (
            O => \N__10205\,
            I => \N__10202\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__10202\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\
        );

    \I__1343\ : InMux
    port map (
            O => \N__10199\,
            I => \N__10196\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__10196\,
            I => \N__10193\
        );

    \I__1341\ : Odrv4
    port map (
            O => \N__10193\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\
        );

    \I__1340\ : CascadeMux
    port map (
            O => \N__10190\,
            I => \N__10187\
        );

    \I__1339\ : InMux
    port map (
            O => \N__10187\,
            I => \N__10184\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__10184\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\
        );

    \I__1337\ : InMux
    port map (
            O => \N__10181\,
            I => \N__10178\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__10178\,
            I => \N__10175\
        );

    \I__1335\ : Span4Mux_v
    port map (
            O => \N__10175\,
            I => \N__10172\
        );

    \I__1334\ : Odrv4
    port map (
            O => \N__10172\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\
        );

    \I__1333\ : CascadeMux
    port map (
            O => \N__10169\,
            I => \N__10166\
        );

    \I__1332\ : InMux
    port map (
            O => \N__10166\,
            I => \N__10163\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__10163\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\
        );

    \I__1330\ : InMux
    port map (
            O => \N__10160\,
            I => \N__10152\
        );

    \I__1329\ : InMux
    port map (
            O => \N__10159\,
            I => \N__10152\
        );

    \I__1328\ : InMux
    port map (
            O => \N__10158\,
            I => \N__10147\
        );

    \I__1327\ : InMux
    port map (
            O => \N__10157\,
            I => \N__10147\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__10152\,
            I => \N__10144\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__10147\,
            I => \N__10141\
        );

    \I__1324\ : Odrv4
    port map (
            O => \N__10144\,
            I => \phase_controller_inst1.stoper_tr.un1_start\
        );

    \I__1323\ : Odrv4
    port map (
            O => \N__10141\,
            I => \phase_controller_inst1.stoper_tr.un1_start\
        );

    \I__1322\ : InMux
    port map (
            O => \N__10136\,
            I => \N__10133\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__10133\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\
        );

    \I__1320\ : CascadeMux
    port map (
            O => \N__10130\,
            I => \N__10127\
        );

    \I__1319\ : InMux
    port map (
            O => \N__10127\,
            I => \N__10124\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__10124\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\
        );

    \I__1317\ : InMux
    port map (
            O => \N__10121\,
            I => \N__10118\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__10118\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\
        );

    \I__1315\ : CascadeMux
    port map (
            O => \N__10115\,
            I => \N__10112\
        );

    \I__1314\ : InMux
    port map (
            O => \N__10112\,
            I => \N__10109\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__10109\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\
        );

    \I__1312\ : InMux
    port map (
            O => \N__10106\,
            I => \N__10103\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__10103\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\
        );

    \I__1310\ : CascadeMux
    port map (
            O => \N__10100\,
            I => \N__10097\
        );

    \I__1309\ : InMux
    port map (
            O => \N__10097\,
            I => \N__10094\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__10094\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\
        );

    \I__1307\ : CascadeMux
    port map (
            O => \N__10091\,
            I => \N__10088\
        );

    \I__1306\ : InMux
    port map (
            O => \N__10088\,
            I => \N__10085\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__10085\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\
        );

    \I__1304\ : InMux
    port map (
            O => \N__10082\,
            I => \N__10079\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__10079\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\
        );

    \I__1302\ : CascadeMux
    port map (
            O => \N__10076\,
            I => \N__10073\
        );

    \I__1301\ : InMux
    port map (
            O => \N__10073\,
            I => \N__10070\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__10070\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\
        );

    \I__1299\ : InMux
    port map (
            O => \N__10067\,
            I => \N__10064\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__10064\,
            I => \N__10061\
        );

    \I__1297\ : Odrv4
    port map (
            O => \N__10061\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ1Z_6\
        );

    \I__1296\ : CascadeMux
    port map (
            O => \N__10058\,
            I => \N__10055\
        );

    \I__1295\ : InMux
    port map (
            O => \N__10055\,
            I => \N__10052\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__10052\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\
        );

    \I__1293\ : CascadeMux
    port map (
            O => \N__10049\,
            I => \phase_controller_inst1.stoper_tr.un2_startlto6Z0Z_0_cascade_\
        );

    \I__1292\ : InMux
    port map (
            O => \N__10046\,
            I => \N__10043\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__10043\,
            I => \phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_4\
        );

    \I__1290\ : CascadeMux
    port map (
            O => \N__10040\,
            I => \phase_controller_inst1.stoper_tr.un2_startlt19_0_cascade_\
        );

    \I__1289\ : InMux
    port map (
            O => \N__10037\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14\
        );

    \I__1288\ : InMux
    port map (
            O => \N__10034\,
            I => \bfn_7_19_0_\
        );

    \I__1287\ : InMux
    port map (
            O => \N__10031\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16\
        );

    \I__1286\ : InMux
    port map (
            O => \N__10028\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17\
        );

    \I__1285\ : CascadeMux
    port map (
            O => \N__10025\,
            I => \phase_controller_inst1.stoper_tr.un1_startlt8_cascade_\
        );

    \I__1284\ : InMux
    port map (
            O => \N__10022\,
            I => \N__10019\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__10019\,
            I => \phase_controller_inst1.stoper_tr.un1_startlto5Z0Z_1\
        );

    \I__1282\ : InMux
    port map (
            O => \N__10016\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5\
        );

    \I__1281\ : InMux
    port map (
            O => \N__10013\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6\
        );

    \I__1280\ : InMux
    port map (
            O => \N__10010\,
            I => \bfn_7_18_0_\
        );

    \I__1279\ : InMux
    port map (
            O => \N__10007\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8\
        );

    \I__1278\ : InMux
    port map (
            O => \N__10004\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9\
        );

    \I__1277\ : InMux
    port map (
            O => \N__10001\,
            I => \N__9998\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__9998\,
            I => \N__9995\
        );

    \I__1275\ : Odrv4
    port map (
            O => \N__9995\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12\
        );

    \I__1274\ : InMux
    port map (
            O => \N__9992\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10\
        );

    \I__1273\ : InMux
    port map (
            O => \N__9989\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11\
        );

    \I__1272\ : InMux
    port map (
            O => \N__9986\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12\
        );

    \I__1271\ : InMux
    port map (
            O => \N__9983\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13\
        );

    \I__1270\ : InMux
    port map (
            O => \N__9980\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_26\
        );

    \I__1269\ : InMux
    port map (
            O => \N__9977\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_27\
        );

    \I__1268\ : InMux
    port map (
            O => \N__9974\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_28\
        );

    \I__1267\ : InMux
    port map (
            O => \N__9971\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0\
        );

    \I__1266\ : InMux
    port map (
            O => \N__9968\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1\
        );

    \I__1265\ : InMux
    port map (
            O => \N__9965\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2\
        );

    \I__1264\ : InMux
    port map (
            O => \N__9962\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3\
        );

    \I__1263\ : InMux
    port map (
            O => \N__9959\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4\
        );

    \I__1262\ : InMux
    port map (
            O => \N__9956\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_17\
        );

    \I__1261\ : InMux
    port map (
            O => \N__9953\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_18\
        );

    \I__1260\ : InMux
    port map (
            O => \N__9950\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_19\
        );

    \I__1259\ : InMux
    port map (
            O => \N__9947\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_20\
        );

    \I__1258\ : InMux
    port map (
            O => \N__9944\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_21\
        );

    \I__1257\ : InMux
    port map (
            O => \N__9941\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_22\
        );

    \I__1256\ : InMux
    port map (
            O => \N__9938\,
            I => \bfn_7_16_0_\
        );

    \I__1255\ : InMux
    port map (
            O => \N__9935\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_24\
        );

    \I__1254\ : InMux
    port map (
            O => \N__9932\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_25\
        );

    \I__1253\ : InMux
    port map (
            O => \N__9929\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_8\
        );

    \I__1252\ : InMux
    port map (
            O => \N__9926\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_9\
        );

    \I__1251\ : InMux
    port map (
            O => \N__9923\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_10\
        );

    \I__1250\ : InMux
    port map (
            O => \N__9920\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_11\
        );

    \I__1249\ : InMux
    port map (
            O => \N__9917\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_12\
        );

    \I__1248\ : InMux
    port map (
            O => \N__9914\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_13\
        );

    \I__1247\ : InMux
    port map (
            O => \N__9911\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_14\
        );

    \I__1246\ : InMux
    port map (
            O => \N__9908\,
            I => \bfn_7_15_0_\
        );

    \I__1245\ : InMux
    port map (
            O => \N__9905\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_16\
        );

    \I__1244\ : InMux
    port map (
            O => \N__9902\,
            I => \bfn_7_13_0_\
        );

    \I__1243\ : InMux
    port map (
            O => \N__9899\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_0\
        );

    \I__1242\ : InMux
    port map (
            O => \N__9896\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_1\
        );

    \I__1241\ : InMux
    port map (
            O => \N__9893\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_2\
        );

    \I__1240\ : InMux
    port map (
            O => \N__9890\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_3\
        );

    \I__1239\ : InMux
    port map (
            O => \N__9887\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_4\
        );

    \I__1238\ : InMux
    port map (
            O => \N__9884\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_5\
        );

    \I__1237\ : InMux
    port map (
            O => \N__9881\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_6\
        );

    \I__1236\ : InMux
    port map (
            O => \N__9878\,
            I => \bfn_7_14_0_\
        );

    \I__1235\ : CascadeMux
    port map (
            O => \N__9875\,
            I => \N__9872\
        );

    \I__1234\ : InMux
    port map (
            O => \N__9872\,
            I => \N__9869\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__9869\,
            I => \phase_controller_slave.stoper_hc.N_60\
        );

    \I__1232\ : InMux
    port map (
            O => \N__9866\,
            I => \N__9858\
        );

    \I__1231\ : InMux
    port map (
            O => \N__9865\,
            I => \N__9858\
        );

    \I__1230\ : InMux
    port map (
            O => \N__9864\,
            I => \N__9855\
        );

    \I__1229\ : InMux
    port map (
            O => \N__9863\,
            I => \N__9852\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__9858\,
            I => \N__9847\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__9855\,
            I => \N__9847\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__9852\,
            I => \phase_controller_slave.hc_time_passed\
        );

    \I__1225\ : Odrv4
    port map (
            O => \N__9847\,
            I => \phase_controller_slave.hc_time_passed\
        );

    \I__1224\ : InMux
    port map (
            O => \N__9842\,
            I => \N__9839\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__9839\,
            I => \N__9835\
        );

    \I__1222\ : InMux
    port map (
            O => \N__9838\,
            I => \N__9832\
        );

    \I__1221\ : Odrv4
    port map (
            O => \N__9835\,
            I => \phase_controller_slave.state_RNIVDE2Z0Z_0\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__9832\,
            I => \phase_controller_slave.state_RNIVDE2Z0Z_0\
        );

    \I__1219\ : CascadeMux
    port map (
            O => \N__9827\,
            I => \N__9824\
        );

    \I__1218\ : InMux
    port map (
            O => \N__9824\,
            I => \N__9819\
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__9823\,
            I => \N__9816\
        );

    \I__1216\ : CascadeMux
    port map (
            O => \N__9822\,
            I => \N__9813\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__9819\,
            I => \N__9809\
        );

    \I__1214\ : InMux
    port map (
            O => \N__9816\,
            I => \N__9806\
        );

    \I__1213\ : InMux
    port map (
            O => \N__9813\,
            I => \N__9801\
        );

    \I__1212\ : InMux
    port map (
            O => \N__9812\,
            I => \N__9801\
        );

    \I__1211\ : Span4Mux_h
    port map (
            O => \N__9809\,
            I => \N__9798\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__9806\,
            I => \N__9795\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__9801\,
            I => \N__9792\
        );

    \I__1208\ : Odrv4
    port map (
            O => \N__9798\,
            I => \phase_controller_slave.stateZ0Z_4\
        );

    \I__1207\ : Odrv4
    port map (
            O => \N__9795\,
            I => \phase_controller_slave.stateZ0Z_4\
        );

    \I__1206\ : Odrv4
    port map (
            O => \N__9792\,
            I => \phase_controller_slave.stateZ0Z_4\
        );

    \I__1205\ : InMux
    port map (
            O => \N__9785\,
            I => \N__9782\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__9782\,
            I => \phase_controller_slave.state_RNO_0Z0Z_3\
        );

    \I__1203\ : InMux
    port map (
            O => \N__9779\,
            I => \N__9775\
        );

    \I__1202\ : CascadeMux
    port map (
            O => \N__9778\,
            I => \N__9772\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__9775\,
            I => \N__9768\
        );

    \I__1200\ : InMux
    port map (
            O => \N__9772\,
            I => \N__9765\
        );

    \I__1199\ : InMux
    port map (
            O => \N__9771\,
            I => \N__9762\
        );

    \I__1198\ : Odrv4
    port map (
            O => \N__9768\,
            I => shift_flag_start
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__9765\,
            I => shift_flag_start
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__9762\,
            I => shift_flag_start
        );

    \I__1195\ : InMux
    port map (
            O => \N__9755\,
            I => \N__9752\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__9752\,
            I => \N__9746\
        );

    \I__1193\ : InMux
    port map (
            O => \N__9751\,
            I => \N__9743\
        );

    \I__1192\ : InMux
    port map (
            O => \N__9750\,
            I => \N__9740\
        );

    \I__1191\ : InMux
    port map (
            O => \N__9749\,
            I => \N__9737\
        );

    \I__1190\ : Odrv12
    port map (
            O => \N__9746\,
            I => \phase_controller_slave.stateZ0Z_1\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__9743\,
            I => \phase_controller_slave.stateZ0Z_1\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__9740\,
            I => \phase_controller_slave.stateZ0Z_1\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__9737\,
            I => \phase_controller_slave.stateZ0Z_1\
        );

    \I__1186\ : IoInMux
    port map (
            O => \N__9728\,
            I => \N__9725\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__9725\,
            I => \N__9722\
        );

    \I__1184\ : IoSpan4Mux
    port map (
            O => \N__9722\,
            I => \N__9719\
        );

    \I__1183\ : Span4Mux_s2_v
    port map (
            O => \N__9719\,
            I => \N__9716\
        );

    \I__1182\ : Span4Mux_v
    port map (
            O => \N__9716\,
            I => \N__9713\
        );

    \I__1181\ : Odrv4
    port map (
            O => \N__9713\,
            I => s4_phy_c
        );

    \I__1180\ : InMux
    port map (
            O => \N__9710\,
            I => \N__9707\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__9707\,
            I => \N__9704\
        );

    \I__1178\ : Odrv4
    port map (
            O => \N__9704\,
            I => \il_max_comp2_D1\
        );

    \I__1177\ : InMux
    port map (
            O => \N__9701\,
            I => \N__9698\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__9698\,
            I => \N__9695\
        );

    \I__1175\ : Odrv4
    port map (
            O => \N__9695\,
            I => \phase_controller_slave.start_timer_hc_0_sqmuxa\
        );

    \I__1174\ : InMux
    port map (
            O => \N__9692\,
            I => \N__9689\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__9689\,
            I => \phase_controller_slave.start_timer_hc_RNOZ0Z_0\
        );

    \I__1172\ : InMux
    port map (
            O => \N__9686\,
            I => \N__9681\
        );

    \I__1171\ : InMux
    port map (
            O => \N__9685\,
            I => \N__9678\
        );

    \I__1170\ : InMux
    port map (
            O => \N__9684\,
            I => \N__9675\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__9681\,
            I => \N__9668\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__9678\,
            I => \N__9668\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__9675\,
            I => \N__9668\
        );

    \I__1166\ : Span4Mux_v
    port map (
            O => \N__9668\,
            I => \N__9665\
        );

    \I__1165\ : Odrv4
    port map (
            O => \N__9665\,
            I => \il_min_comp2_D2\
        );

    \I__1164\ : CascadeMux
    port map (
            O => \N__9662\,
            I => \N__9659\
        );

    \I__1163\ : InMux
    port map (
            O => \N__9659\,
            I => \N__9652\
        );

    \I__1162\ : InMux
    port map (
            O => \N__9658\,
            I => \N__9652\
        );

    \I__1161\ : InMux
    port map (
            O => \N__9657\,
            I => \N__9649\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__9652\,
            I => \phase_controller_slave.stateZ0Z_2\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__9649\,
            I => \phase_controller_slave.stateZ0Z_2\
        );

    \I__1158\ : InMux
    port map (
            O => \N__9644\,
            I => \N__9640\
        );

    \I__1157\ : InMux
    port map (
            O => \N__9643\,
            I => \N__9637\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__9640\,
            I => \N__9631\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__9637\,
            I => \N__9631\
        );

    \I__1154\ : InMux
    port map (
            O => \N__9636\,
            I => \N__9628\
        );

    \I__1153\ : Odrv12
    port map (
            O => \N__9631\,
            I => \il_max_comp2_D2\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__9628\,
            I => \il_max_comp2_D2\
        );

    \I__1151\ : InMux
    port map (
            O => \N__9623\,
            I => \N__9620\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__9620\,
            I => \N__9617\
        );

    \I__1149\ : Odrv4
    port map (
            O => \N__9617\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_16\
        );

    \I__1148\ : InMux
    port map (
            O => \N__9614\,
            I => \N__9611\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__9611\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_11\
        );

    \I__1146\ : InMux
    port map (
            O => \N__9608\,
            I => \N__9605\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__9605\,
            I => \N__9602\
        );

    \I__1144\ : Odrv4
    port map (
            O => \N__9602\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_10\
        );

    \I__1143\ : InMux
    port map (
            O => \N__9599\,
            I => \N__9596\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__9596\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_12\
        );

    \I__1141\ : InMux
    port map (
            O => \N__9593\,
            I => \N__9590\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__9590\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_19\
        );

    \I__1139\ : CEMux
    port map (
            O => \N__9587\,
            I => \N__9584\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__9584\,
            I => \N__9579\
        );

    \I__1137\ : CEMux
    port map (
            O => \N__9583\,
            I => \N__9576\
        );

    \I__1136\ : CEMux
    port map (
            O => \N__9582\,
            I => \N__9572\
        );

    \I__1135\ : Span4Mux_h
    port map (
            O => \N__9579\,
            I => \N__9567\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__9576\,
            I => \N__9567\
        );

    \I__1133\ : CEMux
    port map (
            O => \N__9575\,
            I => \N__9564\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__9572\,
            I => \N__9561\
        );

    \I__1131\ : Span4Mux_v
    port map (
            O => \N__9567\,
            I => \N__9558\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__9564\,
            I => \N__9555\
        );

    \I__1129\ : Span4Mux_h
    port map (
            O => \N__9561\,
            I => \N__9552\
        );

    \I__1128\ : Span4Mux_h
    port map (
            O => \N__9558\,
            I => \N__9549\
        );

    \I__1127\ : Span4Mux_h
    port map (
            O => \N__9555\,
            I => \N__9546\
        );

    \I__1126\ : Odrv4
    port map (
            O => \N__9552\,
            I => \phase_controller_slave.stoper_tr.stoper_state_RNII60DZ0Z_1\
        );

    \I__1125\ : Odrv4
    port map (
            O => \N__9549\,
            I => \phase_controller_slave.stoper_tr.stoper_state_RNII60DZ0Z_1\
        );

    \I__1124\ : Odrv4
    port map (
            O => \N__9546\,
            I => \phase_controller_slave.stoper_tr.stoper_state_RNII60DZ0Z_1\
        );

    \I__1123\ : InMux
    port map (
            O => \N__9539\,
            I => \N__9536\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__9536\,
            I => \N__9533\
        );

    \I__1121\ : Span12Mux_v
    port map (
            O => \N__9533\,
            I => \N__9530\
        );

    \I__1120\ : Odrv12
    port map (
            O => \N__9530\,
            I => il_max_comp2_c
        );

    \I__1119\ : InMux
    port map (
            O => \N__9527\,
            I => \N__9524\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__9524\,
            I => \N__9521\
        );

    \I__1117\ : Span4Mux_h
    port map (
            O => \N__9521\,
            I => \N__9518\
        );

    \I__1116\ : Span4Mux_v
    port map (
            O => \N__9518\,
            I => \N__9515\
        );

    \I__1115\ : Span4Mux_v
    port map (
            O => \N__9515\,
            I => \N__9512\
        );

    \I__1114\ : Odrv4
    port map (
            O => \N__9512\,
            I => il_min_comp2_c
        );

    \I__1113\ : InMux
    port map (
            O => \N__9509\,
            I => \N__9506\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__9506\,
            I => \il_min_comp2_D1\
        );

    \I__1111\ : InMux
    port map (
            O => \N__9503\,
            I => \N__9500\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__9500\,
            I => \N__9497\
        );

    \I__1109\ : Odrv4
    port map (
            O => \N__9497\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_2\
        );

    \I__1108\ : InMux
    port map (
            O => \N__9494\,
            I => \N__9491\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__9491\,
            I => \N__9488\
        );

    \I__1106\ : Odrv4
    port map (
            O => \N__9488\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_13\
        );

    \I__1105\ : InMux
    port map (
            O => \N__9485\,
            I => \N__9482\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__9482\,
            I => \N__9479\
        );

    \I__1103\ : Odrv4
    port map (
            O => \N__9479\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_5\
        );

    \I__1102\ : InMux
    port map (
            O => \N__9476\,
            I => \N__9473\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__9473\,
            I => \N__9470\
        );

    \I__1100\ : Span4Mux_h
    port map (
            O => \N__9470\,
            I => \N__9467\
        );

    \I__1099\ : Odrv4
    port map (
            O => \N__9467\,
            I => \phase_controller_slave.stoper_tr.target_timeZ1Z_6\
        );

    \I__1098\ : InMux
    port map (
            O => \N__9464\,
            I => \N__9461\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__9461\,
            I => \N__9458\
        );

    \I__1096\ : Odrv4
    port map (
            O => \N__9458\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_14\
        );

    \I__1095\ : InMux
    port map (
            O => \N__9455\,
            I => \N__9452\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__9452\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_15\
        );

    \I__1093\ : InMux
    port map (
            O => \N__9449\,
            I => \N__9446\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__9446\,
            I => \N__9443\
        );

    \I__1091\ : Span4Mux_v
    port map (
            O => \N__9443\,
            I => \N__9440\
        );

    \I__1090\ : Odrv4
    port map (
            O => \N__9440\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_9\
        );

    \I__1089\ : InMux
    port map (
            O => \N__9437\,
            I => \N__9434\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__9434\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_17\
        );

    \I__1087\ : InMux
    port map (
            O => \N__9431\,
            I => \N__9428\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__9428\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_18\
        );

    \I__1085\ : InMux
    port map (
            O => \N__9425\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__1084\ : InMux
    port map (
            O => \N__9422\,
            I => \N__9419\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__9419\,
            I => \N__9411\
        );

    \I__1082\ : InMux
    port map (
            O => \N__9418\,
            I => \N__9400\
        );

    \I__1081\ : InMux
    port map (
            O => \N__9417\,
            I => \N__9400\
        );

    \I__1080\ : InMux
    port map (
            O => \N__9416\,
            I => \N__9400\
        );

    \I__1079\ : InMux
    port map (
            O => \N__9415\,
            I => \N__9400\
        );

    \I__1078\ : InMux
    port map (
            O => \N__9414\,
            I => \N__9400\
        );

    \I__1077\ : Odrv4
    port map (
            O => \N__9411\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__9400\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__1075\ : CascadeMux
    port map (
            O => \N__9395\,
            I => \N__9392\
        );

    \I__1074\ : InMux
    port map (
            O => \N__9392\,
            I => \N__9387\
        );

    \I__1073\ : InMux
    port map (
            O => \N__9391\,
            I => \N__9384\
        );

    \I__1072\ : InMux
    port map (
            O => \N__9390\,
            I => \N__9381\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__9387\,
            I => \phase_controller_slave.tr_time_passed\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__9384\,
            I => \phase_controller_slave.tr_time_passed\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__9381\,
            I => \phase_controller_slave.tr_time_passed\
        );

    \I__1068\ : InMux
    port map (
            O => \N__9374\,
            I => \N__9370\
        );

    \I__1067\ : InMux
    port map (
            O => \N__9373\,
            I => \N__9367\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__9370\,
            I => \phase_controller_slave.stateZ0Z_0\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__9367\,
            I => \phase_controller_slave.stateZ0Z_0\
        );

    \I__1064\ : InMux
    port map (
            O => \N__9362\,
            I => \N__9359\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__9359\,
            I => \phase_controller_slave.start_timer_tr_0_sqmuxa\
        );

    \I__1062\ : InMux
    port map (
            O => \N__9356\,
            I => \N__9353\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__9353\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_7\
        );

    \I__1060\ : InMux
    port map (
            O => \N__9350\,
            I => \N__9347\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__9347\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_3\
        );

    \I__1058\ : InMux
    port map (
            O => \N__9344\,
            I => \N__9341\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__9341\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_1\
        );

    \I__1056\ : InMux
    port map (
            O => \N__9338\,
            I => \N__9335\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__9335\,
            I => \N__9332\
        );

    \I__1054\ : Odrv4
    port map (
            O => \N__9332\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_8\
        );

    \I__1053\ : InMux
    port map (
            O => \N__9329\,
            I => \N__9326\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__9326\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_4\
        );

    \I__1051\ : InMux
    port map (
            O => \N__9323\,
            I => \N__9319\
        );

    \I__1050\ : InMux
    port map (
            O => \N__9322\,
            I => \N__9316\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__9319\,
            I => \N__9313\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__9316\,
            I => \N__9310\
        );

    \I__1047\ : Span4Mux_v
    port map (
            O => \N__9313\,
            I => \N__9307\
        );

    \I__1046\ : Span4Mux_v
    port map (
            O => \N__9310\,
            I => \N__9304\
        );

    \I__1045\ : Odrv4
    port map (
            O => \N__9307\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__1044\ : Odrv4
    port map (
            O => \N__9304\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__1043\ : CascadeMux
    port map (
            O => \N__9299\,
            I => \N__9296\
        );

    \I__1042\ : InMux
    port map (
            O => \N__9296\,
            I => \N__9293\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__9293\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_12\
        );

    \I__1040\ : InMux
    port map (
            O => \N__9290\,
            I => \N__9286\
        );

    \I__1039\ : InMux
    port map (
            O => \N__9289\,
            I => \N__9283\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__9286\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__9283\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__1036\ : CascadeMux
    port map (
            O => \N__9278\,
            I => \N__9275\
        );

    \I__1035\ : InMux
    port map (
            O => \N__9275\,
            I => \N__9272\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__9272\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_13\
        );

    \I__1033\ : InMux
    port map (
            O => \N__9269\,
            I => \N__9265\
        );

    \I__1032\ : InMux
    port map (
            O => \N__9268\,
            I => \N__9262\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__9265\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__9262\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__1029\ : CascadeMux
    port map (
            O => \N__9257\,
            I => \N__9254\
        );

    \I__1028\ : InMux
    port map (
            O => \N__9254\,
            I => \N__9251\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__9251\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_14\
        );

    \I__1026\ : InMux
    port map (
            O => \N__9248\,
            I => \N__9244\
        );

    \I__1025\ : InMux
    port map (
            O => \N__9247\,
            I => \N__9241\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__9244\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__9241\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__1022\ : CascadeMux
    port map (
            O => \N__9236\,
            I => \N__9233\
        );

    \I__1021\ : InMux
    port map (
            O => \N__9233\,
            I => \N__9230\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__9230\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_15\
        );

    \I__1019\ : InMux
    port map (
            O => \N__9227\,
            I => \N__9223\
        );

    \I__1018\ : InMux
    port map (
            O => \N__9226\,
            I => \N__9220\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__9223\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__9220\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__1015\ : CascadeMux
    port map (
            O => \N__9215\,
            I => \N__9212\
        );

    \I__1014\ : InMux
    port map (
            O => \N__9212\,
            I => \N__9209\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__9209\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_16\
        );

    \I__1012\ : InMux
    port map (
            O => \N__9206\,
            I => \N__9202\
        );

    \I__1011\ : InMux
    port map (
            O => \N__9205\,
            I => \N__9199\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__9202\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__9199\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__1008\ : CascadeMux
    port map (
            O => \N__9194\,
            I => \N__9191\
        );

    \I__1007\ : InMux
    port map (
            O => \N__9191\,
            I => \N__9188\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__9188\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_17\
        );

    \I__1005\ : InMux
    port map (
            O => \N__9185\,
            I => \N__9181\
        );

    \I__1004\ : InMux
    port map (
            O => \N__9184\,
            I => \N__9178\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__9181\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__9178\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__1001\ : CascadeMux
    port map (
            O => \N__9173\,
            I => \N__9170\
        );

    \I__1000\ : InMux
    port map (
            O => \N__9170\,
            I => \N__9167\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__9167\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_18\
        );

    \I__998\ : InMux
    port map (
            O => \N__9164\,
            I => \N__9160\
        );

    \I__997\ : InMux
    port map (
            O => \N__9163\,
            I => \N__9157\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__9160\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__9157\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__994\ : CascadeMux
    port map (
            O => \N__9152\,
            I => \N__9149\
        );

    \I__993\ : InMux
    port map (
            O => \N__9149\,
            I => \N__9146\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__9146\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_19\
        );

    \I__991\ : InMux
    port map (
            O => \N__9143\,
            I => \N__9139\
        );

    \I__990\ : InMux
    port map (
            O => \N__9142\,
            I => \N__9136\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__9139\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__9136\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__987\ : CascadeMux
    port map (
            O => \N__9131\,
            I => \N__9128\
        );

    \I__986\ : InMux
    port map (
            O => \N__9128\,
            I => \N__9125\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__9125\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_4\
        );

    \I__984\ : InMux
    port map (
            O => \N__9122\,
            I => \N__9119\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__9119\,
            I => \N__9115\
        );

    \I__982\ : InMux
    port map (
            O => \N__9118\,
            I => \N__9112\
        );

    \I__981\ : Odrv4
    port map (
            O => \N__9115\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__9112\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__979\ : CascadeMux
    port map (
            O => \N__9107\,
            I => \N__9104\
        );

    \I__978\ : InMux
    port map (
            O => \N__9104\,
            I => \N__9101\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__9101\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_5\
        );

    \I__976\ : CascadeMux
    port map (
            O => \N__9098\,
            I => \N__9095\
        );

    \I__975\ : InMux
    port map (
            O => \N__9095\,
            I => \N__9091\
        );

    \I__974\ : InMux
    port map (
            O => \N__9094\,
            I => \N__9088\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__9091\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__9088\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__971\ : CascadeMux
    port map (
            O => \N__9083\,
            I => \N__9080\
        );

    \I__970\ : InMux
    port map (
            O => \N__9080\,
            I => \N__9077\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__9077\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_6\
        );

    \I__968\ : InMux
    port map (
            O => \N__9074\,
            I => \N__9070\
        );

    \I__967\ : InMux
    port map (
            O => \N__9073\,
            I => \N__9067\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__9070\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__9067\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__964\ : CascadeMux
    port map (
            O => \N__9062\,
            I => \N__9059\
        );

    \I__963\ : InMux
    port map (
            O => \N__9059\,
            I => \N__9056\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__9056\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_7\
        );

    \I__961\ : CascadeMux
    port map (
            O => \N__9053\,
            I => \N__9050\
        );

    \I__960\ : InMux
    port map (
            O => \N__9050\,
            I => \N__9046\
        );

    \I__959\ : InMux
    port map (
            O => \N__9049\,
            I => \N__9043\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__9046\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__9043\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__956\ : CascadeMux
    port map (
            O => \N__9038\,
            I => \N__9035\
        );

    \I__955\ : InMux
    port map (
            O => \N__9035\,
            I => \N__9032\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__9032\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_8\
        );

    \I__953\ : InMux
    port map (
            O => \N__9029\,
            I => \N__9025\
        );

    \I__952\ : InMux
    port map (
            O => \N__9028\,
            I => \N__9022\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__9025\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__9022\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__949\ : CascadeMux
    port map (
            O => \N__9017\,
            I => \N__9014\
        );

    \I__948\ : InMux
    port map (
            O => \N__9014\,
            I => \N__9011\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__9011\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_9\
        );

    \I__946\ : InMux
    port map (
            O => \N__9008\,
            I => \N__9004\
        );

    \I__945\ : InMux
    port map (
            O => \N__9007\,
            I => \N__9001\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__9004\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__9001\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__942\ : CascadeMux
    port map (
            O => \N__8996\,
            I => \N__8993\
        );

    \I__941\ : InMux
    port map (
            O => \N__8993\,
            I => \N__8990\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__8990\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_10\
        );

    \I__939\ : InMux
    port map (
            O => \N__8987\,
            I => \N__8983\
        );

    \I__938\ : InMux
    port map (
            O => \N__8986\,
            I => \N__8980\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__8983\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__8980\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__935\ : CascadeMux
    port map (
            O => \N__8975\,
            I => \N__8972\
        );

    \I__934\ : InMux
    port map (
            O => \N__8972\,
            I => \N__8969\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__8969\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_11\
        );

    \I__932\ : InMux
    port map (
            O => \N__8966\,
            I => \N__8963\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__8963\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18\
        );

    \I__930\ : InMux
    port map (
            O => \N__8960\,
            I => \N__8957\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__8957\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19\
        );

    \I__928\ : CascadeMux
    port map (
            O => \N__8954\,
            I => \N__8942\
        );

    \I__927\ : CascadeMux
    port map (
            O => \N__8953\,
            I => \N__8935\
        );

    \I__926\ : CascadeMux
    port map (
            O => \N__8952\,
            I => \N__8932\
        );

    \I__925\ : CascadeMux
    port map (
            O => \N__8951\,
            I => \N__8929\
        );

    \I__924\ : CascadeMux
    port map (
            O => \N__8950\,
            I => \N__8923\
        );

    \I__923\ : CascadeMux
    port map (
            O => \N__8949\,
            I => \N__8920\
        );

    \I__922\ : CascadeMux
    port map (
            O => \N__8948\,
            I => \N__8917\
        );

    \I__921\ : CascadeMux
    port map (
            O => \N__8947\,
            I => \N__8914\
        );

    \I__920\ : CascadeMux
    port map (
            O => \N__8946\,
            I => \N__8908\
        );

    \I__919\ : CascadeMux
    port map (
            O => \N__8945\,
            I => \N__8905\
        );

    \I__918\ : InMux
    port map (
            O => \N__8942\,
            I => \N__8899\
        );

    \I__917\ : InMux
    port map (
            O => \N__8941\,
            I => \N__8884\
        );

    \I__916\ : InMux
    port map (
            O => \N__8940\,
            I => \N__8884\
        );

    \I__915\ : InMux
    port map (
            O => \N__8939\,
            I => \N__8884\
        );

    \I__914\ : InMux
    port map (
            O => \N__8938\,
            I => \N__8884\
        );

    \I__913\ : InMux
    port map (
            O => \N__8935\,
            I => \N__8884\
        );

    \I__912\ : InMux
    port map (
            O => \N__8932\,
            I => \N__8884\
        );

    \I__911\ : InMux
    port map (
            O => \N__8929\,
            I => \N__8884\
        );

    \I__910\ : InMux
    port map (
            O => \N__8928\,
            I => \N__8881\
        );

    \I__909\ : InMux
    port map (
            O => \N__8927\,
            I => \N__8876\
        );

    \I__908\ : InMux
    port map (
            O => \N__8926\,
            I => \N__8876\
        );

    \I__907\ : InMux
    port map (
            O => \N__8923\,
            I => \N__8861\
        );

    \I__906\ : InMux
    port map (
            O => \N__8920\,
            I => \N__8861\
        );

    \I__905\ : InMux
    port map (
            O => \N__8917\,
            I => \N__8861\
        );

    \I__904\ : InMux
    port map (
            O => \N__8914\,
            I => \N__8861\
        );

    \I__903\ : InMux
    port map (
            O => \N__8913\,
            I => \N__8861\
        );

    \I__902\ : InMux
    port map (
            O => \N__8912\,
            I => \N__8861\
        );

    \I__901\ : InMux
    port map (
            O => \N__8911\,
            I => \N__8861\
        );

    \I__900\ : InMux
    port map (
            O => \N__8908\,
            I => \N__8850\
        );

    \I__899\ : InMux
    port map (
            O => \N__8905\,
            I => \N__8850\
        );

    \I__898\ : InMux
    port map (
            O => \N__8904\,
            I => \N__8850\
        );

    \I__897\ : InMux
    port map (
            O => \N__8903\,
            I => \N__8850\
        );

    \I__896\ : InMux
    port map (
            O => \N__8902\,
            I => \N__8850\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__8899\,
            I => \N__8847\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__8884\,
            I => \N__8840\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__8881\,
            I => \N__8840\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__8876\,
            I => \N__8840\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__8861\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__8850\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__889\ : Odrv4
    port map (
            O => \N__8847\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__888\ : Odrv4
    port map (
            O => \N__8840\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__887\ : InMux
    port map (
            O => \N__8831\,
            I => \N__8828\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__8828\,
            I => \N__8825\
        );

    \I__885\ : Span4Mux_v
    port map (
            O => \N__8825\,
            I => \N__8822\
        );

    \I__884\ : Odrv4
    port map (
            O => \N__8822\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2\
        );

    \I__883\ : CascadeMux
    port map (
            O => \N__8819\,
            I => \N__8813\
        );

    \I__882\ : CascadeMux
    port map (
            O => \N__8818\,
            I => \N__8807\
        );

    \I__881\ : CascadeMux
    port map (
            O => \N__8817\,
            I => \N__8804\
        );

    \I__880\ : CascadeMux
    port map (
            O => \N__8816\,
            I => \N__8801\
        );

    \I__879\ : InMux
    port map (
            O => \N__8813\,
            I => \N__8786\
        );

    \I__878\ : InMux
    port map (
            O => \N__8812\,
            I => \N__8781\
        );

    \I__877\ : InMux
    port map (
            O => \N__8811\,
            I => \N__8781\
        );

    \I__876\ : CascadeMux
    port map (
            O => \N__8810\,
            I => \N__8774\
        );

    \I__875\ : InMux
    port map (
            O => \N__8807\,
            I => \N__8766\
        );

    \I__874\ : InMux
    port map (
            O => \N__8804\,
            I => \N__8766\
        );

    \I__873\ : InMux
    port map (
            O => \N__8801\,
            I => \N__8766\
        );

    \I__872\ : InMux
    port map (
            O => \N__8800\,
            I => \N__8763\
        );

    \I__871\ : InMux
    port map (
            O => \N__8799\,
            I => \N__8746\
        );

    \I__870\ : InMux
    port map (
            O => \N__8798\,
            I => \N__8746\
        );

    \I__869\ : InMux
    port map (
            O => \N__8797\,
            I => \N__8746\
        );

    \I__868\ : InMux
    port map (
            O => \N__8796\,
            I => \N__8746\
        );

    \I__867\ : InMux
    port map (
            O => \N__8795\,
            I => \N__8746\
        );

    \I__866\ : InMux
    port map (
            O => \N__8794\,
            I => \N__8746\
        );

    \I__865\ : InMux
    port map (
            O => \N__8793\,
            I => \N__8746\
        );

    \I__864\ : InMux
    port map (
            O => \N__8792\,
            I => \N__8737\
        );

    \I__863\ : InMux
    port map (
            O => \N__8791\,
            I => \N__8737\
        );

    \I__862\ : InMux
    port map (
            O => \N__8790\,
            I => \N__8737\
        );

    \I__861\ : InMux
    port map (
            O => \N__8789\,
            I => \N__8737\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__8786\,
            I => \N__8734\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__8781\,
            I => \N__8731\
        );

    \I__858\ : InMux
    port map (
            O => \N__8780\,
            I => \N__8718\
        );

    \I__857\ : InMux
    port map (
            O => \N__8779\,
            I => \N__8718\
        );

    \I__856\ : InMux
    port map (
            O => \N__8778\,
            I => \N__8718\
        );

    \I__855\ : InMux
    port map (
            O => \N__8777\,
            I => \N__8718\
        );

    \I__854\ : InMux
    port map (
            O => \N__8774\,
            I => \N__8718\
        );

    \I__853\ : InMux
    port map (
            O => \N__8773\,
            I => \N__8718\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__8766\,
            I => \N__8713\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__8763\,
            I => \N__8713\
        );

    \I__850\ : InMux
    port map (
            O => \N__8762\,
            I => \N__8708\
        );

    \I__849\ : InMux
    port map (
            O => \N__8761\,
            I => \N__8708\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__8746\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__8737\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__846\ : Odrv4
    port map (
            O => \N__8734\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__845\ : Odrv4
    port map (
            O => \N__8731\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__8718\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__843\ : Odrv4
    port map (
            O => \N__8713\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__8708\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__841\ : CascadeMux
    port map (
            O => \N__8693\,
            I => \N__8690\
        );

    \I__840\ : InMux
    port map (
            O => \N__8690\,
            I => \N__8687\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__8687\,
            I => \phase_controller_slave.stoper_tr.N_60\
        );

    \I__838\ : InMux
    port map (
            O => \N__8684\,
            I => \N__8650\
        );

    \I__837\ : InMux
    port map (
            O => \N__8683\,
            I => \N__8650\
        );

    \I__836\ : InMux
    port map (
            O => \N__8682\,
            I => \N__8650\
        );

    \I__835\ : InMux
    port map (
            O => \N__8681\,
            I => \N__8650\
        );

    \I__834\ : InMux
    port map (
            O => \N__8680\,
            I => \N__8650\
        );

    \I__833\ : InMux
    port map (
            O => \N__8679\,
            I => \N__8650\
        );

    \I__832\ : InMux
    port map (
            O => \N__8678\,
            I => \N__8650\
        );

    \I__831\ : InMux
    port map (
            O => \N__8677\,
            I => \N__8633\
        );

    \I__830\ : InMux
    port map (
            O => \N__8676\,
            I => \N__8633\
        );

    \I__829\ : InMux
    port map (
            O => \N__8675\,
            I => \N__8633\
        );

    \I__828\ : InMux
    port map (
            O => \N__8674\,
            I => \N__8633\
        );

    \I__827\ : InMux
    port map (
            O => \N__8673\,
            I => \N__8633\
        );

    \I__826\ : InMux
    port map (
            O => \N__8672\,
            I => \N__8633\
        );

    \I__825\ : InMux
    port map (
            O => \N__8671\,
            I => \N__8633\
        );

    \I__824\ : InMux
    port map (
            O => \N__8670\,
            I => \N__8622\
        );

    \I__823\ : InMux
    port map (
            O => \N__8669\,
            I => \N__8622\
        );

    \I__822\ : InMux
    port map (
            O => \N__8668\,
            I => \N__8622\
        );

    \I__821\ : InMux
    port map (
            O => \N__8667\,
            I => \N__8622\
        );

    \I__820\ : InMux
    port map (
            O => \N__8666\,
            I => \N__8622\
        );

    \I__819\ : InMux
    port map (
            O => \N__8665\,
            I => \N__8617\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__8650\,
            I => \N__8614\
        );

    \I__817\ : InMux
    port map (
            O => \N__8649\,
            I => \N__8611\
        );

    \I__816\ : InMux
    port map (
            O => \N__8648\,
            I => \N__8608\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__8633\,
            I => \N__8603\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__8622\,
            I => \N__8603\
        );

    \I__813\ : InMux
    port map (
            O => \N__8621\,
            I => \N__8598\
        );

    \I__812\ : InMux
    port map (
            O => \N__8620\,
            I => \N__8598\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__8617\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__810\ : Odrv4
    port map (
            O => \N__8614\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__8611\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__8608\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__807\ : Odrv4
    port map (
            O => \N__8603\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__8598\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__805\ : InMux
    port map (
            O => \N__8585\,
            I => \N__8580\
        );

    \I__804\ : InMux
    port map (
            O => \N__8584\,
            I => \N__8577\
        );

    \I__803\ : InMux
    port map (
            O => \N__8583\,
            I => \N__8574\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__8580\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__8577\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__8574\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__799\ : CascadeMux
    port map (
            O => \N__8567\,
            I => \N__8564\
        );

    \I__798\ : InMux
    port map (
            O => \N__8564\,
            I => \N__8561\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__8561\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_1\
        );

    \I__796\ : InMux
    port map (
            O => \N__8558\,
            I => \N__8555\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__8555\,
            I => \N__8552\
        );

    \I__794\ : Span4Mux_s3_h
    port map (
            O => \N__8552\,
            I => \N__8548\
        );

    \I__793\ : InMux
    port map (
            O => \N__8551\,
            I => \N__8545\
        );

    \I__792\ : Odrv4
    port map (
            O => \N__8548\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__8545\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__790\ : CascadeMux
    port map (
            O => \N__8540\,
            I => \N__8537\
        );

    \I__789\ : InMux
    port map (
            O => \N__8537\,
            I => \N__8534\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__8534\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_2\
        );

    \I__787\ : InMux
    port map (
            O => \N__8531\,
            I => \N__8527\
        );

    \I__786\ : InMux
    port map (
            O => \N__8530\,
            I => \N__8524\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__8527\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__8524\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__783\ : CascadeMux
    port map (
            O => \N__8519\,
            I => \N__8516\
        );

    \I__782\ : InMux
    port map (
            O => \N__8516\,
            I => \N__8513\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__8513\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_3\
        );

    \I__780\ : CascadeMux
    port map (
            O => \N__8510\,
            I => \N__8507\
        );

    \I__779\ : InMux
    port map (
            O => \N__8507\,
            I => \N__8504\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__8504\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\
        );

    \I__777\ : CascadeMux
    port map (
            O => \N__8501\,
            I => \N__8498\
        );

    \I__776\ : InMux
    port map (
            O => \N__8498\,
            I => \N__8495\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__8495\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIUSZ0Z53\
        );

    \I__774\ : CascadeMux
    port map (
            O => \N__8492\,
            I => \N__8489\
        );

    \I__773\ : InMux
    port map (
            O => \N__8489\,
            I => \N__8486\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__8486\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10\
        );

    \I__771\ : InMux
    port map (
            O => \N__8483\,
            I => \N__8480\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__8480\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11\
        );

    \I__769\ : InMux
    port map (
            O => \N__8477\,
            I => \N__8474\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__8474\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13\
        );

    \I__767\ : InMux
    port map (
            O => \N__8471\,
            I => \N__8468\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__8468\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14\
        );

    \I__765\ : InMux
    port map (
            O => \N__8465\,
            I => \N__8462\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__8462\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15\
        );

    \I__763\ : InMux
    port map (
            O => \N__8459\,
            I => \N__8456\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__8456\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16\
        );

    \I__761\ : InMux
    port map (
            O => \N__8453\,
            I => \N__8450\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__8450\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17\
        );

    \I__759\ : InMux
    port map (
            O => \N__8447\,
            I => \N__8444\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__8444\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4\
        );

    \I__757\ : CascadeMux
    port map (
            O => \N__8441\,
            I => \N__8438\
        );

    \I__756\ : InMux
    port map (
            O => \N__8438\,
            I => \N__8435\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__8435\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5\
        );

    \I__754\ : InMux
    port map (
            O => \N__8432\,
            I => \N__8429\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__8429\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6\
        );

    \I__752\ : CascadeMux
    port map (
            O => \N__8426\,
            I => \N__8423\
        );

    \I__751\ : InMux
    port map (
            O => \N__8423\,
            I => \N__8420\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__8420\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7\
        );

    \I__749\ : InMux
    port map (
            O => \N__8417\,
            I => \N__8414\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__8414\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8\
        );

    \I__747\ : CascadeMux
    port map (
            O => \N__8411\,
            I => \N__8408\
        );

    \I__746\ : InMux
    port map (
            O => \N__8408\,
            I => \N__8405\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__8405\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9\
        );

    \I__744\ : CascadeMux
    port map (
            O => \N__8402\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\
        );

    \I__743\ : InMux
    port map (
            O => \N__8399\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16\
        );

    \I__742\ : InMux
    port map (
            O => \N__8396\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17\
        );

    \I__741\ : InMux
    port map (
            O => \N__8393\,
            I => \N__8390\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__8390\,
            I => \N_39_i_i\
        );

    \I__739\ : InMux
    port map (
            O => \N__8387\,
            I => \N__8384\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__8384\,
            I => \N__8381\
        );

    \I__737\ : Span12Mux_s3_v
    port map (
            O => \N__8381\,
            I => \N__8378\
        );

    \I__736\ : Span12Mux_h
    port map (
            O => \N__8378\,
            I => \N__8375\
        );

    \I__735\ : Span12Mux_h
    port map (
            O => \N__8375\,
            I => \N__8369\
        );

    \I__734\ : InMux
    port map (
            O => \N__8374\,
            I => \N__8366\
        );

    \I__733\ : InMux
    port map (
            O => \N__8373\,
            I => \N__8363\
        );

    \I__732\ : InMux
    port map (
            O => \N__8372\,
            I => \N__8360\
        );

    \I__731\ : Odrv12
    port map (
            O => \N__8369\,
            I => \CONSTANT_ONE_NET\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__8366\,
            I => \CONSTANT_ONE_NET\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__8363\,
            I => \CONSTANT_ONE_NET\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__8360\,
            I => \CONSTANT_ONE_NET\
        );

    \I__727\ : InMux
    port map (
            O => \N__8351\,
            I => \N__8348\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__8348\,
            I => \rgb_drv_RNOZ0\
        );

    \I__725\ : InMux
    port map (
            O => \N__8345\,
            I => \N__8342\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__8342\,
            I => \N__8339\
        );

    \I__723\ : Odrv4
    port map (
            O => \N__8339\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12\
        );

    \I__722\ : CascadeMux
    port map (
            O => \N__8336\,
            I => \N__8333\
        );

    \I__721\ : InMux
    port map (
            O => \N__8333\,
            I => \N__8330\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__8330\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3\
        );

    \I__719\ : InMux
    port map (
            O => \N__8327\,
            I => \bfn_1_19_0_\
        );

    \I__718\ : InMux
    port map (
            O => \N__8324\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8\
        );

    \I__717\ : InMux
    port map (
            O => \N__8321\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9\
        );

    \I__716\ : InMux
    port map (
            O => \N__8318\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10\
        );

    \I__715\ : InMux
    port map (
            O => \N__8315\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11\
        );

    \I__714\ : InMux
    port map (
            O => \N__8312\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12\
        );

    \I__713\ : InMux
    port map (
            O => \N__8309\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13\
        );

    \I__712\ : InMux
    port map (
            O => \N__8306\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14\
        );

    \I__711\ : InMux
    port map (
            O => \N__8303\,
            I => \bfn_1_20_0_\
        );

    \I__710\ : InMux
    port map (
            O => \N__8300\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0\
        );

    \I__709\ : InMux
    port map (
            O => \N__8297\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1\
        );

    \I__708\ : InMux
    port map (
            O => \N__8294\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2\
        );

    \I__707\ : InMux
    port map (
            O => \N__8291\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3\
        );

    \I__706\ : InMux
    port map (
            O => \N__8288\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4\
        );

    \I__705\ : InMux
    port map (
            O => \N__8285\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5\
        );

    \I__704\ : InMux
    port map (
            O => \N__8282\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6\
        );

    \IN_MUX_bfv_1_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_18_0_\
        );

    \IN_MUX_bfv_1_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_1_19_0_\
        );

    \IN_MUX_bfv_1_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_1_20_0_\
        );

    \IN_MUX_bfv_7_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_17_0_\
        );

    \IN_MUX_bfv_7_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_7_18_0_\
        );

    \IN_MUX_bfv_7_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_7_19_0_\
        );

    \IN_MUX_bfv_8_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_25_0_\
        );

    \IN_MUX_bfv_8_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_8_26_0_\
        );

    \IN_MUX_bfv_8_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_8_27_0_\
        );

    \IN_MUX_bfv_12_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_15_0_\
        );

    \IN_MUX_bfv_12_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_12_16_0_\
        );

    \IN_MUX_bfv_12_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_12_17_0_\
        );

    \IN_MUX_bfv_3_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_18_0_\
        );

    \IN_MUX_bfv_3_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8\,
            carryinitout => \bfn_3_19_0_\
        );

    \IN_MUX_bfv_3_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16\,
            carryinitout => \bfn_3_20_0_\
        );

    \IN_MUX_bfv_9_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_17_0_\
        );

    \IN_MUX_bfv_9_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8\,
            carryinitout => \bfn_9_18_0_\
        );

    \IN_MUX_bfv_9_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16\,
            carryinitout => \bfn_9_19_0_\
        );

    \IN_MUX_bfv_7_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_23_0_\
        );

    \IN_MUX_bfv_7_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            carryinitout => \bfn_7_24_0_\
        );

    \IN_MUX_bfv_7_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            carryinitout => \bfn_7_25_0_\
        );

    \IN_MUX_bfv_10_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_15_0_\
        );

    \IN_MUX_bfv_10_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            carryinitout => \bfn_10_16_0_\
        );

    \IN_MUX_bfv_10_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            carryinitout => \bfn_10_17_0_\
        );

    \IN_MUX_bfv_13_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_19_0_\
        );

    \IN_MUX_bfv_13_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_13_20_0_\
        );

    \IN_MUX_bfv_13_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_13_21_0_\
        );

    \IN_MUX_bfv_13_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_13_22_0_\
        );

    \IN_MUX_bfv_12_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_18_0_\
        );

    \IN_MUX_bfv_12_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            carryinitout => \bfn_12_19_0_\
        );

    \IN_MUX_bfv_12_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            carryinitout => \bfn_12_20_0_\
        );

    \IN_MUX_bfv_12_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            carryinitout => \bfn_12_21_0_\
        );

    \IN_MUX_bfv_8_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_13_0_\
        );

    \IN_MUX_bfv_8_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_8_14_0_\
        );

    \IN_MUX_bfv_8_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_8_15_0_\
        );

    \IN_MUX_bfv_8_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_8_16_0_\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_7_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            carryinitout => \bfn_7_14_0_\
        );

    \IN_MUX_bfv_7_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            carryinitout => \bfn_7_15_0_\
        );

    \IN_MUX_bfv_7_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            carryinitout => \bfn_7_16_0_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQOU9A_0_31\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__14045\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.N_32_g\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__12431\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.delay_tr_timer.N_180_i_g\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__18785\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.delay_hc_timer.N_178_i_g\
        );

    \osc\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b10"
        )
    port map (
            CLKHFPU => \N__8372\,
            CLKHFEN => \N__8374\,
            CLKHF => clk_12mhz
        );

    \rgb_drv\ : SB_RGBA_DRV
    generic map (
            RGB2_CURRENT => "0b111111",
            CURRENT_MODE => "0b0",
            RGB0_CURRENT => "0b111111",
            RGB1_CURRENT => "0b111111"
        )
    port map (
            RGBLEDEN => \N__8373\,
            RGB2PWM => \N__8393\,
            RGB1 => rgb_g_wire,
            CURREN => \N__8387\,
            RGB2 => rgb_b_wire,
            RGB1PWM => \N__8351\,
            RGB0PWM => \N__20902\,
            RGB0 => rgb_r_wire
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__15449\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.delay_tr_timer.N_181_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_1_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8584\,
            in2 => \N__8510\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_18_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_1_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8558\,
            in2 => \_gnd_net_\,
            in3 => \N__8300\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_1_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8531\,
            in2 => \N__8501\,
            in3 => \N__8297\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_1_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9143\,
            in2 => \_gnd_net_\,
            in3 => \N__8294\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_1_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9122\,
            in2 => \_gnd_net_\,
            in3 => \N__8291\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_1_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9098\,
            in3 => \N__8288\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_1_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9074\,
            in2 => \_gnd_net_\,
            in3 => \N__8285\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_1_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9053\,
            in3 => \N__8282\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_1_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9029\,
            in2 => \_gnd_net_\,
            in3 => \N__8327\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9\,
            ltout => OPEN,
            carryin => \bfn_1_19_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_1_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9008\,
            in2 => \_gnd_net_\,
            in3 => \N__8324\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_1_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8987\,
            in2 => \_gnd_net_\,
            in3 => \N__8321\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_1_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9323\,
            in2 => \_gnd_net_\,
            in3 => \N__8318\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_1_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9290\,
            in2 => \_gnd_net_\,
            in3 => \N__8315\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_1_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9269\,
            in2 => \_gnd_net_\,
            in3 => \N__8312\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_1_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9248\,
            in2 => \_gnd_net_\,
            in3 => \N__8309\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_1_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9227\,
            in2 => \_gnd_net_\,
            in3 => \N__8306\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_1_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9206\,
            in2 => \_gnd_net_\,
            in3 => \N__8303\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17\,
            ltout => OPEN,
            carryin => \bfn_1_20_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_1_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9185\,
            in2 => \_gnd_net_\,
            in3 => \N__8399\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_1_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9164\,
            in2 => \_gnd_net_\,
            in3 => \N__8396\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_drv_RNO_0_LC_1_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__21571\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20900\,
            lcout => \N_39_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_1_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_drv_RNO_LC_1_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__20901\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21575\,
            lcout => \rgb_drv_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_12_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__8649\,
            in1 => \N__8928\,
            in2 => \N__8819\,
            in3 => \N__8345\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21189\,
            ce => 'H',
            sr => \N__20820\
        );

    \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8927\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8621\,
            lcout => \phase_controller_slave.stoper_tr.N_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.stoper_state_RNII60D_1_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__8926\,
            in1 => \N__8620\,
            in2 => \_gnd_net_\,
            in3 => \N__8800\,
            lcout => \phase_controller_slave.stoper_tr.stoper_state_RNII60DZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_3_LC_2_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__8678\,
            in1 => \N__8938\,
            in2 => \N__8336\,
            in3 => \N__8796\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21178\,
            ce => 'H',
            sr => \N__20831\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_4_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__8793\,
            in1 => \N__8682\,
            in2 => \N__8951\,
            in3 => \N__8447\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21178\,
            ce => 'H',
            sr => \N__20831\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_5_LC_2_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__8679\,
            in1 => \N__8939\,
            in2 => \N__8441\,
            in3 => \N__8797\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21178\,
            ce => 'H',
            sr => \N__20831\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_6_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__8794\,
            in1 => \N__8683\,
            in2 => \N__8952\,
            in3 => \N__8432\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21178\,
            ce => 'H',
            sr => \N__20831\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_7_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__8680\,
            in1 => \N__8940\,
            in2 => \N__8426\,
            in3 => \N__8798\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21178\,
            ce => 'H',
            sr => \N__20831\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_8_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__8795\,
            in1 => \N__8684\,
            in2 => \N__8953\,
            in3 => \N__8417\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21178\,
            ce => 'H',
            sr => \N__20831\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_9_LC_2_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__8681\,
            in1 => \N__8941\,
            in2 => \N__8411\,
            in3 => \N__8799\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21178\,
            ce => 'H',
            sr => \N__20831\
        );

    \phase_controller_slave.stoper_tr.stoper_state_0_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__9417\,
            in1 => \N__8669\,
            in2 => \N__8945\,
            in3 => \N__8779\,
            lcout => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21173\,
            ce => 'H',
            sr => \N__20837\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_2_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__8773\,
            in1 => \N__8585\,
            in2 => \_gnd_net_\,
            in3 => \N__9416\,
            lcout => OPEN,
            ltout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_1_LC_2_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__8903\,
            in1 => \N__8668\,
            in2 => \N__8402\,
            in3 => \N__8778\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21173\,
            ce => 'H',
            sr => \N__20837\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_2_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8761\,
            in2 => \_gnd_net_\,
            in3 => \N__9414\,
            lcout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.stoper_state_1_LC_2_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010111000000"
        )
    port map (
            in0 => \N__9418\,
            in1 => \N__8670\,
            in2 => \N__8946\,
            in3 => \N__8780\,
            lcout => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21173\,
            ce => 'H',
            sr => \N__20837\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIUS53_LC_2_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8762\,
            in2 => \_gnd_net_\,
            in3 => \N__9415\,
            lcout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIUSZ0Z53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_10_LC_2_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__8902\,
            in1 => \N__8667\,
            in2 => \N__8492\,
            in3 => \N__8777\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21173\,
            ce => 'H',
            sr => \N__20837\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_11_LC_2_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__8666\,
            in1 => \N__8904\,
            in2 => \N__8810\,
            in3 => \N__8483\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21173\,
            ce => 'H',
            sr => \N__20837\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_13_LC_2_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__8789\,
            in1 => \N__8674\,
            in2 => \N__8947\,
            in3 => \N__8477\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21163\,
            ce => 'H',
            sr => \N__20839\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_14_LC_2_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__8671\,
            in1 => \N__8911\,
            in2 => \N__8816\,
            in3 => \N__8471\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21163\,
            ce => 'H',
            sr => \N__20839\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_15_LC_2_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__8790\,
            in1 => \N__8675\,
            in2 => \N__8948\,
            in3 => \N__8465\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21163\,
            ce => 'H',
            sr => \N__20839\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_16_LC_2_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__8672\,
            in1 => \N__8912\,
            in2 => \N__8817\,
            in3 => \N__8459\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21163\,
            ce => 'H',
            sr => \N__20839\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_17_LC_2_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__8791\,
            in1 => \N__8676\,
            in2 => \N__8949\,
            in3 => \N__8453\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21163\,
            ce => 'H',
            sr => \N__20839\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_18_LC_2_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__8673\,
            in1 => \N__8913\,
            in2 => \N__8818\,
            in3 => \N__8966\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21163\,
            ce => 'H',
            sr => \N__20839\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_19_LC_2_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__8792\,
            in1 => \N__8677\,
            in2 => \N__8950\,
            in3 => \N__8960\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21163\,
            ce => 'H',
            sr => \N__20839\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_2_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__8648\,
            in1 => \N__8811\,
            in2 => \N__8954\,
            in3 => \N__8831\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21179\,
            ce => 'H',
            sr => \N__20821\
        );

    \phase_controller_slave.stoper_tr.time_passed_LC_3_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__9391\,
            in1 => \N__8812\,
            in2 => \N__8693\,
            in3 => \N__9422\,
            lcout => \phase_controller_slave.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21179\,
            ce => 'H',
            sr => \N__20821\
        );

    \phase_controller_slave.start_timer_tr_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101110"
        )
    port map (
            in0 => \N__9362\,
            in1 => \N__8665\,
            in2 => \N__9827\,
            in3 => \N__9838\,
            lcout => \phase_controller_slave.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21179\,
            ce => 'H',
            sr => \N__20821\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9344\,
            in2 => \N__8567\,
            in3 => \N__8583\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_3_18_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__8551\,
            in1 => \N__9503\,
            in2 => \N__8540\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__8530\,
            in1 => \N__9350\,
            in2 => \N__8519\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_3_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9329\,
            in2 => \N__9131\,
            in3 => \N__9142\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_3_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9485\,
            in2 => \N__9107\,
            in3 => \N__9118\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_3_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9476\,
            in2 => \N__9083\,
            in3 => \N__9094\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_3_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9356\,
            in2 => \N__9062\,
            in3 => \N__9073\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_3_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9338\,
            in2 => \N__9038\,
            in3 => \N__9049\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9449\,
            in2 => \N__9017\,
            in3 => \N__9028\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_3_19_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_3_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9608\,
            in2 => \N__8996\,
            in3 => \N__9007\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9614\,
            in2 => \N__8975\,
            in3 => \N__8986\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9599\,
            in2 => \N__9299\,
            in3 => \N__9322\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_3_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9289\,
            in1 => \N__9494\,
            in2 => \N__9278\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_3_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9464\,
            in2 => \N__9257\,
            in3 => \N__9268\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9455\,
            in2 => \N__9236\,
            in3 => \N__9247\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_3_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9623\,
            in2 => \N__9215\,
            in3 => \N__9226\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_3_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9437\,
            in2 => \N__9194\,
            in3 => \N__9205\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_3_20_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_3_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9431\,
            in2 => \N__9173\,
            in3 => \N__9184\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_3_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9593\,
            in2 => \N__9152\,
            in3 => \N__9163\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_3_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9425\,
            lcout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.state_0_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000111110001000"
        )
    port map (
            in0 => \N__9751\,
            in1 => \N__9686\,
            in2 => \N__9395\,
            in3 => \N__9374\,
            lcout => \phase_controller_slave.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21180\,
            ce => 'H',
            sr => \N__20813\
        );

    \phase_controller_slave.state_RNIVDE2_0_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9390\,
            in2 => \_gnd_net_\,
            in3 => \N__9373\,
            lcout => \phase_controller_slave.state_RNIVDE2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.start_timer_tr_RNO_0_LC_4_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9749\,
            in2 => \_gnd_net_\,
            in3 => \N__9684\,
            lcout => \phase_controller_slave.start_timer_tr_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.target_time_7_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010000010100000"
        )
    port map (
            in0 => \N__11874\,
            in1 => \N__11614\,
            in2 => \N__13805\,
            in3 => \N__11770\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21164\,
            ce => \N__9575\,
            sr => \N__20822\
        );

    \phase_controller_slave.stoper_tr.target_time_3_LC_4_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100110000000000"
        )
    port map (
            in0 => \N__11612\,
            in1 => \N__15113\,
            in2 => \N__11785\,
            in3 => \N__11877\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21164\,
            ce => \N__9575\,
            sr => \N__20822\
        );

    \phase_controller_slave.stoper_tr.target_time_1_LC_4_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010000010100000"
        )
    port map (
            in0 => \N__11873\,
            in1 => \N__11611\,
            in2 => \N__13544\,
            in3 => \N__11763\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21164\,
            ce => \N__9575\,
            sr => \N__20822\
        );

    \phase_controller_slave.stoper_tr.target_time_8_LC_4_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100110000000000"
        )
    port map (
            in0 => \N__11615\,
            in1 => \N__11876\,
            in2 => \N__11787\,
            in3 => \N__12630\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21164\,
            ce => \N__9575\,
            sr => \N__20822\
        );

    \phase_controller_slave.stoper_tr.target_time_4_LC_4_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100110000000000"
        )
    port map (
            in0 => \N__11613\,
            in1 => \N__11875\,
            in2 => \N__11786\,
            in3 => \N__15032\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21164\,
            ce => \N__9575\,
            sr => \N__20822\
        );

    \phase_controller_slave.stoper_tr.target_time_2_LC_4_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011101010"
        )
    port map (
            in0 => \N__14918\,
            in1 => \N__11202\,
            in2 => \N__11240\,
            in3 => \N__10159\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21157\,
            ce => \N__9583\,
            sr => \N__20827\
        );

    \phase_controller_slave.stoper_tr.target_time_13_LC_4_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__11610\,
            in1 => \N__11761\,
            in2 => \N__11900\,
            in3 => \N__14806\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21157\,
            ce => \N__9583\,
            sr => \N__20827\
        );

    \phase_controller_slave.stoper_tr.target_time_5_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011101100"
        )
    port map (
            in0 => \N__11239\,
            in1 => \N__13430\,
            in2 => \N__11207\,
            in3 => \N__10160\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21157\,
            ce => \N__9583\,
            sr => \N__20827\
        );

    \phase_controller_slave.stoper_tr.target_timeZ0Z_6_LC_4_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111101110111011"
        )
    port map (
            in0 => \N__13649\,
            in1 => \N__11893\,
            in2 => \N__11784\,
            in3 => \N__11609\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21157\,
            ce => \N__9583\,
            sr => \N__20827\
        );

    \phase_controller_slave.stoper_tr.target_time_14_LC_4_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__11762\,
            in1 => \N__13580\,
            in2 => \_gnd_net_\,
            in3 => \N__13727\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21157\,
            ce => \N__9583\,
            sr => \N__20827\
        );

    \phase_controller_slave.stoper_tr.target_time_15_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13718\,
            in2 => \_gnd_net_\,
            in3 => \N__11750\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21151\,
            ce => \N__9582\,
            sr => \N__20832\
        );

    \phase_controller_slave.stoper_tr.target_time_9_LC_4_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001000"
        )
    port map (
            in0 => \N__11582\,
            in1 => \N__11781\,
            in2 => \N__13726\,
            in3 => \N__13468\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21151\,
            ce => \N__9582\,
            sr => \N__20832\
        );

    \phase_controller_slave.stoper_tr.target_time_17_LC_4_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13508\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21151\,
            ce => \N__9582\,
            sr => \N__20832\
        );

    \phase_controller_slave.stoper_tr.target_time_18_LC_4_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15066\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21151\,
            ce => \N__9582\,
            sr => \N__20832\
        );

    \phase_controller_slave.stoper_tr.target_time_16_LC_4_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13760\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21151\,
            ce => \N__9582\,
            sr => \N__20832\
        );

    \phase_controller_slave.stoper_tr.target_time_11_LC_4_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100110000000000"
        )
    port map (
            in0 => \N__11580\,
            in1 => \N__14842\,
            in2 => \N__11782\,
            in3 => \N__11898\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21151\,
            ce => \N__9582\,
            sr => \N__20832\
        );

    \phase_controller_slave.stoper_tr.target_time_10_LC_4_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010000010100000"
        )
    port map (
            in0 => \N__11897\,
            in1 => \N__11751\,
            in2 => \N__14882\,
            in3 => \N__11579\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21151\,
            ce => \N__9582\,
            sr => \N__20832\
        );

    \phase_controller_slave.stoper_tr.target_time_12_LC_4_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100110000000000"
        )
    port map (
            in0 => \N__11581\,
            in1 => \N__13612\,
            in2 => \N__11783\,
            in3 => \N__11899\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21151\,
            ce => \N__9582\,
            sr => \N__20832\
        );

    \phase_controller_slave.stoper_tr.target_time_19_LC_4_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16933\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21145\,
            ce => \N__9587\,
            sr => \N__20838\
        );

    \phase_controller_inst1.stoper_tr.target_time_19_LC_4_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16934\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21138\,
            ce => \N__12035\,
            sr => \N__20843\
        );

    \SB_DFF_inst_PH2_MAX_D1_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9539\,
            lcout => \il_max_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21194\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MIN_D1_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9527\,
            lcout => \il_min_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21192\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MIN_D2_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9509\,
            lcout => \il_min_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21192\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MAX_D2_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9710\,
            lcout => \il_max_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21190\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.start_timer_hc_RNO_1_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13923\,
            in2 => \_gnd_net_\,
            in3 => \N__9636\,
            lcout => \phase_controller_slave.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.start_timer_hc_RNO_0_LC_5_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9657\,
            in2 => \_gnd_net_\,
            in3 => \N__9864\,
            lcout => \phase_controller_slave.start_timer_hc_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.start_timer_hc_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101110101010"
        )
    port map (
            in0 => \N__9701\,
            in1 => \N__9692\,
            in2 => \N__9823\,
            in3 => \N__11428\,
            lcout => \phase_controller_slave.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21165\,
            ce => 'H',
            sr => \N__20814\
        );

    \phase_controller_slave.state_1_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__9866\,
            in1 => \N__9750\,
            in2 => \N__9662\,
            in3 => \N__9685\,
            lcout => \phase_controller_slave.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21165\,
            ce => 'H',
            sr => \N__20814\
        );

    \phase_controller_slave.state_2_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__9644\,
            in1 => \N__9658\,
            in2 => \N__13930\,
            in3 => \N__9865\,
            lcout => \phase_controller_slave.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21165\,
            ce => 'H',
            sr => \N__20814\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_12_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__11427\,
            in1 => \N__11360\,
            in2 => \N__13289\,
            in3 => \N__10001\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21158\,
            ce => 'H',
            sr => \N__20819\
        );

    \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_5_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11426\,
            in2 => \_gnd_net_\,
            in3 => \N__11359\,
            lcout => \phase_controller_slave.stoper_hc.N_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.state_3_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000010101100"
        )
    port map (
            in0 => \N__9785\,
            in1 => \N__13916\,
            in2 => \N__9822\,
            in3 => \N__9643\,
            lcout => \phase_controller_slave.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21152\,
            ce => 'H',
            sr => \N__20823\
        );

    \phase_controller_slave.stoper_hc.time_passed_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__9863\,
            in1 => \N__13288\,
            in2 => \N__9875\,
            in3 => \N__13145\,
            lcout => \phase_controller_slave.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21152\,
            ce => 'H',
            sr => \N__20823\
        );

    \phase_controller_slave.state_4_LC_5_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100111011101110"
        )
    port map (
            in0 => \N__9812\,
            in1 => \N__9842\,
            in2 => \N__21555\,
            in3 => \N__9779\,
            lcout => \phase_controller_slave.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21152\,
            ce => 'H',
            sr => \N__20823\
        );

    \phase_controller_slave.state_RNO_0_3_LC_5_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21556\,
            in2 => \_gnd_net_\,
            in3 => \N__9771\,
            lcout => \phase_controller_slave.state_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.T01_LC_5_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__21487\,
            in1 => \N__19505\,
            in2 => \N__9778\,
            in3 => \N__15215\,
            lcout => shift_flag_start,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21142\,
            ce => 'H',
            sr => \N__20833\
        );

    \phase_controller_slave.S2_LC_5_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9755\,
            lcout => s4_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21142\,
            ce => 'H',
            sr => \N__20833\
        );

    \phase_controller_inst1.stoper_tr.target_time_10_LC_5_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100010001000"
        )
    port map (
            in0 => \N__11890\,
            in1 => \N__14881\,
            in2 => \N__11788\,
            in3 => \N__11616\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21128\,
            ce => \N__12029\,
            sr => \N__20844\
        );

    \phase_controller_inst1.stoper_tr.target_time_11_LC_5_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__11617\,
            in1 => \N__11777\,
            in2 => \N__14849\,
            in3 => \N__11891\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21128\,
            ce => \N__12029\,
            sr => \N__20844\
        );

    \phase_controller_inst1.stoper_tr.target_time_9_LC_5_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110011101100"
        )
    port map (
            in0 => \N__13725\,
            in1 => \N__13472\,
            in2 => \N__11789\,
            in3 => \N__11618\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21128\,
            ce => \N__12029\,
            sr => \N__20844\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10490\,
            lcout => \delay_measurement_inst.elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21186\,
            ce => \N__10889\,
            sr => \N__20783\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10472\,
            lcout => \delay_measurement_inst.elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21186\,
            ce => \N__10889\,
            sr => \N__20783\
        );

    \delay_measurement_inst.delay_hc_timer.counter_0_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17636\,
            in1 => \N__10488\,
            in2 => \_gnd_net_\,
            in3 => \N__9902\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_7_13_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            clk => \N__21181\,
            ce => \N__17498\,
            sr => \N__20788\
        );

    \delay_measurement_inst.delay_hc_timer.counter_1_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17536\,
            in1 => \N__10470\,
            in2 => \_gnd_net_\,
            in3 => \N__9899\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            clk => \N__21181\,
            ce => \N__17498\,
            sr => \N__20788\
        );

    \delay_measurement_inst.delay_hc_timer.counter_2_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17637\,
            in1 => \N__10449\,
            in2 => \_gnd_net_\,
            in3 => \N__9896\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            clk => \N__21181\,
            ce => \N__17498\,
            sr => \N__20788\
        );

    \delay_measurement_inst.delay_hc_timer.counter_3_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17537\,
            in1 => \N__10425\,
            in2 => \_gnd_net_\,
            in3 => \N__9893\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            clk => \N__21181\,
            ce => \N__17498\,
            sr => \N__20788\
        );

    \delay_measurement_inst.delay_hc_timer.counter_4_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17638\,
            in1 => \N__10403\,
            in2 => \_gnd_net_\,
            in3 => \N__9890\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            clk => \N__21181\,
            ce => \N__17498\,
            sr => \N__20788\
        );

    \delay_measurement_inst.delay_hc_timer.counter_5_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17538\,
            in1 => \N__10667\,
            in2 => \_gnd_net_\,
            in3 => \N__9887\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            clk => \N__21181\,
            ce => \N__17498\,
            sr => \N__20788\
        );

    \delay_measurement_inst.delay_hc_timer.counter_6_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17639\,
            in1 => \N__10647\,
            in2 => \_gnd_net_\,
            in3 => \N__9884\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            clk => \N__21181\,
            ce => \N__17498\,
            sr => \N__20788\
        );

    \delay_measurement_inst.delay_hc_timer.counter_7_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17539\,
            in1 => \N__10623\,
            in2 => \_gnd_net_\,
            in3 => \N__9881\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            clk => \N__21181\,
            ce => \N__17498\,
            sr => \N__20788\
        );

    \delay_measurement_inst.delay_hc_timer.counter_8_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17573\,
            in1 => \N__10600\,
            in2 => \_gnd_net_\,
            in3 => \N__9878\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_7_14_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            clk => \N__21174\,
            ce => \N__17500\,
            sr => \N__20793\
        );

    \delay_measurement_inst.delay_hc_timer.counter_9_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17577\,
            in1 => \N__10579\,
            in2 => \_gnd_net_\,
            in3 => \N__9929\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            clk => \N__21174\,
            ce => \N__17500\,
            sr => \N__20793\
        );

    \delay_measurement_inst.delay_hc_timer.counter_10_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17570\,
            in1 => \N__10557\,
            in2 => \_gnd_net_\,
            in3 => \N__9926\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            clk => \N__21174\,
            ce => \N__17500\,
            sr => \N__20793\
        );

    \delay_measurement_inst.delay_hc_timer.counter_11_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17574\,
            in1 => \N__10533\,
            in2 => \_gnd_net_\,
            in3 => \N__9923\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            clk => \N__21174\,
            ce => \N__17500\,
            sr => \N__20793\
        );

    \delay_measurement_inst.delay_hc_timer.counter_12_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17571\,
            in1 => \N__10511\,
            in2 => \_gnd_net_\,
            in3 => \N__9920\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            clk => \N__21174\,
            ce => \N__17500\,
            sr => \N__20793\
        );

    \delay_measurement_inst.delay_hc_timer.counter_13_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17575\,
            in1 => \N__10859\,
            in2 => \_gnd_net_\,
            in3 => \N__9917\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            clk => \N__21174\,
            ce => \N__17500\,
            sr => \N__20793\
        );

    \delay_measurement_inst.delay_hc_timer.counter_14_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17572\,
            in1 => \N__10839\,
            in2 => \_gnd_net_\,
            in3 => \N__9914\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            clk => \N__21174\,
            ce => \N__17500\,
            sr => \N__20793\
        );

    \delay_measurement_inst.delay_hc_timer.counter_15_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17576\,
            in1 => \N__10815\,
            in2 => \_gnd_net_\,
            in3 => \N__9911\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            clk => \N__21174\,
            ce => \N__17500\,
            sr => \N__20793\
        );

    \delay_measurement_inst.delay_hc_timer.counter_16_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17617\,
            in1 => \N__10792\,
            in2 => \_gnd_net_\,
            in3 => \N__9908\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_7_15_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            clk => \N__21166\,
            ce => \N__17499\,
            sr => \N__20800\
        );

    \delay_measurement_inst.delay_hc_timer.counter_17_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17587\,
            in1 => \N__10771\,
            in2 => \_gnd_net_\,
            in3 => \N__9905\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            clk => \N__21166\,
            ce => \N__17499\,
            sr => \N__20800\
        );

    \delay_measurement_inst.delay_hc_timer.counter_18_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17618\,
            in1 => \N__10749\,
            in2 => \_gnd_net_\,
            in3 => \N__9956\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            clk => \N__21166\,
            ce => \N__17499\,
            sr => \N__20800\
        );

    \delay_measurement_inst.delay_hc_timer.counter_19_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17588\,
            in1 => \N__10725\,
            in2 => \_gnd_net_\,
            in3 => \N__9953\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            clk => \N__21166\,
            ce => \N__17499\,
            sr => \N__20800\
        );

    \delay_measurement_inst.delay_hc_timer.counter_20_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17619\,
            in1 => \N__10703\,
            in2 => \_gnd_net_\,
            in3 => \N__9950\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            clk => \N__21166\,
            ce => \N__17499\,
            sr => \N__20800\
        );

    \delay_measurement_inst.delay_hc_timer.counter_21_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17589\,
            in1 => \N__10685\,
            in2 => \_gnd_net_\,
            in3 => \N__9947\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            clk => \N__21166\,
            ce => \N__17499\,
            sr => \N__20800\
        );

    \delay_measurement_inst.delay_hc_timer.counter_22_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17620\,
            in1 => \N__11052\,
            in2 => \_gnd_net_\,
            in3 => \N__9944\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            clk => \N__21166\,
            ce => \N__17499\,
            sr => \N__20800\
        );

    \delay_measurement_inst.delay_hc_timer.counter_23_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17590\,
            in1 => \N__11028\,
            in2 => \_gnd_net_\,
            in3 => \N__9941\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            clk => \N__21166\,
            ce => \N__17499\,
            sr => \N__20800\
        );

    \delay_measurement_inst.delay_hc_timer.counter_24_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17621\,
            in1 => \N__11005\,
            in2 => \_gnd_net_\,
            in3 => \N__9938\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_7_16_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            clk => \N__21159\,
            ce => \N__17501\,
            sr => \N__20805\
        );

    \delay_measurement_inst.delay_hc_timer.counter_25_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17625\,
            in1 => \N__10984\,
            in2 => \_gnd_net_\,
            in3 => \N__9935\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            clk => \N__21159\,
            ce => \N__17501\,
            sr => \N__20805\
        );

    \delay_measurement_inst.delay_hc_timer.counter_26_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17622\,
            in1 => \N__10950\,
            in2 => \_gnd_net_\,
            in3 => \N__9932\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            clk => \N__21159\,
            ce => \N__17501\,
            sr => \N__20805\
        );

    \delay_measurement_inst.delay_hc_timer.counter_27_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17626\,
            in1 => \N__10914\,
            in2 => \_gnd_net_\,
            in3 => \N__9980\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            clk => \N__21159\,
            ce => \N__17501\,
            sr => \N__20805\
        );

    \delay_measurement_inst.delay_hc_timer.counter_28_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17623\,
            in1 => \N__10964\,
            in2 => \_gnd_net_\,
            in3 => \N__9977\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_28\,
            clk => \N__21159\,
            ce => \N__17501\,
            sr => \N__20805\
        );

    \delay_measurement_inst.delay_hc_timer.counter_29_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__10928\,
            in1 => \N__17624\,
            in2 => \_gnd_net_\,
            in3 => \N__9974\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21159\,
            ce => \N__17501\,
            sr => \N__20805\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13162\,
            in2 => \N__11063\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_17_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12902\,
            in2 => \_gnd_net_\,
            in3 => \N__9971\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12866\,
            in2 => \N__11168\,
            in3 => \N__9968\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12833\,
            in2 => \_gnd_net_\,
            in3 => \N__9965\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12803\,
            in2 => \_gnd_net_\,
            in3 => \N__9962\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12776\,
            in3 => \N__9959\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12752\,
            in2 => \_gnd_net_\,
            in3 => \N__10016\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13085\,
            in3 => \N__10013\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13061\,
            in2 => \_gnd_net_\,
            in3 => \N__10010\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9\,
            ltout => OPEN,
            carryin => \bfn_7_18_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13040\,
            in2 => \_gnd_net_\,
            in3 => \N__10007\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13019\,
            in2 => \_gnd_net_\,
            in3 => \N__10004\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12998\,
            in2 => \_gnd_net_\,
            in3 => \N__9992\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12971\,
            in2 => \_gnd_net_\,
            in3 => \N__9989\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12950\,
            in2 => \_gnd_net_\,
            in3 => \N__9986\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13397\,
            in2 => \_gnd_net_\,
            in3 => \N__9983\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13376\,
            in2 => \_gnd_net_\,
            in3 => \N__10037\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13355\,
            in2 => \_gnd_net_\,
            in3 => \N__10034\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17\,
            ltout => OPEN,
            carryin => \bfn_7_19_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13334\,
            in2 => \_gnd_net_\,
            in3 => \N__10031\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13313\,
            in2 => \_gnd_net_\,
            in3 => \N__10028\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_startlto19_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__11707\,
            in1 => \N__11540\,
            in2 => \_gnd_net_\,
            in3 => \N__13712\,
            lcout => \phase_controller_inst1.stoper_tr.un1_start\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_startlto6_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010101010"
        )
    port map (
            in0 => \N__13641\,
            in1 => \N__14906\,
            in2 => \N__15112\,
            in3 => \N__10022\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.un1_startlt8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_startlto9_0_0_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010101010"
        )
    port map (
            in0 => \N__13575\,
            in1 => \N__13467\,
            in2 => \N__10025\,
            in3 => \N__11249\,
            lcout => \phase_controller_inst1.stoper_tr.un1_startlt15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_startlto5_1_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__13418\,
            in1 => \N__13530\,
            in2 => \_gnd_net_\,
            in3 => \N__15020\,
            lcout => \phase_controller_inst1.stoper_tr.un1_startlto5Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un2_startlto19_4_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__15056\,
            in1 => \N__16925\,
            in2 => \_gnd_net_\,
            in3 => \N__13691\,
            lcout => \phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un2_startlto6_0_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13419\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13640\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.un2_startlto6Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un2_startlto6_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__15021\,
            in1 => \N__15107\,
            in2 => \N__10049\,
            in3 => \N__14907\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.un2_startlt19_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un2_startlto19_9_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__10046\,
            in1 => \N__13611\,
            in2 => \N__10040\,
            in3 => \N__14841\,
            lcout => \phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_13_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010000010100000"
        )
    port map (
            in0 => \N__11838\,
            in1 => \N__11541\,
            in2 => \N__14807\,
            in3 => \N__11675\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21133\,
            ce => \N__12031\,
            sr => \N__20824\
        );

    \phase_controller_inst1.stoper_tr.target_time_15_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11674\,
            in2 => \_gnd_net_\,
            in3 => \N__13713\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21133\,
            ce => \N__12031\,
            sr => \N__20824\
        );

    \phase_controller_inst1.stoper_tr.target_time_5_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010101000000"
        )
    port map (
            in0 => \N__10158\,
            in1 => \N__11226\,
            in2 => \N__11206\,
            in3 => \N__13426\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21129\,
            ce => \N__12030\,
            sr => \N__20828\
        );

    \phase_controller_inst1.stoper_tr.target_time_12_LC_7_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__11576\,
            in1 => \N__11701\,
            in2 => \N__11872\,
            in3 => \N__13613\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21129\,
            ce => \N__12030\,
            sr => \N__20828\
        );

    \phase_controller_inst1.stoper_tr.target_time_3_LC_7_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100010001000"
        )
    port map (
            in0 => \N__15111\,
            in1 => \N__11843\,
            in2 => \N__11749\,
            in3 => \N__11578\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21129\,
            ce => \N__12030\,
            sr => \N__20828\
        );

    \phase_controller_inst1.stoper_tr.target_time_14_LC_7_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__11706\,
            in1 => \N__13579\,
            in2 => \_gnd_net_\,
            in3 => \N__13714\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21129\,
            ce => \N__12030\,
            sr => \N__20828\
        );

    \phase_controller_inst1.stoper_tr.target_time_1_LC_7_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000011000000"
        )
    port map (
            in0 => \N__11702\,
            in1 => \N__13537\,
            in2 => \N__11892\,
            in3 => \N__11577\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21129\,
            ce => \N__12030\,
            sr => \N__20828\
        );

    \phase_controller_inst1.stoper_tr.target_time_2_LC_7_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011101010"
        )
    port map (
            in0 => \N__14914\,
            in1 => \N__11198\,
            in2 => \N__11230\,
            in3 => \N__10157\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21129\,
            ce => \N__12030\,
            sr => \N__20828\
        );

    \phase_controller_inst1.stoper_tr.target_timeZ0Z_6_LC_7_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111101110111011"
        )
    port map (
            in0 => \N__13648\,
            in1 => \N__11842\,
            in2 => \N__11748\,
            in3 => \N__11575\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21129\,
            ce => \N__12030\,
            sr => \N__20828\
        );

    \phase_controller_inst1.stoper_tr.target_time_18_LC_7_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15071\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21129\,
            ce => \N__12030\,
            sr => \N__20828\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_7_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10136\,
            in2 => \N__10130\,
            in3 => \N__11973\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_7_23_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_7_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10121\,
            in2 => \N__10115\,
            in3 => \N__11947\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_7_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10106\,
            in2 => \N__10100\,
            in3 => \N__12205\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_7_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11936\,
            in2 => \N__10091\,
            in3 => \N__12169\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_7_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10082\,
            in2 => \N__10076\,
            in3 => \N__12148\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_7_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10067\,
            in2 => \N__10058\,
            in3 => \N__12127\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_7_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11507\,
            in2 => \N__10295\,
            in3 => \N__12106\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_7_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11918\,
            in2 => \N__10286\,
            in3 => \N__12082\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_7_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10277\,
            in2 => \N__10268\,
            in3 => \N__12058\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_7_24_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_7_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10259\,
            in2 => \N__10247\,
            in3 => \N__12397\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_7_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10238\,
            in2 => \N__10229\,
            in3 => \N__12371\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_7_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10220\,
            in2 => \N__10208\,
            in3 => \N__13955\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_7_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10199\,
            in2 => \N__10190\,
            in3 => \N__12344\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_7_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10181\,
            in2 => \N__10169\,
            in3 => \N__12319\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_7_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10376\,
            in2 => \N__10364\,
            in3 => \N__12290\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_7_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11912\,
            in2 => \N__10355\,
            in3 => \N__12266\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_7_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11930\,
            in2 => \N__10346\,
            in3 => \N__12238\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_7_25_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_7_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10337\,
            in2 => \N__10328\,
            in3 => \N__12472\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_7_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10319\,
            in2 => \N__10307\,
            in3 => \N__12451\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_7_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10298\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNI62NA_LC_7_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__15853\,
            in1 => \_gnd_net_\,
            in2 => \N__15935\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNI62NAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_7_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15852\,
            in2 => \_gnd_net_\,
            in3 => \N__15922\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_7_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__15854\,
            in1 => \_gnd_net_\,
            in2 => \N__11984\,
            in3 => \N__15926\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_7_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__15883\,
            in1 => \N__15587\,
            in2 => \N__15740\,
            in3 => \N__12329\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21109\,
            ce => 'H',
            sr => \N__20845\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_7_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__15588\,
            in1 => \N__15729\,
            in2 => \N__12302\,
            in3 => \N__15887\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21109\,
            ce => 'H',
            sr => \N__20845\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_7_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__15884\,
            in1 => \N__15589\,
            in2 => \N__15741\,
            in3 => \N__12275\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21109\,
            ce => 'H',
            sr => \N__20845\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_7_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__15590\,
            in1 => \N__15730\,
            in2 => \N__12251\,
            in3 => \N__15888\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21109\,
            ce => 'H',
            sr => \N__20845\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_7_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__15885\,
            in1 => \N__15591\,
            in2 => \N__15742\,
            in3 => \N__12227\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21109\,
            ce => 'H',
            sr => \N__20845\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_7_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__15592\,
            in1 => \N__15731\,
            in2 => \N__15899\,
            in3 => \N__12461\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21109\,
            ce => 'H',
            sr => \N__20845\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_7_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__15886\,
            in1 => \N__15593\,
            in2 => \N__15743\,
            in3 => \N__12437\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21109\,
            ce => 'H',
            sr => \N__20845\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_7_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__15586\,
            in1 => \N__15728\,
            in2 => \N__15898\,
            in3 => \N__12356\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21109\,
            ce => 'H',
            sr => \N__20845\
        );

    \SB_DFF_inst_PH1_MAX_D1_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10385\,
            lcout => \il_max_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21193\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJHF91_6_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__14005\,
            in1 => \N__14056\,
            in2 => \_gnd_net_\,
            in3 => \N__14341\,
            lcout => \delay_measurement_inst.N_109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17854\,
            in1 => \N__17734\,
            in2 => \N__14326\,
            in3 => \N__13972\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_105\,
            ltout => \delay_measurement_inst.delay_hc_timer.N_105_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4TEU1_9_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010101"
        )
    port map (
            in0 => \N__18031\,
            in1 => \N__14082\,
            in2 => \N__10493\,
            in3 => \N__14116\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_4_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12667\,
            in1 => \N__14182\,
            in2 => \N__12698\,
            in3 => \N__14410\,
            lcout => \delay_measurement_inst.delay_hc_timer.un1_reset_1_i_a2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10489\,
            in2 => \N__10450\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.elapsed_time_hc_3\,
            ltout => OPEN,
            carryin => \bfn_8_13_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__21175\,
            ce => \N__10888\,
            sr => \N__20784\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10471\,
            in2 => \N__10426\,
            in3 => \N__10454\,
            lcout => \delay_measurement_inst.elapsed_time_hc_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__21175\,
            ce => \N__10888\,
            sr => \N__20784\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10401\,
            in2 => \N__10451\,
            in3 => \N__10430\,
            lcout => \delay_measurement_inst.elapsed_time_hc_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__21175\,
            ce => \N__10888\,
            sr => \N__20784\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10665\,
            in2 => \N__10427\,
            in3 => \N__10406\,
            lcout => \delay_measurement_inst.elapsed_time_hc_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__21175\,
            ce => \N__10888\,
            sr => \N__20784\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10402\,
            in2 => \N__10648\,
            in3 => \N__10388\,
            lcout => \delay_measurement_inst.elapsed_time_hc_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__21175\,
            ce => \N__10888\,
            sr => \N__20784\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10666\,
            in2 => \N__10624\,
            in3 => \N__10652\,
            lcout => \delay_measurement_inst.elapsed_time_hc_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__21175\,
            ce => \N__10888\,
            sr => \N__20784\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10599\,
            in2 => \N__10649\,
            in3 => \N__10628\,
            lcout => \delay_measurement_inst.elapsed_time_hc_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__21175\,
            ce => \N__10888\,
            sr => \N__20784\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10578\,
            in2 => \N__10625\,
            in3 => \N__10604\,
            lcout => \delay_measurement_inst.elapsed_time_hc_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__21175\,
            ce => \N__10888\,
            sr => \N__20784\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10601\,
            in2 => \N__10558\,
            in3 => \N__10583\,
            lcout => \delay_measurement_inst.elapsed_time_hc_11\,
            ltout => OPEN,
            carryin => \bfn_8_14_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__21167\,
            ce => \N__10887\,
            sr => \N__20789\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10580\,
            in2 => \N__10534\,
            in3 => \N__10562\,
            lcout => \delay_measurement_inst.elapsed_time_hc_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__21167\,
            ce => \N__10887\,
            sr => \N__20789\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10509\,
            in2 => \N__10559\,
            in3 => \N__10538\,
            lcout => \delay_measurement_inst.elapsed_time_hc_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__21167\,
            ce => \N__10887\,
            sr => \N__20789\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10857\,
            in2 => \N__10535\,
            in3 => \N__10514\,
            lcout => \delay_measurement_inst.elapsed_time_hc_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__21167\,
            ce => \N__10887\,
            sr => \N__20789\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10510\,
            in2 => \N__10840\,
            in3 => \N__10496\,
            lcout => \delay_measurement_inst.elapsed_time_hc_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__21167\,
            ce => \N__10887\,
            sr => \N__20789\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10858\,
            in2 => \N__10816\,
            in3 => \N__10844\,
            lcout => \delay_measurement_inst.elapsed_time_hc_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__21167\,
            ce => \N__10887\,
            sr => \N__20789\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10791\,
            in2 => \N__10841\,
            in3 => \N__10820\,
            lcout => \delay_measurement_inst.elapsed_time_hc_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__21167\,
            ce => \N__10887\,
            sr => \N__20789\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10770\,
            in2 => \N__10817\,
            in3 => \N__10796\,
            lcout => \delay_measurement_inst.elapsed_time_hc_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__21167\,
            ce => \N__10887\,
            sr => \N__20789\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10793\,
            in2 => \N__10750\,
            in3 => \N__10775\,
            lcout => \delay_measurement_inst.elapsed_time_hc_19\,
            ltout => OPEN,
            carryin => \bfn_8_15_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__21160\,
            ce => \N__10886\,
            sr => \N__20794\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10772\,
            in2 => \N__10726\,
            in3 => \N__10754\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__21160\,
            ce => \N__10886\,
            sr => \N__20794\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10701\,
            in2 => \N__10751\,
            in3 => \N__10730\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__21160\,
            ce => \N__10886\,
            sr => \N__20794\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10683\,
            in2 => \N__10727\,
            in3 => \N__10706\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__21160\,
            ce => \N__10886\,
            sr => \N__20794\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10702\,
            in2 => \N__11053\,
            in3 => \N__10688\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__21160\,
            ce => \N__10886\,
            sr => \N__20794\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10684\,
            in2 => \N__11029\,
            in3 => \N__10670\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__21160\,
            ce => \N__10886\,
            sr => \N__20794\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11004\,
            in2 => \N__11054\,
            in3 => \N__11033\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__21160\,
            ce => \N__10886\,
            sr => \N__20794\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10983\,
            in2 => \N__11030\,
            in3 => \N__11009\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__21160\,
            ce => \N__10886\,
            sr => \N__20794\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11006\,
            in2 => \N__10951\,
            in3 => \N__10988\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\,
            ltout => OPEN,
            carryin => \bfn_8_16_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__21153\,
            ce => \N__10885\,
            sr => \N__20801\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10985\,
            in2 => \N__10915\,
            in3 => \N__10967\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__21153\,
            ce => \N__10885\,
            sr => \N__20801\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10963\,
            in2 => \N__10952\,
            in3 => \N__10931\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__21153\,
            ce => \N__10885\,
            sr => \N__20801\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10927\,
            in2 => \N__10916\,
            in3 => \N__10895\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__21153\,
            ce => \N__10885\,
            sr => \N__20801\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10892\,
            lcout => \delay_measurement_inst.elapsed_time_hc_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21153\,
            ce => \N__10885\,
            sr => \N__20801\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_3_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__13281\,
            in1 => \N__11461\,
            in2 => \N__10868\,
            in3 => \N__11322\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21146\,
            ce => 'H',
            sr => \N__20806\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_4_LC_8_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__11458\,
            in1 => \N__13285\,
            in2 => \N__11356\,
            in3 => \N__11108\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21146\,
            ce => 'H',
            sr => \N__20806\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_5_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__13282\,
            in1 => \N__11462\,
            in2 => \N__11102\,
            in3 => \N__11323\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21146\,
            ce => 'H',
            sr => \N__20806\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_6_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__11459\,
            in1 => \N__13286\,
            in2 => \N__11357\,
            in3 => \N__11093\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21146\,
            ce => 'H',
            sr => \N__20806\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_7_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__13283\,
            in1 => \N__11463\,
            in2 => \N__11087\,
            in3 => \N__11324\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21146\,
            ce => 'H',
            sr => \N__20806\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_8_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__11460\,
            in1 => \N__13287\,
            in2 => \N__11358\,
            in3 => \N__11078\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21146\,
            ce => 'H',
            sr => \N__20806\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_9_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__13284\,
            in1 => \N__11464\,
            in2 => \N__11072\,
            in3 => \N__11325\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21146\,
            ce => 'H',
            sr => \N__20806\
        );

    \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_1_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000100"
        )
    port map (
            in0 => \N__11312\,
            in1 => \N__11429\,
            in2 => \N__13274\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_hc.stoper_state_RNI10KLZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_1_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__13228\,
            in1 => \N__11466\,
            in2 => \N__13115\,
            in3 => \N__11337\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21143\,
            ce => 'H',
            sr => \N__20809\
        );

    \phase_controller_slave.stoper_hc.stoper_state_0_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__13139\,
            in1 => \N__11332\,
            in2 => \N__13271\,
            in3 => \N__11468\,
            lcout => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21143\,
            ce => 'H',
            sr => \N__20809\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_8_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13225\,
            in2 => \_gnd_net_\,
            in3 => \N__13137\,
            lcout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.stoper_state_1_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001110000010000"
        )
    port map (
            in0 => \N__13140\,
            in1 => \N__11333\,
            in2 => \N__13272\,
            in3 => \N__11469\,
            lcout => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21143\,
            ce => 'H',
            sr => \N__20809\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNI89DK_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13226\,
            in2 => \_gnd_net_\,
            in3 => \N__13138\,
            lcout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNI89DKZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_10_LC_8_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__13227\,
            in1 => \N__11331\,
            in2 => \N__11159\,
            in3 => \N__11467\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21143\,
            ce => 'H',
            sr => \N__20809\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_11_LC_8_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__11465\,
            in1 => \N__13229\,
            in2 => \N__11361\,
            in3 => \N__11150\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21143\,
            ce => 'H',
            sr => \N__20809\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_13_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__13248\,
            in1 => \N__11474\,
            in2 => \N__11362\,
            in3 => \N__11144\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21139\,
            ce => 'H',
            sr => \N__20810\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_14_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011010000"
        )
    port map (
            in0 => \N__11470\,
            in1 => \N__13252\,
            in2 => \N__11138\,
            in3 => \N__11350\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21139\,
            ce => 'H',
            sr => \N__20810\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_15_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__13249\,
            in1 => \N__11475\,
            in2 => \N__11363\,
            in3 => \N__11129\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21139\,
            ce => 'H',
            sr => \N__20810\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_16_LC_8_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011010000"
        )
    port map (
            in0 => \N__11471\,
            in1 => \N__13253\,
            in2 => \N__11123\,
            in3 => \N__11351\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21139\,
            ce => 'H',
            sr => \N__20810\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_17_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__13250\,
            in1 => \N__11476\,
            in2 => \N__11364\,
            in3 => \N__11114\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21139\,
            ce => 'H',
            sr => \N__20810\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_18_LC_8_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__11472\,
            in1 => \N__13254\,
            in2 => \N__11366\,
            in3 => \N__11489\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21139\,
            ce => 'H',
            sr => \N__20810\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_19_LC_8_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__13251\,
            in1 => \N__11477\,
            in2 => \N__11365\,
            in3 => \N__11483\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21139\,
            ce => 'H',
            sr => \N__20810\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_2_LC_8_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011010000"
        )
    port map (
            in0 => \N__11473\,
            in1 => \N__13255\,
            in2 => \N__11378\,
            in3 => \N__11352\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21139\,
            ce => 'H',
            sr => \N__20810\
        );

    \phase_controller_inst1.stoper_tr.un1_startlto9_c_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__13456\,
            in1 => \N__12623\,
            in2 => \_gnd_net_\,
            in3 => \N__13794\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.un1_startlto9_cZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_startlto13_3_LC_8_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__13601\,
            in1 => \N__14837\,
            in2 => \N__11252\,
            in3 => \N__13816\,
            lcout => \phase_controller_inst1.stoper_tr.un1_startlto13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un2_startlto19_6_LC_8_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12631\,
            in1 => \N__13457\,
            in2 => \N__13798\,
            in3 => \N__13557\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un2_startlto19_8_LC_8_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__13753\,
            in1 => \N__13496\,
            in2 => \N__11243\,
            in3 => \N__13817\,
            lcout => \phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_8\,
            ltout => \phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_start_0_LC_8_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__11673\,
            in1 => \N__13687\,
            in2 => \N__11210\,
            in3 => \N__11181\,
            lcout => \phase_controller_inst1.stoper_tr.un3_start\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_startlto19_2_LC_8_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13752\,
            in1 => \N__16926\,
            in2 => \N__13503\,
            in3 => \N__15067\,
            lcout => \phase_controller_inst1.stoper_tr.un1_startlto19Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_LC_8_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100010001000"
        )
    port map (
            in0 => \N__11839\,
            in1 => \N__15028\,
            in2 => \N__11745\,
            in3 => \N__11583\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21125\,
            ce => \N__12016\,
            sr => \N__20825\
        );

    \phase_controller_inst1.stoper_tr.target_time_17_LC_8_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13504\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21125\,
            ce => \N__12016\,
            sr => \N__20825\
        );

    \phase_controller_inst1.stoper_tr.target_time_8_LC_8_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100010001000"
        )
    port map (
            in0 => \N__11841\,
            in1 => \N__12632\,
            in2 => \N__11747\,
            in3 => \N__11585\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21125\,
            ce => \N__12016\,
            sr => \N__20825\
        );

    \phase_controller_inst1.stoper_tr.target_time_16_LC_8_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13748\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21125\,
            ce => \N__12016\,
            sr => \N__20825\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_LC_8_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100010001000"
        )
    port map (
            in0 => \N__11840\,
            in1 => \N__13792\,
            in2 => \N__11746\,
            in3 => \N__11584\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21125\,
            ce => \N__12016\,
            sr => \N__20825\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_8_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__15560\,
            in1 => \N__15713\,
            in2 => \N__11501\,
            in3 => \N__15851\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21119\,
            ce => 'H',
            sr => \N__20829\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_0_LC_8_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001000000010"
        )
    port map (
            in0 => \N__15562\,
            in1 => \N__15714\,
            in2 => \N__15897\,
            in3 => \N__15936\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21119\,
            ce => 'H',
            sr => \N__20829\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_8_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__15559\,
            in1 => \N__15712\,
            in2 => \N__12386\,
            in3 => \N__15850\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21119\,
            ce => 'H',
            sr => \N__20829\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_8_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__15849\,
            in1 => \N__15561\,
            in2 => \N__15739\,
            in3 => \N__12218\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21119\,
            ce => 'H',
            sr => \N__20829\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_8_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__15828\,
            in1 => \N__15552\,
            in2 => \N__15735\,
            in3 => \N__12179\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21114\,
            ce => 'H',
            sr => \N__20834\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_8_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__15553\,
            in1 => \N__15832\,
            in2 => \N__15732\,
            in3 => \N__12158\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21114\,
            ce => 'H',
            sr => \N__20834\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_8_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__15829\,
            in1 => \N__15554\,
            in2 => \N__15736\,
            in3 => \N__12137\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21114\,
            ce => 'H',
            sr => \N__20834\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_8_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__15555\,
            in1 => \N__15833\,
            in2 => \N__15733\,
            in3 => \N__12116\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21114\,
            ce => 'H',
            sr => \N__20834\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_8_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__15830\,
            in1 => \N__15556\,
            in2 => \N__15737\,
            in3 => \N__12095\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21114\,
            ce => 'H',
            sr => \N__20834\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_8_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__15557\,
            in1 => \N__15834\,
            in2 => \N__15734\,
            in3 => \N__12071\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21114\,
            ce => 'H',
            sr => \N__20834\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_8_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__15831\,
            in1 => \N__15558\,
            in2 => \N__15738\,
            in3 => \N__12047\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21114\,
            ce => 'H',
            sr => \N__20834\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_1_LC_8_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__15687\,
            in1 => \N__15550\,
            in2 => \_gnd_net_\,
            in3 => \N__15827\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJMZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_8_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11980\,
            in2 => \N__11960\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_25_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_8_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11951\,
            in2 => \_gnd_net_\,
            in3 => \N__12209\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_8_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12206\,
            in2 => \N__12188\,
            in3 => \N__12173\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_8_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12170\,
            in2 => \_gnd_net_\,
            in3 => \N__12152\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_8_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12149\,
            in2 => \_gnd_net_\,
            in3 => \N__12131\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_8_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12128\,
            in2 => \_gnd_net_\,
            in3 => \N__12110\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_8_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12107\,
            in2 => \_gnd_net_\,
            in3 => \N__12089\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_8_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12086\,
            in2 => \_gnd_net_\,
            in3 => \N__12065\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_8_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12062\,
            in2 => \_gnd_net_\,
            in3 => \N__12038\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\,
            ltout => OPEN,
            carryin => \bfn_8_26_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_8_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12401\,
            in2 => \_gnd_net_\,
            in3 => \N__12374\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_8_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12370\,
            in2 => \_gnd_net_\,
            in3 => \N__12350\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_8_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13951\,
            in2 => \_gnd_net_\,
            in3 => \N__12347\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_8_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12343\,
            in2 => \_gnd_net_\,
            in3 => \N__12323\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_8_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12320\,
            in3 => \N__12293\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_8_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12289\,
            in2 => \_gnd_net_\,
            in3 => \N__12269\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_8_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12265\,
            in2 => \_gnd_net_\,
            in3 => \N__12242\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_8_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12239\,
            in2 => \_gnd_net_\,
            in3 => \N__12221\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\,
            ltout => OPEN,
            carryin => \bfn_8_27_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_8_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12473\,
            in2 => \_gnd_net_\,
            in3 => \N__12455\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_8_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12452\,
            in2 => \_gnd_net_\,
            in3 => \N__12440\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_tr_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__20892\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13850\,
            lcout => \delay_measurement_inst.stop_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21191\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15477\,
            in2 => \_gnd_net_\,
            in3 => \N__17039\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_180_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D1_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12410\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_min_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21191\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.tr_sync_1_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18857\,
            lcout => \delay_measurement_inst.tr_syncZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21187\,
            ce => 'H',
            sr => \N__20769\
        );

    \delay_measurement_inst.tr_prev_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13883\,
            lcout => \delay_measurement_inst.tr_prevZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21187\,
            ce => 'H',
            sr => \N__20769\
        );

    \delay_measurement_inst.tr_state_0_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000000110"
        )
    port map (
            in0 => \N__13881\,
            in1 => \N__14167\,
            in2 => \N__20903\,
            in3 => \N__14152\,
            lcout => \delay_measurement_inst.tr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21182\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.tr_state_RNIVV8G_0_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__13880\,
            in1 => \N__14166\,
            in2 => \_gnd_net_\,
            in3 => \N__14151\,
            lcout => \delay_measurement_inst.tr_state_RNIVV8GZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJQC01_31_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__20894\,
            in1 => \N__17794\,
            in2 => \_gnd_net_\,
            in3 => \N__15381\,
            lcout => \delay_measurement_inst.delay_hc_timer.un1_reset_1_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__14365\,
            in1 => \N__12696\,
            in2 => \N__12671\,
            in3 => \N__14397\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_81\,
            ltout => \delay_measurement_inst.delay_hc_timer.N_81_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE5L06_31_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111110"
        )
    port map (
            in0 => \N__17798\,
            in1 => \N__12533\,
            in2 => \N__12527\,
            in3 => \N__17962\,
            lcout => \delay_measurement_inst.N_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBM7A4_14_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111010"
        )
    port map (
            in0 => \N__17961\,
            in1 => \N__15400\,
            in2 => \N__18039\,
            in3 => \N__14115\,
            lcout => \delay_measurement_inst.N_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI40E01_17_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14114\,
            in1 => \N__14364\,
            in2 => \N__14399\,
            in3 => \N__18024\,
            lcout => \delay_measurement_inst.delay_hc_timer.un1_reset_1_i_a2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKF324_15_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__17963\,
            in1 => \_gnd_net_\,
            in2 => \N__18038\,
            in3 => \N__12509\,
            lcout => \delay_measurement_inst.N_107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE9BL2_2_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000000"
        )
    port map (
            in0 => \N__12643\,
            in1 => \N__12487\,
            in2 => \N__14086\,
            in3 => \N__12524\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un1_reset_1_i_a2_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJTHF5_17_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__15388\,
            in1 => \N__14279\,
            in2 => \N__12518\,
            in3 => \N__12515\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un1_reset_1_i_a2_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQOU9A_31_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__12508\,
            in1 => \N__12500\,
            in2 => \N__12494\,
            in3 => \N__17960\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_esr_2_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__14283\,
            in1 => \N__14253\,
            in2 => \N__14223\,
            in3 => \N__12491\,
            lcout => measured_delay_hc_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21168\,
            ce => \N__17686\,
            sr => \N__17658\
        );

    \delay_measurement_inst.delay_hc_reg_esr_19_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__17965\,
            in1 => \N__17796\,
            in2 => \_gnd_net_\,
            in3 => \N__12697\,
            lcout => measured_delay_hc_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21168\,
            ce => \N__17686\,
            sr => \N__17658\
        );

    \delay_measurement_inst.delay_hc_reg_esr_16_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__17795\,
            in1 => \N__17964\,
            in2 => \_gnd_net_\,
            in3 => \N__12666\,
            lcout => measured_delay_hc_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21168\,
            ce => \N__17686\,
            sr => \N__17658\
        );

    \delay_measurement_inst.delay_hc_reg_ess_3_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__14254\,
            in1 => \N__12644\,
            in2 => \N__14303\,
            in3 => \N__14211\,
            lcout => measured_delay_hc_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21168\,
            ce => \N__17686\,
            sr => \N__17658\
        );

    \delay_measurement_inst.delay_tr_reg_8_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__14996\,
            in1 => \N__19850\,
            in2 => \N__15332\,
            in3 => \N__12611\,
            lcout => measured_delay_tr_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21161\,
            ce => 'H',
            sr => \N__17185\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__12587\,
            in1 => \N__12581\,
            in2 => \N__12575\,
            in3 => \N__12566\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg_5_0_o2_0_7_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_16_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16261\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21154\,
            ce => \N__18772\,
            sr => \N__20790\
        );

    \phase_controller_inst1.stoper_hc.target_time_17_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16195\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21154\,
            ce => \N__18772\,
            sr => \N__20790\
        );

    \phase_controller_inst1.stoper_hc.target_time_18_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16166\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21154\,
            ce => \N__18772\,
            sr => \N__20790\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAAI01_25_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__12560\,
            in1 => \N__12554\,
            in2 => \N__12548\,
            in3 => \N__12539\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg_5_0_o2_0_6_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__12731\,
            in1 => \N__12725\,
            in2 => \N__12719\,
            in3 => \N__12704\,
            lcout => \delay_measurement_inst.N_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI23AG_29_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12716\,
            in2 => \_gnd_net_\,
            in3 => \N__12710\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg_5_0_o2_0_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_19_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16228\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21154\,
            ce => \N__18772\,
            sr => \N__20790\
        );

    \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111101110111011"
        )
    port map (
            in0 => \N__16846\,
            in1 => \N__16609\,
            in2 => \N__16442\,
            in3 => \N__16717\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21147\,
            ce => \N__15141\,
            sr => \N__20795\
        );

    \phase_controller_slave.stoper_hc.target_time_4_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__16720\,
            in1 => \N__16436\,
            in2 => \N__16622\,
            in3 => \N__17362\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21147\,
            ce => \N__15141\,
            sr => \N__20795\
        );

    \phase_controller_slave.stoper_hc.target_time_8_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000011000000"
        )
    port map (
            in0 => \N__16437\,
            in1 => \N__16610\,
            in2 => \N__16106\,
            in3 => \N__16721\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21147\,
            ce => \N__15141\,
            sr => \N__20795\
        );

    \phase_controller_slave.stoper_hc.target_time_2_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011101010"
        )
    port map (
            in0 => \N__17453\,
            in1 => \N__17238\,
            in2 => \N__16016\,
            in3 => \N__16132\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21147\,
            ce => \N__15141\,
            sr => \N__20795\
        );

    \phase_controller_slave.stoper_hc.target_time_5_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010101000000"
        )
    port map (
            in0 => \N__16133\,
            in1 => \N__16015\,
            in2 => \N__17243\,
            in3 => \N__16289\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21147\,
            ce => \N__15141\,
            sr => \N__20795\
        );

    \phase_controller_slave.stoper_hc.target_time_1_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__16718\,
            in1 => \N__16434\,
            in2 => \N__16620\,
            in3 => \N__15980\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21147\,
            ce => \N__15141\,
            sr => \N__20795\
        );

    \phase_controller_slave.stoper_hc.target_time_3_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__16719\,
            in1 => \N__16435\,
            in2 => \N__16621\,
            in3 => \N__17399\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21147\,
            ce => \N__15141\,
            sr => \N__20795\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12929\,
            in2 => \N__12920\,
            in3 => \N__13161\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_9_17_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12911\,
            in2 => \N__12884\,
            in3 => \N__12901\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12875\,
            in2 => \N__12851\,
            in3 => \N__12862\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12842\,
            in2 => \N__12821\,
            in3 => \N__12832\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12812\,
            in2 => \N__12791\,
            in3 => \N__12802\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12782\,
            in2 => \N__12761\,
            in3 => \N__12772\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14756\,
            in2 => \N__12740\,
            in3 => \N__12751\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13094\,
            in2 => \N__13070\,
            in3 => \N__13081\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14750\,
            in2 => \N__13049\,
            in3 => \N__13060\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_9_18_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14744\,
            in2 => \N__13028\,
            in3 => \N__13039\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14765\,
            in2 => \N__13007\,
            in3 => \N__13018\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14609\,
            in2 => \N__12980\,
            in3 => \N__12997\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15149\,
            in2 => \N__12959\,
            in3 => \N__12970\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14726\,
            in2 => \N__12938\,
            in3 => \N__12949\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14735\,
            in2 => \N__13385\,
            in3 => \N__13396\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14717\,
            in2 => \N__13364\,
            in3 => \N__13375\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14708\,
            in2 => \N__13343\,
            in3 => \N__13354\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_9_19_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14702\,
            in2 => \N__13322\,
            in3 => \N__13333\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14603\,
            in2 => \N__13301\,
            in3 => \N__13312\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13292\,
            lcout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__13273\,
            in1 => \N__13163\,
            in2 => \_gnd_net_\,
            in3 => \N__13141\,
            lcout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI43GB_6_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__19021\,
            in1 => \N__19843\,
            in2 => \_gnd_net_\,
            in3 => \N__19891\,
            lcout => \delay_measurement_inst.N_172\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D2_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13106\,
            lcout => \il_min_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21134\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_15_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011010000"
        )
    port map (
            in0 => \N__16980\,
            in1 => \N__21679\,
            in2 => \N__20261\,
            in3 => \N__15343\,
            lcout => measured_delay_tr_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21130\,
            ce => \N__16892\,
            sr => \N__17179\
        );

    \delay_measurement_inst.delay_tr_reg_esr_6_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001110101111"
        )
    port map (
            in0 => \N__19025\,
            in1 => \N__15280\,
            in2 => \N__14995\,
            in3 => \N__14946\,
            lcout => measured_delay_tr_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21130\,
            ce => \N__16892\,
            sr => \N__17179\
        );

    \delay_measurement_inst.delay_tr_reg_esr_12_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__21670\,
            in1 => \N__19657\,
            in2 => \_gnd_net_\,
            in3 => \N__15364\,
            lcout => measured_delay_tr_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21130\,
            ce => \N__16892\,
            sr => \N__17179\
        );

    \delay_measurement_inst.delay_tr_reg_esr_14_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__19556\,
            in1 => \N__21671\,
            in2 => \N__15344\,
            in3 => \N__16982\,
            lcout => measured_delay_tr_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21130\,
            ce => \N__16892\,
            sr => \N__17179\
        );

    \delay_measurement_inst.delay_tr_reg_ess_1_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111000010000000"
        )
    port map (
            in0 => \N__14947\,
            in1 => \N__15279\,
            in2 => \N__17018\,
            in3 => \N__14987\,
            lcout => measured_delay_tr_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21130\,
            ce => \N__16892\,
            sr => \N__17179\
        );

    \delay_measurement_inst.delay_tr_reg_esr_17_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__21678\,
            in1 => \N__16981\,
            in2 => \_gnd_net_\,
            in3 => \N__20130\,
            lcout => measured_delay_tr_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21130\,
            ce => \N__16892\,
            sr => \N__17179\
        );

    \delay_measurement_inst.delay_tr_reg_esr_9_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000100"
        )
    port map (
            in0 => \N__15281\,
            in1 => \N__15365\,
            in2 => \N__21683\,
            in3 => \N__19802\,
            lcout => measured_delay_tr_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21130\,
            ce => \N__16892\,
            sr => \N__17179\
        );

    \delay_measurement_inst.delay_tr_reg_esr_5_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101000000000"
        )
    port map (
            in0 => \N__14983\,
            in1 => \N__14945\,
            in2 => \N__15284\,
            in3 => \N__19073\,
            lcout => measured_delay_tr_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21130\,
            ce => \N__16892\,
            sr => \N__17179\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIF26P1_16_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20188\,
            in1 => \N__20259\,
            in2 => \N__20083\,
            in3 => \N__19557\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.un1_reset_i_a2_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUEN44_2_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__14951\,
            in1 => \N__13852\,
            in2 => \N__13862\,
            in3 => \N__14771\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.un1_reset_i_a2_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6L42C_31_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__15300\,
            in1 => \N__13823\,
            in2 => \N__13859\,
            in3 => \N__16974\,
            lcout => \delay_measurement_inst.elapsed_time_ns_1_RNI6L42C_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.tr_state_RNIVV8G_0_0_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13853\,
            lcout => \delay_measurement_inst.N_134_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010101"
        )
    port map (
            in0 => \N__20260\,
            in1 => \N__19797\,
            in2 => \N__15302\,
            in3 => \N__19558\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.N_160_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111010"
        )
    port map (
            in0 => \N__21665\,
            in1 => \N__16975\,
            in2 => \N__13856\,
            in3 => \N__17108\,
            lcout => \delay_measurement_inst.N_129\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVOI61_31_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__20898\,
            in1 => \N__21664\,
            in2 => \_gnd_net_\,
            in3 => \N__13851\,
            lcout => \delay_measurement_inst.delay_tr_timer.un1_reset_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un2_startlto19_2_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14787\,
            in2 => \_gnd_net_\,
            in3 => \N__14862\,
            lcout => \phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_7_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__15325\,
            in1 => \N__14991\,
            in2 => \N__19898\,
            in3 => \N__13793\,
            lcout => measured_delay_tr_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21120\,
            ce => 'H',
            sr => \N__17186\
        );

    \delay_measurement_inst.delay_tr_reg_esr_16_LC_9_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__16985\,
            in1 => \N__21682\,
            in2 => \_gnd_net_\,
            in3 => \N__20189\,
            lcout => measured_delay_tr_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21115\,
            ce => \N__16891\,
            sr => \N__17172\
        );

    \phase_controller_inst1.start_timer_tr_LC_9_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000100"
        )
    port map (
            in0 => \N__18547\,
            in1 => \N__15566\,
            in2 => \N__21488\,
            in3 => \N__15210\,
            lcout => \phase_controller_inst1.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21110\,
            ce => 'H',
            sr => \N__20830\
        );

    \phase_controller_inst1.state_RNI7NN7_0_LC_9_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15761\,
            in2 => \_gnd_net_\,
            in3 => \N__15189\,
            lcout => \phase_controller_inst1.N_108\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_0_LC_9_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001000100010"
        )
    port map (
            in0 => \N__15190\,
            in1 => \N__15762\,
            in2 => \N__15245\,
            in3 => \N__18976\,
            lcout => \phase_controller_inst1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21106\,
            ce => 'H',
            sr => \N__20835\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_9_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__15551\,
            in1 => \N__15882\,
            in2 => \N__15686\,
            in3 => \N__13961\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21106\,
            ce => 'H',
            sr => \N__20835\
        );

    \phase_controller_slave.S1_LC_9_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13937\,
            lcout => s3_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21100\,
            ce => 'H',
            sr => \N__20846\
        );

    \delay_measurement_inst.delay_tr_timer.running_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__15481\,
            in1 => \N__15461\,
            in2 => \_gnd_net_\,
            in3 => \N__17044\,
            lcout => \delay_measurement_inst.delay_tr_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21183\,
            ce => 'H',
            sr => \N__20760\
        );

    \delay_measurement_inst.hc_state_RNIE29G_0_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__15419\,
            in1 => \N__14130\,
            in2 => \_gnd_net_\,
            in3 => \N__15432\,
            lcout => \delay_measurement_inst.N_54\,
            ltout => \delay_measurement_inst.N_54_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.hc_state_RNIE29G_0_0_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13886\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.N_54_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.start_timer_hc_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__15434\,
            in1 => \N__20890\,
            in2 => \N__14138\,
            in3 => \N__15421\,
            lcout => \delay_measurement_inst.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21177\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.start_timer_tr_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__13882\,
            in1 => \N__20891\,
            in2 => \N__14171\,
            in3 => \N__14153\,
            lcout => \delay_measurement_inst.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21177\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.hc_state_0_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000100110000"
        )
    port map (
            in0 => \N__15433\,
            in1 => \N__20889\,
            in2 => \N__14137\,
            in3 => \N__15420\,
            lcout => \delay_measurement_inst.hc_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21177\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_esr_14_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__17833\,
            in1 => \N__14120\,
            in2 => \N__17996\,
            in3 => \N__17974\,
            lcout => measured_delay_hc_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21170\,
            ce => \N__17681\,
            sr => \N__17656\
        );

    \delay_measurement_inst.delay_hc_reg_esr_9_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000100"
        )
    port map (
            in0 => \N__14210\,
            in1 => \N__17710\,
            in2 => \N__17837\,
            in3 => \N__14090\,
            lcout => measured_delay_hc_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21170\,
            ce => \N__17681\,
            sr => \N__17656\
        );

    \delay_measurement_inst.delay_hc_reg_7_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__14251\,
            in1 => \N__14063\,
            in2 => \N__16064\,
            in3 => \N__14026\,
            lcout => measured_delay_hc_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21162\,
            ce => 'H',
            sr => \N__17657\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8R7QA_31_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14025\,
            in2 => \_gnd_net_\,
            in3 => \N__14041\,
            lcout => \delay_measurement_inst.N_54_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_8_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__14027\,
            in1 => \N__14012\,
            in2 => \N__16102\,
            in3 => \N__14252\,
            lcout => measured_delay_hc_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21162\,
            ce => 'H',
            sr => \N__17657\
        );

    \delay_measurement_inst.delay_hc_reg_ess_1_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110000010100000"
        )
    port map (
            in0 => \N__14258\,
            in1 => \N__14215\,
            in2 => \N__13994\,
            in3 => \N__14302\,
            lcout => measured_delay_hc_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21155\,
            ce => \N__17682\,
            sr => \N__17659\
        );

    \delay_measurement_inst.delay_hc_reg_esr_10_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__13976\,
            in1 => \N__17821\,
            in2 => \_gnd_net_\,
            in3 => \N__17708\,
            lcout => measured_delay_hc_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21155\,
            ce => \N__17682\,
            sr => \N__17659\
        );

    \delay_measurement_inst.delay_hc_reg_esr_4_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000010100000"
        )
    port map (
            in0 => \N__14255\,
            in1 => \N__14301\,
            in2 => \N__14417\,
            in3 => \N__14222\,
            lcout => measured_delay_hc_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21155\,
            ce => \N__17682\,
            sr => \N__17659\
        );

    \delay_measurement_inst.delay_hc_reg_esr_18_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__17973\,
            in1 => \N__17826\,
            in2 => \_gnd_net_\,
            in3 => \N__14398\,
            lcout => measured_delay_hc_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21155\,
            ce => \N__17682\,
            sr => \N__17659\
        );

    \delay_measurement_inst.delay_hc_reg_esr_17_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__17825\,
            in1 => \N__14369\,
            in2 => \_gnd_net_\,
            in3 => \N__17972\,
            lcout => measured_delay_hc_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21155\,
            ce => \N__17682\,
            sr => \N__17659\
        );

    \delay_measurement_inst.delay_hc_reg_esr_6_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111100010011"
        )
    port map (
            in0 => \N__14300\,
            in1 => \N__14257\,
            in2 => \N__14225\,
            in3 => \N__14345\,
            lcout => measured_delay_hc_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21155\,
            ce => \N__17682\,
            sr => \N__17659\
        );

    \delay_measurement_inst.delay_hc_reg_esr_13_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010100000000"
        )
    port map (
            in0 => \N__17709\,
            in1 => \_gnd_net_\,
            in2 => \N__17832\,
            in3 => \N__14330\,
            lcout => measured_delay_hc_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21155\,
            ce => \N__17682\,
            sr => \N__17659\
        );

    \delay_measurement_inst.delay_hc_reg_esr_5_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__14299\,
            in1 => \N__14256\,
            in2 => \N__14224\,
            in3 => \N__14186\,
            lcout => measured_delay_hc_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21155\,
            ce => \N__17682\,
            sr => \N__17659\
        );

    \phase_controller_inst1.stoper_hc.target_time_3_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010000010100000"
        )
    port map (
            in0 => \N__16562\,
            in1 => \N__16355\,
            in2 => \N__17400\,
            in3 => \N__16682\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21149\,
            ce => \N__18773\,
            sr => \N__20779\
        );

    \phase_controller_inst1.stoper_hc.target_time_5_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010101000000"
        )
    port map (
            in0 => \N__16123\,
            in1 => \N__16005\,
            in2 => \N__17242\,
            in3 => \N__16285\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21149\,
            ce => \N__18773\,
            sr => \N__20779\
        );

    \phase_controller_inst1.stoper_hc.target_time_8_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100110000000000"
        )
    port map (
            in0 => \N__16685\,
            in1 => \N__16565\,
            in2 => \N__16400\,
            in3 => \N__16101\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21149\,
            ce => \N__18773\,
            sr => \N__20779\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010000010100000"
        )
    port map (
            in0 => \N__16563\,
            in1 => \N__16356\,
            in2 => \N__17363\,
            in3 => \N__16683\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21149\,
            ce => \N__18773\,
            sr => \N__20779\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100110000000000"
        )
    port map (
            in0 => \N__16684\,
            in1 => \N__16564\,
            in2 => \N__16399\,
            in3 => \N__16063\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21149\,
            ce => \N__18773\,
            sr => \N__20779\
        );

    \phase_controller_inst1.stoper_hc.target_time_2_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011101010"
        )
    port map (
            in0 => \N__17438\,
            in1 => \N__17234\,
            in2 => \N__16011\,
            in3 => \N__16122\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21149\,
            ce => \N__18773\,
            sr => \N__20779\
        );

    \phase_controller_inst1.stoper_hc.target_time_1_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100110000000000"
        )
    port map (
            in0 => \N__16681\,
            in1 => \N__15973\,
            in2 => \N__16398\,
            in3 => \N__16566\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21149\,
            ce => \N__18773\,
            sr => \N__20779\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14498\,
            in2 => \N__14492\,
            in3 => \N__18246\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_10_15_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14483\,
            in2 => \N__14474\,
            in3 => \N__18220\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14465\,
            in2 => \N__14456\,
            in3 => \N__18196\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14447\,
            in2 => \N__14441\,
            in3 => \N__18163\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14432\,
            in2 => \N__14426\,
            in3 => \N__18139\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16814\,
            in2 => \N__14597\,
            in3 => \N__18112\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14588\,
            in2 => \N__14579\,
            in3 => \N__18091\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14570\,
            in2 => \N__14561\,
            in3 => \N__18064\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__18400\,
            in1 => \N__16769\,
            in2 => \N__14552\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_10_16_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16490\,
            in2 => \N__14543\,
            in3 => \N__18376\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16808\,
            in2 => \N__14534\,
            in3 => \N__18355\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16763\,
            in2 => \N__14525\,
            in3 => \N__19520\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16727\,
            in2 => \N__14516\,
            in3 => \N__18331\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16451\,
            in2 => \N__14507\,
            in3 => \N__18310\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16298\,
            in2 => \N__14696\,
            in3 => \N__18289\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14687\,
            in2 => \N__14675\,
            in3 => \N__18268\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14666\,
            in2 => \N__14657\,
            in3 => \N__18478\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_10_17_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14648\,
            in2 => \N__14639\,
            in3 => \N__18457\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14630\,
            in2 => \N__14621\,
            in3 => \N__18436\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14612\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.target_time_12_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100010001000"
        )
    port map (
            in0 => \N__16603\,
            in1 => \N__17321\,
            in2 => \N__16440\,
            in3 => \N__16713\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21131\,
            ce => \N__15142\,
            sr => \N__20796\
        );

    \phase_controller_slave.stoper_hc.target_time_19_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16232\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21131\,
            ce => \N__15142\,
            sr => \N__20796\
        );

    \phase_controller_slave.stoper_hc.target_time_11_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100010001000"
        )
    port map (
            in0 => \N__16602\,
            in1 => \N__17282\,
            in2 => \N__16439\,
            in3 => \N__16712\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21131\,
            ce => \N__15142\,
            sr => \N__20796\
        );

    \phase_controller_slave.stoper_hc.target_time_7_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100010001000"
        )
    port map (
            in0 => \N__16604\,
            in1 => \N__16062\,
            in2 => \N__16441\,
            in3 => \N__16714\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21131\,
            ce => \N__15142\,
            sr => \N__20796\
        );

    \phase_controller_slave.stoper_hc.target_time_9_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111011001100"
        )
    port map (
            in0 => \N__16715\,
            in1 => \N__16801\,
            in2 => \N__17921\,
            in3 => \N__16428\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21131\,
            ce => \N__15142\,
            sr => \N__20796\
        );

    \phase_controller_slave.stoper_hc.target_time_10_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100010001000"
        )
    port map (
            in0 => \N__16601\,
            in1 => \N__16514\,
            in2 => \N__16438\,
            in3 => \N__16711\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21131\,
            ce => \N__15142\,
            sr => \N__20796\
        );

    \phase_controller_slave.stoper_hc.target_time_15_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__17920\,
            in1 => \N__16415\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21131\,
            ce => \N__15142\,
            sr => \N__20796\
        );

    \phase_controller_slave.stoper_hc.target_time_14_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__17916\,
            in1 => \N__16430\,
            in2 => \_gnd_net_\,
            in3 => \N__16484\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21126\,
            ce => \N__15143\,
            sr => \N__20802\
        );

    \phase_controller_slave.stoper_hc.target_time_16_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16265\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21126\,
            ce => \N__15143\,
            sr => \N__20802\
        );

    \phase_controller_slave.stoper_hc.target_time_17_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16199\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21126\,
            ce => \N__15143\,
            sr => \N__20802\
        );

    \phase_controller_slave.stoper_hc.target_time_18_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16165\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21126\,
            ce => \N__15143\,
            sr => \N__20802\
        );

    \phase_controller_slave.stoper_hc.target_time_13_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000011000000"
        )
    port map (
            in0 => \N__16716\,
            in1 => \N__16605\,
            in2 => \N__16756\,
            in3 => \N__16429\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21126\,
            ce => \N__15143\,
            sr => \N__20802\
        );

    \delay_measurement_inst.delay_tr_reg_ess_3_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__14989\,
            in1 => \N__19166\,
            in2 => \N__15283\,
            in3 => \N__14950\,
            lcout => measured_delay_tr_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21122\,
            ce => \N__16886\,
            sr => \N__17184\
        );

    \delay_measurement_inst.delay_tr_reg_esr_18_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__21676\,
            in1 => \N__20076\,
            in2 => \_gnd_net_\,
            in3 => \N__16984\,
            lcout => measured_delay_tr_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21122\,
            ce => \N__16886\,
            sr => \N__17184\
        );

    \delay_measurement_inst.delay_tr_reg_esr_4_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__14949\,
            in1 => \N__14990\,
            in2 => \N__19124\,
            in3 => \N__15272\,
            lcout => measured_delay_tr_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21122\,
            ce => \N__16886\,
            sr => \N__17184\
        );

    \delay_measurement_inst.delay_tr_reg_esr_2_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__14988\,
            in1 => \N__16999\,
            in2 => \N__15282\,
            in3 => \N__14948\,
            lcout => measured_delay_tr_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21122\,
            ce => \N__16886\,
            sr => \N__17184\
        );

    \delay_measurement_inst.delay_tr_reg_esr_10_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__19748\,
            in1 => \N__21680\,
            in2 => \_gnd_net_\,
            in3 => \N__15361\,
            lcout => measured_delay_tr_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21122\,
            ce => \N__16886\,
            sr => \N__17184\
        );

    \delay_measurement_inst.delay_tr_reg_esr_11_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__15362\,
            in1 => \N__21677\,
            in2 => \_gnd_net_\,
            in3 => \N__19702\,
            lcout => measured_delay_tr_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21122\,
            ce => \N__16886\,
            sr => \N__17184\
        );

    \delay_measurement_inst.delay_tr_reg_esr_13_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__21675\,
            in1 => \N__19612\,
            in2 => \_gnd_net_\,
            in3 => \N__15363\,
            lcout => measured_delay_tr_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21122\,
            ce => \N__16886\,
            sr => \N__17184\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIC9OF1_2_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000000"
        )
    port map (
            in0 => \N__17000\,
            in1 => \N__19165\,
            in2 => \N__19801\,
            in3 => \N__17114\,
            lcout => \delay_measurement_inst.delay_tr_timer.un1_reset_i_a2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110010"
        )
    port map (
            in0 => \N__20257\,
            in1 => \N__17104\,
            in2 => \N__19562\,
            in3 => \N__16976\,
            lcout => \delay_measurement_inst.N_132\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19658\,
            in1 => \N__19703\,
            in2 => \N__19613\,
            in3 => \N__19744\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_167\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIA9RL2_15_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__17103\,
            in1 => \N__21666\,
            in2 => \_gnd_net_\,
            in3 => \N__20258\,
            lcout => \delay_measurement_inst.N_139\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.tr_state_RNI5LDIC_0_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__15321\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17145\,
            lcout => \delay_measurement_inst.N_134_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17090\,
            in1 => \N__17120\,
            in2 => \N__19979\,
            in3 => \N__17084\,
            lcout => \delay_measurement_inst.N_201\,
            ltout => \delay_measurement_inst.N_201_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4T357_15_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__20256\,
            in1 => \_gnd_net_\,
            in2 => \N__15305\,
            in3 => \N__15301\,
            lcout => \delay_measurement_inst.N_170\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_1_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010001000100"
        )
    port map (
            in0 => \N__15244\,
            in1 => \N__18969\,
            in2 => \N__19504\,
            in3 => \N__21227\,
            lcout => \phase_controller_inst1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21112\,
            ce => 'H',
            sr => \N__20811\
        );

    \phase_controller_inst1.state_RNIR0JF_1_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18968\,
            in2 => \_gnd_net_\,
            in3 => \N__15243\,
            lcout => \phase_controller_inst1.T01_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.T12_LC_10_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010111000"
        )
    port map (
            in0 => \N__15763\,
            in1 => \N__15214\,
            in2 => \N__15166\,
            in3 => \N__15191\,
            lcout => \T12_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21103\,
            ce => 'H',
            sr => \N__20826\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_1_LC_10_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010000000101100"
        )
    port map (
            in0 => \N__15567\,
            in1 => \N__15889\,
            in2 => \N__15715\,
            in3 => \N__15938\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21103\,
            ce => 'H',
            sr => \N__20826\
        );

    \phase_controller_inst1.stoper_tr.time_passed_LC_10_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000111000000"
        )
    port map (
            in0 => \N__15937\,
            in1 => \N__15488\,
            in2 => \N__15767\,
            in3 => \N__15890\,
            lcout => \phase_controller_inst1.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21103\,
            ce => 'H',
            sr => \N__20826\
        );

    \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_10_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15626\,
            in2 => \_gnd_net_\,
            in3 => \N__15568\,
            lcout => \phase_controller_inst1.stoper_tr.N_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__15482\,
            in1 => \N__15460\,
            in2 => \_gnd_net_\,
            in3 => \N__17040\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_181_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.hc_prev_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15422\,
            lcout => \delay_measurement_inst.hc_prevZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21171\,
            ce => 'H',
            sr => \N__20761\
        );

    \delay_measurement_inst.hc_sync_1_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17054\,
            lcout => \delay_measurement_inst.hc_syncZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21171\,
            ce => 'H',
            sr => \N__20761\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI84NG1_15_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__15404\,
            in1 => \N__17797\,
            in2 => \_gnd_net_\,
            in3 => \N__18040\,
            lcout => \delay_measurement_inst.N_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto19_6_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16052\,
            in1 => \N__16467\,
            in2 => \N__16097\,
            in3 => \N__16790\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_hc_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15389\,
            in2 => \_gnd_net_\,
            in3 => \N__20893\,
            lcout => \delay_measurement_inst.stop_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21156\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto6_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010101010"
        )
    port map (
            in0 => \N__16836\,
            in1 => \N__17451\,
            in2 => \N__17408\,
            in3 => \N__15956\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un1_startlt8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto9_0_0_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010101010"
        )
    port map (
            in0 => \N__16468\,
            in1 => \N__16791\,
            in2 => \N__16109\,
            in3 => \N__16028\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlt15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto9_c_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__16789\,
            in1 => \N__16084\,
            in2 => \_gnd_net_\,
            in3 => \N__16051\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un1_startlto9_cZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto13_3_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__17313\,
            in1 => \N__17264\,
            in2 => \N__16031\,
            in3 => \N__15949\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto19_8_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__16260\,
            in1 => \N__16022\,
            in2 => \N__16194\,
            in3 => \N__15950\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_8\,
            ltout => \phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_start_0_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__16329\,
            in1 => \N__17879\,
            in2 => \N__15983\,
            in3 => \N__17217\,
            lcout => \phase_controller_inst1.stoper_hc.un3_start\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto5_1_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__16283\,
            in1 => \N__17345\,
            in2 => \_gnd_net_\,
            in3 => \N__15972\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto19_2_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16743\,
            in2 => \_gnd_net_\,
            in3 => \N__16506\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto19_4_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__17878\,
            in1 => \N__16226\,
            in2 => \_gnd_net_\,
            in3 => \N__16160\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto6_0_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__16835\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16284\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto6Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16259\,
            in1 => \N__16227\,
            in2 => \N__16193\,
            in3 => \N__16161\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2\,
            ltout => \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto19_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17880\,
            in2 => \N__16136\,
            in3 => \N__16642\,
            lcout => \phase_controller_inst1.stoper_hc.un1_start\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__19302\,
            in1 => \N__19456\,
            in2 => \N__18176\,
            in3 => \N__21371\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21144\,
            ce => 'H',
            sr => \N__20776\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__21367\,
            in1 => \N__19305\,
            in2 => \N__19461\,
            in3 => \N__18152\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21144\,
            ce => 'H',
            sr => \N__20776\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__19303\,
            in1 => \N__19457\,
            in2 => \N__18128\,
            in3 => \N__21372\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21144\,
            ce => 'H',
            sr => \N__20776\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__21368\,
            in1 => \N__19306\,
            in2 => \N__19462\,
            in3 => \N__18101\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21144\,
            ce => 'H',
            sr => \N__20776\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__19304\,
            in1 => \N__19458\,
            in2 => \N__18080\,
            in3 => \N__21373\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21144\,
            ce => 'H',
            sr => \N__20776\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__21369\,
            in1 => \N__19307\,
            in2 => \N__19463\,
            in3 => \N__18053\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21144\,
            ce => 'H',
            sr => \N__20776\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__19301\,
            in1 => \N__19455\,
            in2 => \N__18209\,
            in3 => \N__21370\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21144\,
            ce => 'H',
            sr => \N__20776\
        );

    \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111101110111011"
        )
    port map (
            in0 => \N__16847\,
            in1 => \N__16579\,
            in2 => \N__16412\,
            in3 => \N__16675\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21141\,
            ce => \N__18765\,
            sr => \N__20780\
        );

    \phase_controller_inst1.stoper_hc.target_time_11_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__16677\,
            in1 => \N__16371\,
            in2 => \N__16607\,
            in3 => \N__17278\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21141\,
            ce => \N__18765\,
            sr => \N__20780\
        );

    \phase_controller_inst1.stoper_hc.target_time_9_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110011101100"
        )
    port map (
            in0 => \N__17915\,
            in1 => \N__16802\,
            in2 => \N__16414\,
            in3 => \N__16680\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21141\,
            ce => \N__18765\,
            sr => \N__20780\
        );

    \phase_controller_inst1.stoper_hc.target_time_12_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__16678\,
            in1 => \N__16372\,
            in2 => \N__16608\,
            in3 => \N__17320\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21141\,
            ce => \N__18765\,
            sr => \N__20780\
        );

    \phase_controller_inst1.stoper_hc.target_time_13_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000011000000"
        )
    port map (
            in0 => \N__16373\,
            in1 => \N__16580\,
            in2 => \N__16757\,
            in3 => \N__16679\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21141\,
            ce => \N__18765\,
            sr => \N__20780\
        );

    \phase_controller_inst1.stoper_hc.target_time_10_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__16676\,
            in1 => \N__16370\,
            in2 => \N__16606\,
            in3 => \N__16513\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21141\,
            ce => \N__18765\,
            sr => \N__20780\
        );

    \phase_controller_inst1.stoper_hc.target_time_14_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17913\,
            in2 => \N__16413\,
            in3 => \N__16480\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21141\,
            ce => \N__18765\,
            sr => \N__20780\
        );

    \phase_controller_inst1.stoper_hc.target_time_15_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__17914\,
            in1 => \N__16366\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21141\,
            ce => \N__18765\,
            sr => \N__20780\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_0_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__21249\,
            in1 => \N__19284\,
            in2 => \N__19433\,
            in3 => \N__21344\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21135\,
            ce => 'H',
            sr => \N__20781\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__21338\,
            in1 => \N__18248\,
            in2 => \_gnd_net_\,
            in3 => \N__21248\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__19381\,
            in1 => \N__19283\,
            in2 => \N__16850\,
            in3 => \N__21343\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21135\,
            ce => 'H',
            sr => \N__20781\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21311\,
            in2 => \_gnd_net_\,
            in3 => \N__21246\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_1_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010111000000"
        )
    port map (
            in0 => \N__21250\,
            in1 => \N__19285\,
            in2 => \N__19434\,
            in3 => \N__21345\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21135\,
            ce => 'H',
            sr => \N__20781\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIGEUB_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21312\,
            in2 => \_gnd_net_\,
            in3 => \N__21247\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIGEUBZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__19281\,
            in1 => \N__21339\,
            in2 => \N__19432\,
            in3 => \N__18365\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21135\,
            ce => 'H',
            sr => \N__20781\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__19282\,
            in1 => \N__19382\,
            in2 => \N__21374\,
            in3 => \N__18344\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21135\,
            ce => 'H',
            sr => \N__20781\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__21346\,
            in1 => \N__19277\,
            in2 => \N__19435\,
            in3 => \N__18320\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21132\,
            ce => 'H',
            sr => \N__20785\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__19273\,
            in1 => \N__19392\,
            in2 => \N__21387\,
            in3 => \N__18299\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21132\,
            ce => 'H',
            sr => \N__20785\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__21347\,
            in1 => \N__19278\,
            in2 => \N__19436\,
            in3 => \N__18278\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21132\,
            ce => 'H',
            sr => \N__20785\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__19274\,
            in1 => \N__19393\,
            in2 => \N__21388\,
            in3 => \N__18257\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21132\,
            ce => 'H',
            sr => \N__20785\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__21348\,
            in1 => \N__19279\,
            in2 => \N__19437\,
            in3 => \N__18467\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21132\,
            ce => 'H',
            sr => \N__20785\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__19275\,
            in1 => \N__19394\,
            in2 => \N__21389\,
            in3 => \N__18446\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21132\,
            ce => 'H',
            sr => \N__20785\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__21349\,
            in1 => \N__19280\,
            in2 => \N__19438\,
            in3 => \N__18422\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21132\,
            ce => 'H',
            sr => \N__20785\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011010000"
        )
    port map (
            in0 => \N__19276\,
            in1 => \N__21350\,
            in2 => \N__18389\,
            in3 => \N__19407\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21132\,
            ce => 'H',
            sr => \N__20785\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19184\,
            lcout => \delay_measurement_inst.elapsed_time_tr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21123\,
            ce => \N__21593\,
            sr => \N__20797\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19142\,
            lcout => \delay_measurement_inst.elapsed_time_tr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21123\,
            ce => \N__21593\,
            sr => \N__20797\
        );

    \delay_measurement_inst.delay_tr_reg_esr_19_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__21681\,
            in1 => \N__16983\,
            in2 => \_gnd_net_\,
            in3 => \N__20027\,
            lcout => measured_delay_tr_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21117\,
            ce => \N__16887\,
            sr => \N__17183\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19943\,
            in1 => \N__20534\,
            in2 => \N__20570\,
            in3 => \N__19910\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_0_o2_0_7_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFD841_4_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20131\,
            in1 => \N__19072\,
            in2 => \N__20026\,
            in3 => \N__19120\,
            lcout => \delay_measurement_inst.delay_tr_timer.un1_reset_i_a2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__20187\,
            in1 => \N__20022\,
            in2 => \N__20084\,
            in3 => \N__20132\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_127\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20432\,
            in1 => \N__20465\,
            in2 => \N__20396\,
            in3 => \N__20498\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_0_o2_0_6_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20294\,
            in2 => \_gnd_net_\,
            in3 => \N__20342\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_0_o2_0_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_11_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17078\,
            lcout => \GB_BUFFER_clk_12mhz_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_HC2_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18863\,
            lcout => delay_hc_d2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21176\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.hc_sync_0_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17060\,
            lcout => \delay_measurement_inst.hc_syncZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21169\,
            ce => 'H',
            sr => \N__20758\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17048\,
            lcout => \delay_measurement_inst.delay_tr_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_esr_15_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000001100"
        )
    port map (
            in0 => \N__17820\,
            in1 => \N__18044\,
            in2 => \N__17995\,
            in3 => \N__17978\,
            lcout => measured_delay_hc_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21148\,
            ce => \N__17690\,
            sr => \N__17660\
        );

    \delay_measurement_inst.delay_hc_reg_esr_12_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001000100"
        )
    port map (
            in0 => \N__17717\,
            in1 => \N__17858\,
            in2 => \_gnd_net_\,
            in3 => \N__17819\,
            lcout => measured_delay_hc_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21148\,
            ce => \N__17690\,
            sr => \N__17660\
        );

    \delay_measurement_inst.delay_hc_reg_esr_11_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__17818\,
            in1 => \N__17738\,
            in2 => \_gnd_net_\,
            in3 => \N__17716\,
            lcout => measured_delay_hc_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21148\,
            ce => \N__17690\,
            sr => \N__17660\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18804\,
            lcout => \delay_measurement_inst.delay_hc_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__18805\,
            in1 => \N__18847\,
            in2 => \_gnd_net_\,
            in3 => \N__18822\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_179_i_g\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto6_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__17452\,
            in1 => \N__17414\,
            in2 => \N__17407\,
            in3 => \N__17355\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un2_startlt19_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto19_9_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__17327\,
            in1 => \N__17309\,
            in2 => \N__17285\,
            in3 => \N__17265\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D2_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17201\,
            lcout => \il_max_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21140\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18247\,
            in2 => \N__18230\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_15_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18221\,
            in2 => \_gnd_net_\,
            in3 => \N__18200\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18197\,
            in2 => \N__18185\,
            in3 => \N__18167\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18164\,
            in2 => \_gnd_net_\,
            in3 => \N__18146\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18143\,
            in3 => \N__18119\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18116\,
            in3 => \N__18095\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18092\,
            in2 => \_gnd_net_\,
            in3 => \N__18071\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18068\,
            in3 => \N__18047\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18401\,
            in2 => \_gnd_net_\,
            in3 => \N__18380\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_12_16_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18377\,
            in2 => \_gnd_net_\,
            in3 => \N__18359\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18356\,
            in2 => \_gnd_net_\,
            in3 => \N__18338\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19519\,
            in2 => \_gnd_net_\,
            in3 => \N__18335\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18332\,
            in2 => \_gnd_net_\,
            in3 => \N__18314\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18311\,
            in2 => \_gnd_net_\,
            in3 => \N__18293\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18290\,
            in2 => \_gnd_net_\,
            in3 => \N__18272\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18269\,
            in2 => \_gnd_net_\,
            in3 => \N__18251\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18479\,
            in2 => \_gnd_net_\,
            in3 => \N__18461\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_12_17_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18458\,
            in2 => \_gnd_net_\,
            in3 => \N__18440\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18437\,
            in2 => \_gnd_net_\,
            in3 => \N__18425\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.counter_0_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18705\,
            in1 => \N__19182\,
            in2 => \_gnd_net_\,
            in3 => \N__18416\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_12_18_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            clk => \N__21121\,
            ce => \N__18593\,
            sr => \N__20786\
        );

    \delay_measurement_inst.delay_tr_timer.counter_1_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18700\,
            in1 => \N__19140\,
            in2 => \_gnd_net_\,
            in3 => \N__18413\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            clk => \N__21121\,
            ce => \N__18593\,
            sr => \N__20786\
        );

    \delay_measurement_inst.delay_tr_timer.counter_2_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18706\,
            in1 => \N__19092\,
            in2 => \_gnd_net_\,
            in3 => \N__18410\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            clk => \N__21121\,
            ce => \N__18593\,
            sr => \N__20786\
        );

    \delay_measurement_inst.delay_tr_timer.counter_3_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18701\,
            in1 => \N__19044\,
            in2 => \_gnd_net_\,
            in3 => \N__18407\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            clk => \N__21121\,
            ce => \N__18593\,
            sr => \N__20786\
        );

    \delay_measurement_inst.delay_tr_timer.counter_4_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18707\,
            in1 => \N__18999\,
            in2 => \_gnd_net_\,
            in3 => \N__18404\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            clk => \N__21121\,
            ce => \N__18593\,
            sr => \N__20786\
        );

    \delay_measurement_inst.delay_tr_timer.counter_5_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18702\,
            in1 => \N__19869\,
            in2 => \_gnd_net_\,
            in3 => \N__18506\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            clk => \N__21121\,
            ce => \N__18593\,
            sr => \N__20786\
        );

    \delay_measurement_inst.delay_tr_timer.counter_6_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18704\,
            in1 => \N__19821\,
            in2 => \_gnd_net_\,
            in3 => \N__18503\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            clk => \N__21121\,
            ce => \N__18593\,
            sr => \N__20786\
        );

    \delay_measurement_inst.delay_tr_timer.counter_7_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18703\,
            in1 => \N__19767\,
            in2 => \_gnd_net_\,
            in3 => \N__18500\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            clk => \N__21121\,
            ce => \N__18593\,
            sr => \N__20786\
        );

    \delay_measurement_inst.delay_tr_timer.counter_8_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18699\,
            in1 => \N__19722\,
            in2 => \_gnd_net_\,
            in3 => \N__18497\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_12_19_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            clk => \N__21116\,
            ce => \N__18594\,
            sr => \N__20791\
        );

    \delay_measurement_inst.delay_tr_timer.counter_9_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18711\,
            in1 => \N__19677\,
            in2 => \_gnd_net_\,
            in3 => \N__18494\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            clk => \N__21116\,
            ce => \N__18594\,
            sr => \N__20791\
        );

    \delay_measurement_inst.delay_tr_timer.counter_10_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18696\,
            in1 => \N__19632\,
            in2 => \_gnd_net_\,
            in3 => \N__18491\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            clk => \N__21116\,
            ce => \N__18594\,
            sr => \N__20791\
        );

    \delay_measurement_inst.delay_tr_timer.counter_11_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18708\,
            in1 => \N__19581\,
            in2 => \_gnd_net_\,
            in3 => \N__18488\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            clk => \N__21116\,
            ce => \N__18594\,
            sr => \N__20791\
        );

    \delay_measurement_inst.delay_tr_timer.counter_12_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18697\,
            in1 => \N__20280\,
            in2 => \_gnd_net_\,
            in3 => \N__18485\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            clk => \N__21116\,
            ce => \N__18594\,
            sr => \N__20791\
        );

    \delay_measurement_inst.delay_tr_timer.counter_13_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18709\,
            in1 => \N__20208\,
            in2 => \_gnd_net_\,
            in3 => \N__18482\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            clk => \N__21116\,
            ce => \N__18594\,
            sr => \N__20791\
        );

    \delay_measurement_inst.delay_tr_timer.counter_14_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18698\,
            in1 => \N__20151\,
            in2 => \_gnd_net_\,
            in3 => \N__18536\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            clk => \N__21116\,
            ce => \N__18594\,
            sr => \N__20791\
        );

    \delay_measurement_inst.delay_tr_timer.counter_15_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18710\,
            in1 => \N__20103\,
            in2 => \_gnd_net_\,
            in3 => \N__18533\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            clk => \N__21116\,
            ce => \N__18594\,
            sr => \N__20791\
        );

    \delay_measurement_inst.delay_tr_timer.counter_16_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18714\,
            in1 => \N__20046\,
            in2 => \_gnd_net_\,
            in3 => \N__18530\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_12_20_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            clk => \N__21111\,
            ce => \N__18595\,
            sr => \N__20798\
        );

    \delay_measurement_inst.delay_tr_timer.counter_17_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18718\,
            in1 => \N__19998\,
            in2 => \_gnd_net_\,
            in3 => \N__18527\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            clk => \N__21111\,
            ce => \N__18595\,
            sr => \N__20798\
        );

    \delay_measurement_inst.delay_tr_timer.counter_18_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18715\,
            in1 => \N__19962\,
            in2 => \_gnd_net_\,
            in3 => \N__18524\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            clk => \N__21111\,
            ce => \N__18595\,
            sr => \N__20798\
        );

    \delay_measurement_inst.delay_tr_timer.counter_19_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18719\,
            in1 => \N__19929\,
            in2 => \_gnd_net_\,
            in3 => \N__18521\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            clk => \N__21111\,
            ce => \N__18595\,
            sr => \N__20798\
        );

    \delay_measurement_inst.delay_tr_timer.counter_20_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18716\,
            in1 => \N__20589\,
            in2 => \_gnd_net_\,
            in3 => \N__18518\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            clk => \N__21111\,
            ce => \N__18595\,
            sr => \N__20798\
        );

    \delay_measurement_inst.delay_tr_timer.counter_21_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18720\,
            in1 => \N__20553\,
            in2 => \_gnd_net_\,
            in3 => \N__18515\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            clk => \N__21111\,
            ce => \N__18595\,
            sr => \N__20798\
        );

    \delay_measurement_inst.delay_tr_timer.counter_22_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18717\,
            in1 => \N__20517\,
            in2 => \_gnd_net_\,
            in3 => \N__18512\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            clk => \N__21111\,
            ce => \N__18595\,
            sr => \N__20798\
        );

    \delay_measurement_inst.delay_tr_timer.counter_23_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18721\,
            in1 => \N__20484\,
            in2 => \_gnd_net_\,
            in3 => \N__18509\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            clk => \N__21111\,
            ce => \N__18595\,
            sr => \N__20798\
        );

    \delay_measurement_inst.delay_tr_timer.counter_24_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18722\,
            in1 => \N__20451\,
            in2 => \_gnd_net_\,
            in3 => \N__18740\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_12_21_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            clk => \N__21107\,
            ce => \N__18596\,
            sr => \N__20803\
        );

    \delay_measurement_inst.delay_tr_timer.counter_25_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18712\,
            in1 => \N__20415\,
            in2 => \_gnd_net_\,
            in3 => \N__18737\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            clk => \N__21107\,
            ce => \N__18596\,
            sr => \N__20803\
        );

    \delay_measurement_inst.delay_tr_timer.counter_26_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18723\,
            in1 => \N__20376\,
            in2 => \_gnd_net_\,
            in3 => \N__18734\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            clk => \N__21107\,
            ce => \N__18596\,
            sr => \N__20803\
        );

    \delay_measurement_inst.delay_tr_timer.counter_27_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18713\,
            in1 => \N__20328\,
            in2 => \_gnd_net_\,
            in3 => \N__18731\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            clk => \N__21107\,
            ce => \N__18596\,
            sr => \N__20803\
        );

    \delay_measurement_inst.delay_tr_timer.counter_28_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18724\,
            in1 => \N__20356\,
            in2 => \_gnd_net_\,
            in3 => \N__18728\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_28\,
            clk => \N__21107\,
            ce => \N__18596\,
            sr => \N__20803\
        );

    \delay_measurement_inst.delay_tr_timer.counter_29_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__20308\,
            in1 => \N__18725\,
            in2 => \_gnd_net_\,
            in3 => \N__18599\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21107\,
            ce => \N__18596\,
            sr => \N__20803\
        );

    \phase_controller_inst1.state_2_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__18578\,
            in1 => \N__19484\,
            in2 => \N__18937\,
            in3 => \N__21226\,
            lcout => \phase_controller_inst1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21104\,
            ce => 'H',
            sr => \N__20807\
        );

    \phase_controller_inst1.start_timer_hc_RNO_1_LC_12_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18920\,
            in2 => \_gnd_net_\,
            in3 => \N__18576\,
            lcout => \phase_controller_inst1.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_3_LC_12_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110111010"
        )
    port map (
            in0 => \N__21440\,
            in1 => \N__18577\,
            in2 => \N__18936\,
            in3 => \N__18554\,
            lcout => \phase_controller_inst1.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21102\,
            ce => 'H',
            sr => \N__20812\
        );

    \phase_controller_inst1.S2_LC_12_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18980\,
            lcout => s2_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21101\,
            ce => 'H',
            sr => \N__20818\
        );

    \phase_controller_inst1.S1_LC_12_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18938\,
            lcout => s1_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21099\,
            ce => 'H',
            sr => \N__20836\
        );

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20899\,
            lcout => \pll_inst.red_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_HC1_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__18878\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => delay_hc_d1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21184\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.tr_sync_0_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21400\,
            lcout => \delay_measurement_inst.tr_syncZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21172\,
            ce => 'H',
            sr => \N__20759\
        );

    \delay_measurement_inst.delay_hc_timer.running_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__18848\,
            in1 => \N__18830\,
            in2 => \_gnd_net_\,
            in3 => \N__18806\,
            lcout => \delay_measurement_inst.delay_hc_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21150\,
            ce => 'H',
            sr => \N__20762\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18829\,
            in2 => \_gnd_net_\,
            in3 => \N__18803\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_178_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_1_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__19445\,
            in1 => \N__19238\,
            in2 => \_gnd_net_\,
            in3 => \N__21375\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_state_RNITN7VZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__19239\,
            in1 => \N__21376\,
            in2 => \N__19460\,
            in3 => \N__19526\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21136\,
            ce => 'H',
            sr => \N__20777\
        );

    \phase_controller_inst1.start_timer_hc_RNO_0_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19500\,
            in2 => \_gnd_net_\,
            in3 => \N__21210\,
            lcout => \phase_controller_inst1.N_112\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19459\,
            in2 => \_gnd_net_\,
            in3 => \N__19223\,
            lcout => \phase_controller_inst1.stoper_hc.N_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__21480\,
            in1 => \N__19325\,
            in2 => \N__19272\,
            in3 => \N__19313\,
            lcout => \phase_controller_inst1.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21127\,
            ce => 'H',
            sr => \N__20782\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19183\,
            in2 => \N__19094\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.elapsed_time_tr_3\,
            ltout => OPEN,
            carryin => \bfn_13_19_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__21124\,
            ce => \N__21596\,
            sr => \N__20787\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19141\,
            in2 => \N__19046\,
            in3 => \N__19097\,
            lcout => \delay_measurement_inst.elapsed_time_tr_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__21124\,
            ce => \N__21596\,
            sr => \N__20787\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19093\,
            in2 => \N__19001\,
            in3 => \N__19049\,
            lcout => \delay_measurement_inst.elapsed_time_tr_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__21124\,
            ce => \N__21596\,
            sr => \N__20787\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19045\,
            in2 => \N__19871\,
            in3 => \N__19004\,
            lcout => \delay_measurement_inst.elapsed_time_tr_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__21124\,
            ce => \N__21596\,
            sr => \N__20787\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19000\,
            in2 => \N__19823\,
            in3 => \N__19874\,
            lcout => \delay_measurement_inst.elapsed_time_tr_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__21124\,
            ce => \N__21596\,
            sr => \N__20787\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19870\,
            in2 => \N__19769\,
            in3 => \N__19826\,
            lcout => \delay_measurement_inst.elapsed_time_tr_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__21124\,
            ce => \N__21596\,
            sr => \N__20787\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19822\,
            in2 => \N__19724\,
            in3 => \N__19772\,
            lcout => \delay_measurement_inst.elapsed_time_tr_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__21124\,
            ce => \N__21596\,
            sr => \N__20787\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19768\,
            in2 => \N__19679\,
            in3 => \N__19727\,
            lcout => \delay_measurement_inst.elapsed_time_tr_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__21124\,
            ce => \N__21596\,
            sr => \N__20787\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19723\,
            in2 => \N__19634\,
            in3 => \N__19682\,
            lcout => \delay_measurement_inst.elapsed_time_tr_11\,
            ltout => OPEN,
            carryin => \bfn_13_20_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__21118\,
            ce => \N__21595\,
            sr => \N__20792\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19678\,
            in2 => \N__19583\,
            in3 => \N__19637\,
            lcout => \delay_measurement_inst.elapsed_time_tr_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__21118\,
            ce => \N__21595\,
            sr => \N__20792\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19633\,
            in2 => \N__20282\,
            in3 => \N__19586\,
            lcout => \delay_measurement_inst.elapsed_time_tr_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__21118\,
            ce => \N__21595\,
            sr => \N__20792\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19582\,
            in2 => \N__20210\,
            in3 => \N__19529\,
            lcout => \delay_measurement_inst.elapsed_time_tr_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__21118\,
            ce => \N__21595\,
            sr => \N__20792\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20281\,
            in2 => \N__20153\,
            in3 => \N__20213\,
            lcout => \delay_measurement_inst.elapsed_time_tr_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__21118\,
            ce => \N__21595\,
            sr => \N__20792\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20209\,
            in2 => \N__20105\,
            in3 => \N__20156\,
            lcout => \delay_measurement_inst.elapsed_time_tr_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__21118\,
            ce => \N__21595\,
            sr => \N__20792\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20152\,
            in2 => \N__20048\,
            in3 => \N__20108\,
            lcout => \delay_measurement_inst.elapsed_time_tr_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__21118\,
            ce => \N__21595\,
            sr => \N__20792\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20104\,
            in2 => \N__20000\,
            in3 => \N__20051\,
            lcout => \delay_measurement_inst.elapsed_time_tr_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__21118\,
            ce => \N__21595\,
            sr => \N__20792\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20047\,
            in2 => \N__19964\,
            in3 => \N__20003\,
            lcout => \delay_measurement_inst.elapsed_time_tr_19\,
            ltout => OPEN,
            carryin => \bfn_13_21_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__21113\,
            ce => \N__21594\,
            sr => \N__20799\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19999\,
            in2 => \N__19931\,
            in3 => \N__19967\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__21113\,
            ce => \N__21594\,
            sr => \N__20799\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19963\,
            in2 => \N__20591\,
            in3 => \N__19934\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__21113\,
            ce => \N__21594\,
            sr => \N__20799\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19930\,
            in2 => \N__20555\,
            in3 => \N__19901\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__21113\,
            ce => \N__21594\,
            sr => \N__20799\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20590\,
            in2 => \N__20519\,
            in3 => \N__20558\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__21113\,
            ce => \N__21594\,
            sr => \N__20799\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20554\,
            in2 => \N__20486\,
            in3 => \N__20522\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__21113\,
            ce => \N__21594\,
            sr => \N__20799\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20518\,
            in2 => \N__20453\,
            in3 => \N__20489\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__21113\,
            ce => \N__21594\,
            sr => \N__20799\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_13_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20485\,
            in2 => \N__20417\,
            in3 => \N__20456\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__21113\,
            ce => \N__21594\,
            sr => \N__20799\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20452\,
            in2 => \N__20378\,
            in3 => \N__20420\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\,
            ltout => OPEN,
            carryin => \bfn_13_22_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__21108\,
            ce => \N__21592\,
            sr => \N__20804\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20416\,
            in2 => \N__20330\,
            in3 => \N__20381\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__21108\,
            ce => \N__21592\,
            sr => \N__20804\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20377\,
            in2 => \N__20357\,
            in3 => \N__20333\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__21108\,
            ce => \N__21592\,
            sr => \N__20804\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20329\,
            in2 => \N__20309\,
            in3 => \N__20285\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__21108\,
            ce => \N__21592\,
            sr => \N__20804\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21686\,
            lcout => \delay_measurement_inst.elapsed_time_tr_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21108\,
            ce => \N__21592\,
            sr => \N__20804\
        );

    \phase_controller_inst1.state_4_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21530\,
            in2 => \_gnd_net_\,
            in3 => \N__21464\,
            lcout => \phase_controller_inst1.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21105\,
            ce => 'H',
            sr => \N__20808\
        );

    \phase_controller_inst1.state_RNO_0_3_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21554\,
            in2 => \_gnd_net_\,
            in3 => \N__21463\,
            lcout => \phase_controller_inst1.N_110\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_TR1_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21434\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => delay_tr_d1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21188\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_TR2_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21422\,
            lcout => \T23_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__21214\,
            in1 => \N__21377\,
            in2 => \N__21263\,
            in3 => \N__21254\,
            lcout => \phase_controller_inst1.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21137\,
            ce => 'H',
            sr => \N__20778\
        );
end \INTERFACE\;
