-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Mar 2 2025 23:51:14

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MAIN" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MAIN
entity MAIN is
port (
    start_stop : in std_logic;
    s2_phy : out std_logic;
    T23 : out std_logic;
    s3_phy : out std_logic;
    il_min_comp2 : in std_logic;
    il_max_comp1 : in std_logic;
    s1_phy : out std_logic;
    reset : in std_logic;
    il_min_comp1 : in std_logic;
    delay_tr_input : in std_logic;
    T45 : out std_logic;
    T12 : out std_logic;
    s4_phy : out std_logic;
    rgb_g : out std_logic;
    T01 : out std_logic;
    rgb_r : out std_logic;
    rgb_b : out std_logic;
    pwm_output : out std_logic;
    il_max_comp2 : in std_logic;
    delay_hc_input : in std_logic);
end MAIN;

-- Architecture of MAIN
-- View name is \INTERFACE\
architecture \INTERFACE\ of MAIN is

signal \N__48452\ : std_logic;
signal \N__48451\ : std_logic;
signal \N__48450\ : std_logic;
signal \N__48441\ : std_logic;
signal \N__48440\ : std_logic;
signal \N__48439\ : std_logic;
signal \N__48432\ : std_logic;
signal \N__48431\ : std_logic;
signal \N__48430\ : std_logic;
signal \N__48423\ : std_logic;
signal \N__48422\ : std_logic;
signal \N__48421\ : std_logic;
signal \N__48414\ : std_logic;
signal \N__48413\ : std_logic;
signal \N__48412\ : std_logic;
signal \N__48405\ : std_logic;
signal \N__48404\ : std_logic;
signal \N__48403\ : std_logic;
signal \N__48396\ : std_logic;
signal \N__48395\ : std_logic;
signal \N__48394\ : std_logic;
signal \N__48387\ : std_logic;
signal \N__48386\ : std_logic;
signal \N__48385\ : std_logic;
signal \N__48378\ : std_logic;
signal \N__48377\ : std_logic;
signal \N__48376\ : std_logic;
signal \N__48369\ : std_logic;
signal \N__48368\ : std_logic;
signal \N__48367\ : std_logic;
signal \N__48360\ : std_logic;
signal \N__48359\ : std_logic;
signal \N__48358\ : std_logic;
signal \N__48351\ : std_logic;
signal \N__48350\ : std_logic;
signal \N__48349\ : std_logic;
signal \N__48342\ : std_logic;
signal \N__48341\ : std_logic;
signal \N__48340\ : std_logic;
signal \N__48333\ : std_logic;
signal \N__48332\ : std_logic;
signal \N__48331\ : std_logic;
signal \N__48324\ : std_logic;
signal \N__48323\ : std_logic;
signal \N__48322\ : std_logic;
signal \N__48315\ : std_logic;
signal \N__48314\ : std_logic;
signal \N__48313\ : std_logic;
signal \N__48306\ : std_logic;
signal \N__48305\ : std_logic;
signal \N__48304\ : std_logic;
signal \N__48287\ : std_logic;
signal \N__48286\ : std_logic;
signal \N__48285\ : std_logic;
signal \N__48284\ : std_logic;
signal \N__48281\ : std_logic;
signal \N__48278\ : std_logic;
signal \N__48275\ : std_logic;
signal \N__48272\ : std_logic;
signal \N__48269\ : std_logic;
signal \N__48266\ : std_logic;
signal \N__48263\ : std_logic;
signal \N__48260\ : std_logic;
signal \N__48257\ : std_logic;
signal \N__48254\ : std_logic;
signal \N__48251\ : std_logic;
signal \N__48248\ : std_logic;
signal \N__48245\ : std_logic;
signal \N__48242\ : std_logic;
signal \N__48239\ : std_logic;
signal \N__48236\ : std_logic;
signal \N__48227\ : std_logic;
signal \N__48226\ : std_logic;
signal \N__48223\ : std_logic;
signal \N__48222\ : std_logic;
signal \N__48219\ : std_logic;
signal \N__48216\ : std_logic;
signal \N__48213\ : std_logic;
signal \N__48206\ : std_logic;
signal \N__48205\ : std_logic;
signal \N__48204\ : std_logic;
signal \N__48203\ : std_logic;
signal \N__48202\ : std_logic;
signal \N__48201\ : std_logic;
signal \N__48200\ : std_logic;
signal \N__48199\ : std_logic;
signal \N__48198\ : std_logic;
signal \N__48197\ : std_logic;
signal \N__48196\ : std_logic;
signal \N__48195\ : std_logic;
signal \N__48194\ : std_logic;
signal \N__48193\ : std_logic;
signal \N__48190\ : std_logic;
signal \N__48189\ : std_logic;
signal \N__48188\ : std_logic;
signal \N__48187\ : std_logic;
signal \N__48186\ : std_logic;
signal \N__48185\ : std_logic;
signal \N__48184\ : std_logic;
signal \N__48183\ : std_logic;
signal \N__48182\ : std_logic;
signal \N__48181\ : std_logic;
signal \N__48180\ : std_logic;
signal \N__48179\ : std_logic;
signal \N__48178\ : std_logic;
signal \N__48177\ : std_logic;
signal \N__48176\ : std_logic;
signal \N__48173\ : std_logic;
signal \N__48170\ : std_logic;
signal \N__48169\ : std_logic;
signal \N__48160\ : std_logic;
signal \N__48155\ : std_logic;
signal \N__48154\ : std_logic;
signal \N__48153\ : std_logic;
signal \N__48152\ : std_logic;
signal \N__48151\ : std_logic;
signal \N__48150\ : std_logic;
signal \N__48149\ : std_logic;
signal \N__48148\ : std_logic;
signal \N__48147\ : std_logic;
signal \N__48146\ : std_logic;
signal \N__48145\ : std_logic;
signal \N__48144\ : std_logic;
signal \N__48133\ : std_logic;
signal \N__48132\ : std_logic;
signal \N__48131\ : std_logic;
signal \N__48130\ : std_logic;
signal \N__48129\ : std_logic;
signal \N__48118\ : std_logic;
signal \N__48117\ : std_logic;
signal \N__48116\ : std_logic;
signal \N__48105\ : std_logic;
signal \N__48102\ : std_logic;
signal \N__48101\ : std_logic;
signal \N__48100\ : std_logic;
signal \N__48099\ : std_logic;
signal \N__48098\ : std_logic;
signal \N__48097\ : std_logic;
signal \N__48096\ : std_logic;
signal \N__48095\ : std_logic;
signal \N__48092\ : std_logic;
signal \N__48091\ : std_logic;
signal \N__48090\ : std_logic;
signal \N__48089\ : std_logic;
signal \N__48088\ : std_logic;
signal \N__48087\ : std_logic;
signal \N__48080\ : std_logic;
signal \N__48073\ : std_logic;
signal \N__48068\ : std_logic;
signal \N__48063\ : std_logic;
signal \N__48060\ : std_logic;
signal \N__48057\ : std_logic;
signal \N__48052\ : std_logic;
signal \N__48051\ : std_logic;
signal \N__48042\ : std_logic;
signal \N__48039\ : std_logic;
signal \N__48036\ : std_logic;
signal \N__48027\ : std_logic;
signal \N__48026\ : std_logic;
signal \N__48025\ : std_logic;
signal \N__48024\ : std_logic;
signal \N__48023\ : std_logic;
signal \N__48022\ : std_logic;
signal \N__48021\ : std_logic;
signal \N__48020\ : std_logic;
signal \N__48019\ : std_logic;
signal \N__48016\ : std_logic;
signal \N__48011\ : std_logic;
signal \N__48010\ : std_logic;
signal \N__48009\ : std_logic;
signal \N__48008\ : std_logic;
signal \N__48007\ : std_logic;
signal \N__48006\ : std_logic;
signal \N__48005\ : std_logic;
signal \N__48004\ : std_logic;
signal \N__48003\ : std_logic;
signal \N__48002\ : std_logic;
signal \N__48001\ : std_logic;
signal \N__48000\ : std_logic;
signal \N__47999\ : std_logic;
signal \N__47998\ : std_logic;
signal \N__47997\ : std_logic;
signal \N__47996\ : std_logic;
signal \N__47995\ : std_logic;
signal \N__47992\ : std_logic;
signal \N__47989\ : std_logic;
signal \N__47988\ : std_logic;
signal \N__47987\ : std_logic;
signal \N__47986\ : std_logic;
signal \N__47985\ : std_logic;
signal \N__47984\ : std_logic;
signal \N__47983\ : std_logic;
signal \N__47982\ : std_logic;
signal \N__47981\ : std_logic;
signal \N__47980\ : std_logic;
signal \N__47971\ : std_logic;
signal \N__47960\ : std_logic;
signal \N__47951\ : std_logic;
signal \N__47936\ : std_logic;
signal \N__47933\ : std_logic;
signal \N__47928\ : std_logic;
signal \N__47925\ : std_logic;
signal \N__47922\ : std_logic;
signal \N__47917\ : std_logic;
signal \N__47910\ : std_logic;
signal \N__47903\ : std_logic;
signal \N__47898\ : std_logic;
signal \N__47895\ : std_logic;
signal \N__47886\ : std_logic;
signal \N__47879\ : std_logic;
signal \N__47870\ : std_logic;
signal \N__47861\ : std_logic;
signal \N__47856\ : std_logic;
signal \N__47853\ : std_logic;
signal \N__47848\ : std_logic;
signal \N__47839\ : std_logic;
signal \N__47834\ : std_logic;
signal \N__47827\ : std_logic;
signal \N__47824\ : std_logic;
signal \N__47813\ : std_logic;
signal \N__47806\ : std_logic;
signal \N__47777\ : std_logic;
signal \N__47776\ : std_logic;
signal \N__47775\ : std_logic;
signal \N__47772\ : std_logic;
signal \N__47769\ : std_logic;
signal \N__47766\ : std_logic;
signal \N__47763\ : std_logic;
signal \N__47762\ : std_logic;
signal \N__47759\ : std_logic;
signal \N__47756\ : std_logic;
signal \N__47753\ : std_logic;
signal \N__47750\ : std_logic;
signal \N__47747\ : std_logic;
signal \N__47744\ : std_logic;
signal \N__47741\ : std_logic;
signal \N__47738\ : std_logic;
signal \N__47735\ : std_logic;
signal \N__47730\ : std_logic;
signal \N__47723\ : std_logic;
signal \N__47722\ : std_logic;
signal \N__47719\ : std_logic;
signal \N__47718\ : std_logic;
signal \N__47715\ : std_logic;
signal \N__47712\ : std_logic;
signal \N__47709\ : std_logic;
signal \N__47702\ : std_logic;
signal \N__47701\ : std_logic;
signal \N__47700\ : std_logic;
signal \N__47699\ : std_logic;
signal \N__47698\ : std_logic;
signal \N__47697\ : std_logic;
signal \N__47696\ : std_logic;
signal \N__47695\ : std_logic;
signal \N__47694\ : std_logic;
signal \N__47693\ : std_logic;
signal \N__47692\ : std_logic;
signal \N__47691\ : std_logic;
signal \N__47690\ : std_logic;
signal \N__47689\ : std_logic;
signal \N__47688\ : std_logic;
signal \N__47687\ : std_logic;
signal \N__47686\ : std_logic;
signal \N__47685\ : std_logic;
signal \N__47684\ : std_logic;
signal \N__47683\ : std_logic;
signal \N__47682\ : std_logic;
signal \N__47681\ : std_logic;
signal \N__47680\ : std_logic;
signal \N__47679\ : std_logic;
signal \N__47678\ : std_logic;
signal \N__47677\ : std_logic;
signal \N__47676\ : std_logic;
signal \N__47675\ : std_logic;
signal \N__47674\ : std_logic;
signal \N__47673\ : std_logic;
signal \N__47672\ : std_logic;
signal \N__47671\ : std_logic;
signal \N__47670\ : std_logic;
signal \N__47669\ : std_logic;
signal \N__47668\ : std_logic;
signal \N__47667\ : std_logic;
signal \N__47666\ : std_logic;
signal \N__47665\ : std_logic;
signal \N__47664\ : std_logic;
signal \N__47663\ : std_logic;
signal \N__47662\ : std_logic;
signal \N__47661\ : std_logic;
signal \N__47660\ : std_logic;
signal \N__47659\ : std_logic;
signal \N__47658\ : std_logic;
signal \N__47657\ : std_logic;
signal \N__47656\ : std_logic;
signal \N__47655\ : std_logic;
signal \N__47654\ : std_logic;
signal \N__47653\ : std_logic;
signal \N__47652\ : std_logic;
signal \N__47651\ : std_logic;
signal \N__47650\ : std_logic;
signal \N__47649\ : std_logic;
signal \N__47648\ : std_logic;
signal \N__47647\ : std_logic;
signal \N__47646\ : std_logic;
signal \N__47645\ : std_logic;
signal \N__47644\ : std_logic;
signal \N__47643\ : std_logic;
signal \N__47642\ : std_logic;
signal \N__47641\ : std_logic;
signal \N__47640\ : std_logic;
signal \N__47639\ : std_logic;
signal \N__47638\ : std_logic;
signal \N__47637\ : std_logic;
signal \N__47636\ : std_logic;
signal \N__47635\ : std_logic;
signal \N__47634\ : std_logic;
signal \N__47633\ : std_logic;
signal \N__47632\ : std_logic;
signal \N__47631\ : std_logic;
signal \N__47630\ : std_logic;
signal \N__47629\ : std_logic;
signal \N__47628\ : std_logic;
signal \N__47627\ : std_logic;
signal \N__47626\ : std_logic;
signal \N__47625\ : std_logic;
signal \N__47624\ : std_logic;
signal \N__47623\ : std_logic;
signal \N__47622\ : std_logic;
signal \N__47621\ : std_logic;
signal \N__47620\ : std_logic;
signal \N__47619\ : std_logic;
signal \N__47618\ : std_logic;
signal \N__47617\ : std_logic;
signal \N__47616\ : std_logic;
signal \N__47615\ : std_logic;
signal \N__47614\ : std_logic;
signal \N__47613\ : std_logic;
signal \N__47612\ : std_logic;
signal \N__47611\ : std_logic;
signal \N__47610\ : std_logic;
signal \N__47609\ : std_logic;
signal \N__47608\ : std_logic;
signal \N__47607\ : std_logic;
signal \N__47606\ : std_logic;
signal \N__47605\ : std_logic;
signal \N__47604\ : std_logic;
signal \N__47603\ : std_logic;
signal \N__47602\ : std_logic;
signal \N__47601\ : std_logic;
signal \N__47600\ : std_logic;
signal \N__47599\ : std_logic;
signal \N__47598\ : std_logic;
signal \N__47597\ : std_logic;
signal \N__47596\ : std_logic;
signal \N__47595\ : std_logic;
signal \N__47594\ : std_logic;
signal \N__47593\ : std_logic;
signal \N__47592\ : std_logic;
signal \N__47591\ : std_logic;
signal \N__47590\ : std_logic;
signal \N__47589\ : std_logic;
signal \N__47588\ : std_logic;
signal \N__47587\ : std_logic;
signal \N__47586\ : std_logic;
signal \N__47585\ : std_logic;
signal \N__47584\ : std_logic;
signal \N__47583\ : std_logic;
signal \N__47582\ : std_logic;
signal \N__47581\ : std_logic;
signal \N__47580\ : std_logic;
signal \N__47579\ : std_logic;
signal \N__47578\ : std_logic;
signal \N__47577\ : std_logic;
signal \N__47576\ : std_logic;
signal \N__47575\ : std_logic;
signal \N__47574\ : std_logic;
signal \N__47573\ : std_logic;
signal \N__47572\ : std_logic;
signal \N__47571\ : std_logic;
signal \N__47570\ : std_logic;
signal \N__47569\ : std_logic;
signal \N__47568\ : std_logic;
signal \N__47567\ : std_logic;
signal \N__47566\ : std_logic;
signal \N__47565\ : std_logic;
signal \N__47564\ : std_logic;
signal \N__47563\ : std_logic;
signal \N__47562\ : std_logic;
signal \N__47561\ : std_logic;
signal \N__47560\ : std_logic;
signal \N__47559\ : std_logic;
signal \N__47558\ : std_logic;
signal \N__47557\ : std_logic;
signal \N__47556\ : std_logic;
signal \N__47555\ : std_logic;
signal \N__47554\ : std_logic;
signal \N__47553\ : std_logic;
signal \N__47552\ : std_logic;
signal \N__47551\ : std_logic;
signal \N__47550\ : std_logic;
signal \N__47549\ : std_logic;
signal \N__47240\ : std_logic;
signal \N__47237\ : std_logic;
signal \N__47236\ : std_logic;
signal \N__47233\ : std_logic;
signal \N__47230\ : std_logic;
signal \N__47229\ : std_logic;
signal \N__47224\ : std_logic;
signal \N__47221\ : std_logic;
signal \N__47220\ : std_logic;
signal \N__47219\ : std_logic;
signal \N__47216\ : std_logic;
signal \N__47213\ : std_logic;
signal \N__47210\ : std_logic;
signal \N__47209\ : std_logic;
signal \N__47208\ : std_logic;
signal \N__47205\ : std_logic;
signal \N__47204\ : std_logic;
signal \N__47203\ : std_logic;
signal \N__47202\ : std_logic;
signal \N__47195\ : std_logic;
signal \N__47192\ : std_logic;
signal \N__47191\ : std_logic;
signal \N__47190\ : std_logic;
signal \N__47189\ : std_logic;
signal \N__47188\ : std_logic;
signal \N__47185\ : std_logic;
signal \N__47182\ : std_logic;
signal \N__47179\ : std_logic;
signal \N__47176\ : std_logic;
signal \N__47173\ : std_logic;
signal \N__47172\ : std_logic;
signal \N__47171\ : std_logic;
signal \N__47166\ : std_logic;
signal \N__47165\ : std_logic;
signal \N__47164\ : std_logic;
signal \N__47163\ : std_logic;
signal \N__47162\ : std_logic;
signal \N__47161\ : std_logic;
signal \N__47160\ : std_logic;
signal \N__47159\ : std_logic;
signal \N__47158\ : std_logic;
signal \N__47157\ : std_logic;
signal \N__47156\ : std_logic;
signal \N__47155\ : std_logic;
signal \N__47154\ : std_logic;
signal \N__47153\ : std_logic;
signal \N__47152\ : std_logic;
signal \N__47151\ : std_logic;
signal \N__47150\ : std_logic;
signal \N__47147\ : std_logic;
signal \N__47140\ : std_logic;
signal \N__47137\ : std_logic;
signal \N__47134\ : std_logic;
signal \N__47131\ : std_logic;
signal \N__47126\ : std_logic;
signal \N__47123\ : std_logic;
signal \N__47120\ : std_logic;
signal \N__47119\ : std_logic;
signal \N__47118\ : std_logic;
signal \N__47117\ : std_logic;
signal \N__47116\ : std_logic;
signal \N__47115\ : std_logic;
signal \N__47114\ : std_logic;
signal \N__47113\ : std_logic;
signal \N__47110\ : std_logic;
signal \N__47101\ : std_logic;
signal \N__47092\ : std_logic;
signal \N__47083\ : std_logic;
signal \N__47074\ : std_logic;
signal \N__47071\ : std_logic;
signal \N__47070\ : std_logic;
signal \N__47069\ : std_logic;
signal \N__47068\ : std_logic;
signal \N__47067\ : std_logic;
signal \N__47062\ : std_logic;
signal \N__47053\ : std_logic;
signal \N__47050\ : std_logic;
signal \N__47043\ : std_logic;
signal \N__47034\ : std_logic;
signal \N__47029\ : std_logic;
signal \N__47026\ : std_logic;
signal \N__47019\ : std_logic;
signal \N__47010\ : std_logic;
signal \N__47005\ : std_logic;
signal \N__46998\ : std_logic;
signal \N__46993\ : std_logic;
signal \N__46990\ : std_logic;
signal \N__46987\ : std_logic;
signal \N__46984\ : std_logic;
signal \N__46981\ : std_logic;
signal \N__46978\ : std_logic;
signal \N__46975\ : std_logic;
signal \N__46970\ : std_logic;
signal \N__46961\ : std_logic;
signal \N__46960\ : std_logic;
signal \N__46959\ : std_logic;
signal \N__46958\ : std_logic;
signal \N__46955\ : std_logic;
signal \N__46950\ : std_logic;
signal \N__46947\ : std_logic;
signal \N__46944\ : std_logic;
signal \N__46941\ : std_logic;
signal \N__46940\ : std_logic;
signal \N__46939\ : std_logic;
signal \N__46938\ : std_logic;
signal \N__46937\ : std_logic;
signal \N__46936\ : std_logic;
signal \N__46933\ : std_logic;
signal \N__46932\ : std_logic;
signal \N__46931\ : std_logic;
signal \N__46930\ : std_logic;
signal \N__46929\ : std_logic;
signal \N__46928\ : std_logic;
signal \N__46927\ : std_logic;
signal \N__46926\ : std_logic;
signal \N__46925\ : std_logic;
signal \N__46924\ : std_logic;
signal \N__46923\ : std_logic;
signal \N__46922\ : std_logic;
signal \N__46921\ : std_logic;
signal \N__46920\ : std_logic;
signal \N__46919\ : std_logic;
signal \N__46918\ : std_logic;
signal \N__46917\ : std_logic;
signal \N__46916\ : std_logic;
signal \N__46915\ : std_logic;
signal \N__46914\ : std_logic;
signal \N__46913\ : std_logic;
signal \N__46912\ : std_logic;
signal \N__46911\ : std_logic;
signal \N__46910\ : std_logic;
signal \N__46909\ : std_logic;
signal \N__46908\ : std_logic;
signal \N__46907\ : std_logic;
signal \N__46906\ : std_logic;
signal \N__46905\ : std_logic;
signal \N__46904\ : std_logic;
signal \N__46903\ : std_logic;
signal \N__46902\ : std_logic;
signal \N__46901\ : std_logic;
signal \N__46900\ : std_logic;
signal \N__46899\ : std_logic;
signal \N__46898\ : std_logic;
signal \N__46897\ : std_logic;
signal \N__46896\ : std_logic;
signal \N__46895\ : std_logic;
signal \N__46894\ : std_logic;
signal \N__46893\ : std_logic;
signal \N__46892\ : std_logic;
signal \N__46891\ : std_logic;
signal \N__46890\ : std_logic;
signal \N__46889\ : std_logic;
signal \N__46888\ : std_logic;
signal \N__46887\ : std_logic;
signal \N__46886\ : std_logic;
signal \N__46885\ : std_logic;
signal \N__46884\ : std_logic;
signal \N__46883\ : std_logic;
signal \N__46882\ : std_logic;
signal \N__46881\ : std_logic;
signal \N__46880\ : std_logic;
signal \N__46879\ : std_logic;
signal \N__46878\ : std_logic;
signal \N__46877\ : std_logic;
signal \N__46876\ : std_logic;
signal \N__46875\ : std_logic;
signal \N__46874\ : std_logic;
signal \N__46873\ : std_logic;
signal \N__46872\ : std_logic;
signal \N__46871\ : std_logic;
signal \N__46870\ : std_logic;
signal \N__46869\ : std_logic;
signal \N__46868\ : std_logic;
signal \N__46867\ : std_logic;
signal \N__46866\ : std_logic;
signal \N__46865\ : std_logic;
signal \N__46864\ : std_logic;
signal \N__46863\ : std_logic;
signal \N__46862\ : std_logic;
signal \N__46861\ : std_logic;
signal \N__46860\ : std_logic;
signal \N__46859\ : std_logic;
signal \N__46858\ : std_logic;
signal \N__46857\ : std_logic;
signal \N__46856\ : std_logic;
signal \N__46855\ : std_logic;
signal \N__46854\ : std_logic;
signal \N__46853\ : std_logic;
signal \N__46852\ : std_logic;
signal \N__46851\ : std_logic;
signal \N__46850\ : std_logic;
signal \N__46849\ : std_logic;
signal \N__46848\ : std_logic;
signal \N__46847\ : std_logic;
signal \N__46846\ : std_logic;
signal \N__46845\ : std_logic;
signal \N__46844\ : std_logic;
signal \N__46843\ : std_logic;
signal \N__46842\ : std_logic;
signal \N__46841\ : std_logic;
signal \N__46840\ : std_logic;
signal \N__46839\ : std_logic;
signal \N__46838\ : std_logic;
signal \N__46837\ : std_logic;
signal \N__46836\ : std_logic;
signal \N__46835\ : std_logic;
signal \N__46834\ : std_logic;
signal \N__46833\ : std_logic;
signal \N__46832\ : std_logic;
signal \N__46831\ : std_logic;
signal \N__46830\ : std_logic;
signal \N__46829\ : std_logic;
signal \N__46828\ : std_logic;
signal \N__46827\ : std_logic;
signal \N__46826\ : std_logic;
signal \N__46825\ : std_logic;
signal \N__46824\ : std_logic;
signal \N__46823\ : std_logic;
signal \N__46822\ : std_logic;
signal \N__46821\ : std_logic;
signal \N__46820\ : std_logic;
signal \N__46819\ : std_logic;
signal \N__46818\ : std_logic;
signal \N__46817\ : std_logic;
signal \N__46816\ : std_logic;
signal \N__46815\ : std_logic;
signal \N__46814\ : std_logic;
signal \N__46813\ : std_logic;
signal \N__46812\ : std_logic;
signal \N__46811\ : std_logic;
signal \N__46810\ : std_logic;
signal \N__46809\ : std_logic;
signal \N__46808\ : std_logic;
signal \N__46807\ : std_logic;
signal \N__46806\ : std_logic;
signal \N__46805\ : std_logic;
signal \N__46804\ : std_logic;
signal \N__46803\ : std_logic;
signal \N__46802\ : std_logic;
signal \N__46801\ : std_logic;
signal \N__46800\ : std_logic;
signal \N__46799\ : std_logic;
signal \N__46798\ : std_logic;
signal \N__46797\ : std_logic;
signal \N__46796\ : std_logic;
signal \N__46795\ : std_logic;
signal \N__46794\ : std_logic;
signal \N__46793\ : std_logic;
signal \N__46792\ : std_logic;
signal \N__46791\ : std_logic;
signal \N__46790\ : std_logic;
signal \N__46789\ : std_logic;
signal \N__46788\ : std_logic;
signal \N__46787\ : std_logic;
signal \N__46786\ : std_logic;
signal \N__46785\ : std_logic;
signal \N__46784\ : std_logic;
signal \N__46783\ : std_logic;
signal \N__46466\ : std_logic;
signal \N__46463\ : std_logic;
signal \N__46460\ : std_logic;
signal \N__46457\ : std_logic;
signal \N__46454\ : std_logic;
signal \N__46451\ : std_logic;
signal \N__46448\ : std_logic;
signal \N__46445\ : std_logic;
signal \N__46444\ : std_logic;
signal \N__46439\ : std_logic;
signal \N__46436\ : std_logic;
signal \N__46435\ : std_logic;
signal \N__46434\ : std_logic;
signal \N__46429\ : std_logic;
signal \N__46426\ : std_logic;
signal \N__46423\ : std_logic;
signal \N__46418\ : std_logic;
signal \N__46415\ : std_logic;
signal \N__46414\ : std_logic;
signal \N__46411\ : std_logic;
signal \N__46408\ : std_logic;
signal \N__46403\ : std_logic;
signal \N__46402\ : std_logic;
signal \N__46399\ : std_logic;
signal \N__46396\ : std_logic;
signal \N__46393\ : std_logic;
signal \N__46388\ : std_logic;
signal \N__46387\ : std_logic;
signal \N__46382\ : std_logic;
signal \N__46379\ : std_logic;
signal \N__46376\ : std_logic;
signal \N__46373\ : std_logic;
signal \N__46370\ : std_logic;
signal \N__46367\ : std_logic;
signal \N__46366\ : std_logic;
signal \N__46365\ : std_logic;
signal \N__46362\ : std_logic;
signal \N__46359\ : std_logic;
signal \N__46356\ : std_logic;
signal \N__46351\ : std_logic;
signal \N__46346\ : std_logic;
signal \N__46345\ : std_logic;
signal \N__46342\ : std_logic;
signal \N__46339\ : std_logic;
signal \N__46334\ : std_logic;
signal \N__46331\ : std_logic;
signal \N__46330\ : std_logic;
signal \N__46329\ : std_logic;
signal \N__46326\ : std_logic;
signal \N__46323\ : std_logic;
signal \N__46320\ : std_logic;
signal \N__46317\ : std_logic;
signal \N__46314\ : std_logic;
signal \N__46307\ : std_logic;
signal \N__46306\ : std_logic;
signal \N__46303\ : std_logic;
signal \N__46300\ : std_logic;
signal \N__46295\ : std_logic;
signal \N__46292\ : std_logic;
signal \N__46289\ : std_logic;
signal \N__46286\ : std_logic;
signal \N__46283\ : std_logic;
signal \N__46280\ : std_logic;
signal \N__46277\ : std_logic;
signal \N__46274\ : std_logic;
signal \N__46271\ : std_logic;
signal \N__46270\ : std_logic;
signal \N__46267\ : std_logic;
signal \N__46264\ : std_logic;
signal \N__46259\ : std_logic;
signal \N__46256\ : std_logic;
signal \N__46255\ : std_logic;
signal \N__46254\ : std_logic;
signal \N__46253\ : std_logic;
signal \N__46250\ : std_logic;
signal \N__46249\ : std_logic;
signal \N__46248\ : std_logic;
signal \N__46247\ : std_logic;
signal \N__46244\ : std_logic;
signal \N__46243\ : std_logic;
signal \N__46242\ : std_logic;
signal \N__46239\ : std_logic;
signal \N__46236\ : std_logic;
signal \N__46235\ : std_logic;
signal \N__46234\ : std_logic;
signal \N__46233\ : std_logic;
signal \N__46232\ : std_logic;
signal \N__46231\ : std_logic;
signal \N__46228\ : std_logic;
signal \N__46219\ : std_logic;
signal \N__46210\ : std_logic;
signal \N__46209\ : std_logic;
signal \N__46208\ : std_logic;
signal \N__46203\ : std_logic;
signal \N__46196\ : std_logic;
signal \N__46191\ : std_logic;
signal \N__46188\ : std_logic;
signal \N__46185\ : std_logic;
signal \N__46184\ : std_logic;
signal \N__46183\ : std_logic;
signal \N__46182\ : std_logic;
signal \N__46181\ : std_logic;
signal \N__46180\ : std_logic;
signal \N__46179\ : std_logic;
signal \N__46178\ : std_logic;
signal \N__46177\ : std_logic;
signal \N__46176\ : std_logic;
signal \N__46175\ : std_logic;
signal \N__46174\ : std_logic;
signal \N__46173\ : std_logic;
signal \N__46172\ : std_logic;
signal \N__46171\ : std_logic;
signal \N__46170\ : std_logic;
signal \N__46169\ : std_logic;
signal \N__46166\ : std_logic;
signal \N__46163\ : std_logic;
signal \N__46160\ : std_logic;
signal \N__46155\ : std_logic;
signal \N__46152\ : std_logic;
signal \N__46135\ : std_logic;
signal \N__46120\ : std_logic;
signal \N__46117\ : std_logic;
signal \N__46114\ : std_logic;
signal \N__46111\ : std_logic;
signal \N__46108\ : std_logic;
signal \N__46105\ : std_logic;
signal \N__46098\ : std_logic;
signal \N__46089\ : std_logic;
signal \N__46082\ : std_logic;
signal \N__46079\ : std_logic;
signal \N__46076\ : std_logic;
signal \N__46075\ : std_logic;
signal \N__46074\ : std_logic;
signal \N__46073\ : std_logic;
signal \N__46072\ : std_logic;
signal \N__46071\ : std_logic;
signal \N__46068\ : std_logic;
signal \N__46065\ : std_logic;
signal \N__46064\ : std_logic;
signal \N__46061\ : std_logic;
signal \N__46058\ : std_logic;
signal \N__46057\ : std_logic;
signal \N__46054\ : std_logic;
signal \N__46051\ : std_logic;
signal \N__46048\ : std_logic;
signal \N__46045\ : std_logic;
signal \N__46038\ : std_logic;
signal \N__46031\ : std_logic;
signal \N__46028\ : std_logic;
signal \N__46021\ : std_logic;
signal \N__46018\ : std_logic;
signal \N__46015\ : std_logic;
signal \N__46010\ : std_logic;
signal \N__46007\ : std_logic;
signal \N__46004\ : std_logic;
signal \N__46001\ : std_logic;
signal \N__45998\ : std_logic;
signal \N__45995\ : std_logic;
signal \N__45992\ : std_logic;
signal \N__45991\ : std_logic;
signal \N__45986\ : std_logic;
signal \N__45983\ : std_logic;
signal \N__45980\ : std_logic;
signal \N__45979\ : std_logic;
signal \N__45974\ : std_logic;
signal \N__45971\ : std_logic;
signal \N__45970\ : std_logic;
signal \N__45967\ : std_logic;
signal \N__45964\ : std_logic;
signal \N__45959\ : std_logic;
signal \N__45958\ : std_logic;
signal \N__45957\ : std_logic;
signal \N__45956\ : std_logic;
signal \N__45955\ : std_logic;
signal \N__45954\ : std_logic;
signal \N__45953\ : std_logic;
signal \N__45952\ : std_logic;
signal \N__45935\ : std_logic;
signal \N__45932\ : std_logic;
signal \N__45929\ : std_logic;
signal \N__45928\ : std_logic;
signal \N__45927\ : std_logic;
signal \N__45926\ : std_logic;
signal \N__45923\ : std_logic;
signal \N__45920\ : std_logic;
signal \N__45917\ : std_logic;
signal \N__45914\ : std_logic;
signal \N__45911\ : std_logic;
signal \N__45906\ : std_logic;
signal \N__45903\ : std_logic;
signal \N__45900\ : std_logic;
signal \N__45895\ : std_logic;
signal \N__45892\ : std_logic;
signal \N__45889\ : std_logic;
signal \N__45884\ : std_logic;
signal \N__45883\ : std_logic;
signal \N__45882\ : std_logic;
signal \N__45879\ : std_logic;
signal \N__45876\ : std_logic;
signal \N__45873\ : std_logic;
signal \N__45868\ : std_logic;
signal \N__45863\ : std_logic;
signal \N__45862\ : std_logic;
signal \N__45859\ : std_logic;
signal \N__45858\ : std_logic;
signal \N__45855\ : std_logic;
signal \N__45852\ : std_logic;
signal \N__45849\ : std_logic;
signal \N__45842\ : std_logic;
signal \N__45841\ : std_logic;
signal \N__45840\ : std_logic;
signal \N__45837\ : std_logic;
signal \N__45834\ : std_logic;
signal \N__45831\ : std_logic;
signal \N__45830\ : std_logic;
signal \N__45827\ : std_logic;
signal \N__45824\ : std_logic;
signal \N__45821\ : std_logic;
signal \N__45818\ : std_logic;
signal \N__45815\ : std_logic;
signal \N__45812\ : std_logic;
signal \N__45809\ : std_logic;
signal \N__45806\ : std_logic;
signal \N__45803\ : std_logic;
signal \N__45800\ : std_logic;
signal \N__45797\ : std_logic;
signal \N__45788\ : std_logic;
signal \N__45787\ : std_logic;
signal \N__45786\ : std_logic;
signal \N__45783\ : std_logic;
signal \N__45780\ : std_logic;
signal \N__45777\ : std_logic;
signal \N__45770\ : std_logic;
signal \N__45769\ : std_logic;
signal \N__45766\ : std_logic;
signal \N__45763\ : std_logic;
signal \N__45758\ : std_logic;
signal \N__45757\ : std_logic;
signal \N__45756\ : std_logic;
signal \N__45753\ : std_logic;
signal \N__45750\ : std_logic;
signal \N__45747\ : std_logic;
signal \N__45742\ : std_logic;
signal \N__45739\ : std_logic;
signal \N__45736\ : std_logic;
signal \N__45731\ : std_logic;
signal \N__45728\ : std_logic;
signal \N__45725\ : std_logic;
signal \N__45722\ : std_logic;
signal \N__45719\ : std_logic;
signal \N__45716\ : std_logic;
signal \N__45713\ : std_logic;
signal \N__45712\ : std_logic;
signal \N__45709\ : std_logic;
signal \N__45706\ : std_logic;
signal \N__45705\ : std_logic;
signal \N__45704\ : std_logic;
signal \N__45699\ : std_logic;
signal \N__45696\ : std_logic;
signal \N__45693\ : std_logic;
signal \N__45688\ : std_logic;
signal \N__45685\ : std_logic;
signal \N__45682\ : std_logic;
signal \N__45679\ : std_logic;
signal \N__45676\ : std_logic;
signal \N__45673\ : std_logic;
signal \N__45668\ : std_logic;
signal \N__45667\ : std_logic;
signal \N__45664\ : std_logic;
signal \N__45663\ : std_logic;
signal \N__45660\ : std_logic;
signal \N__45657\ : std_logic;
signal \N__45654\ : std_logic;
signal \N__45647\ : std_logic;
signal \N__45644\ : std_logic;
signal \N__45641\ : std_logic;
signal \N__45638\ : std_logic;
signal \N__45637\ : std_logic;
signal \N__45632\ : std_logic;
signal \N__45629\ : std_logic;
signal \N__45628\ : std_logic;
signal \N__45623\ : std_logic;
signal \N__45620\ : std_logic;
signal \N__45619\ : std_logic;
signal \N__45616\ : std_logic;
signal \N__45615\ : std_logic;
signal \N__45610\ : std_logic;
signal \N__45607\ : std_logic;
signal \N__45604\ : std_logic;
signal \N__45599\ : std_logic;
signal \N__45598\ : std_logic;
signal \N__45595\ : std_logic;
signal \N__45594\ : std_logic;
signal \N__45589\ : std_logic;
signal \N__45586\ : std_logic;
signal \N__45583\ : std_logic;
signal \N__45578\ : std_logic;
signal \N__45575\ : std_logic;
signal \N__45572\ : std_logic;
signal \N__45569\ : std_logic;
signal \N__45566\ : std_logic;
signal \N__45563\ : std_logic;
signal \N__45560\ : std_logic;
signal \N__45557\ : std_logic;
signal \N__45556\ : std_logic;
signal \N__45555\ : std_logic;
signal \N__45552\ : std_logic;
signal \N__45549\ : std_logic;
signal \N__45546\ : std_logic;
signal \N__45543\ : std_logic;
signal \N__45540\ : std_logic;
signal \N__45539\ : std_logic;
signal \N__45536\ : std_logic;
signal \N__45531\ : std_logic;
signal \N__45528\ : std_logic;
signal \N__45525\ : std_logic;
signal \N__45522\ : std_logic;
signal \N__45519\ : std_logic;
signal \N__45516\ : std_logic;
signal \N__45513\ : std_logic;
signal \N__45506\ : std_logic;
signal \N__45503\ : std_logic;
signal \N__45500\ : std_logic;
signal \N__45499\ : std_logic;
signal \N__45498\ : std_logic;
signal \N__45497\ : std_logic;
signal \N__45494\ : std_logic;
signal \N__45489\ : std_logic;
signal \N__45488\ : std_logic;
signal \N__45485\ : std_logic;
signal \N__45482\ : std_logic;
signal \N__45479\ : std_logic;
signal \N__45476\ : std_logic;
signal \N__45473\ : std_logic;
signal \N__45470\ : std_logic;
signal \N__45467\ : std_logic;
signal \N__45462\ : std_logic;
signal \N__45457\ : std_logic;
signal \N__45454\ : std_logic;
signal \N__45449\ : std_logic;
signal \N__45448\ : std_logic;
signal \N__45445\ : std_logic;
signal \N__45440\ : std_logic;
signal \N__45437\ : std_logic;
signal \N__45436\ : std_logic;
signal \N__45433\ : std_logic;
signal \N__45430\ : std_logic;
signal \N__45427\ : std_logic;
signal \N__45422\ : std_logic;
signal \N__45419\ : std_logic;
signal \N__45418\ : std_logic;
signal \N__45415\ : std_logic;
signal \N__45412\ : std_logic;
signal \N__45407\ : std_logic;
signal \N__45406\ : std_logic;
signal \N__45403\ : std_logic;
signal \N__45400\ : std_logic;
signal \N__45397\ : std_logic;
signal \N__45392\ : std_logic;
signal \N__45389\ : std_logic;
signal \N__45386\ : std_logic;
signal \N__45383\ : std_logic;
signal \N__45380\ : std_logic;
signal \N__45377\ : std_logic;
signal \N__45374\ : std_logic;
signal \N__45371\ : std_logic;
signal \N__45370\ : std_logic;
signal \N__45365\ : std_logic;
signal \N__45362\ : std_logic;
signal \N__45361\ : std_logic;
signal \N__45358\ : std_logic;
signal \N__45355\ : std_logic;
signal \N__45352\ : std_logic;
signal \N__45347\ : std_logic;
signal \N__45346\ : std_logic;
signal \N__45343\ : std_logic;
signal \N__45338\ : std_logic;
signal \N__45337\ : std_logic;
signal \N__45334\ : std_logic;
signal \N__45331\ : std_logic;
signal \N__45328\ : std_logic;
signal \N__45323\ : std_logic;
signal \N__45320\ : std_logic;
signal \N__45317\ : std_logic;
signal \N__45314\ : std_logic;
signal \N__45311\ : std_logic;
signal \N__45310\ : std_logic;
signal \N__45305\ : std_logic;
signal \N__45302\ : std_logic;
signal \N__45299\ : std_logic;
signal \N__45296\ : std_logic;
signal \N__45293\ : std_logic;
signal \N__45290\ : std_logic;
signal \N__45287\ : std_logic;
signal \N__45286\ : std_logic;
signal \N__45281\ : std_logic;
signal \N__45278\ : std_logic;
signal \N__45277\ : std_logic;
signal \N__45276\ : std_logic;
signal \N__45273\ : std_logic;
signal \N__45270\ : std_logic;
signal \N__45267\ : std_logic;
signal \N__45262\ : std_logic;
signal \N__45257\ : std_logic;
signal \N__45256\ : std_logic;
signal \N__45253\ : std_logic;
signal \N__45250\ : std_logic;
signal \N__45247\ : std_logic;
signal \N__45244\ : std_logic;
signal \N__45243\ : std_logic;
signal \N__45238\ : std_logic;
signal \N__45235\ : std_logic;
signal \N__45232\ : std_logic;
signal \N__45227\ : std_logic;
signal \N__45226\ : std_logic;
signal \N__45221\ : std_logic;
signal \N__45218\ : std_logic;
signal \N__45217\ : std_logic;
signal \N__45212\ : std_logic;
signal \N__45211\ : std_logic;
signal \N__45208\ : std_logic;
signal \N__45205\ : std_logic;
signal \N__45202\ : std_logic;
signal \N__45199\ : std_logic;
signal \N__45194\ : std_logic;
signal \N__45191\ : std_logic;
signal \N__45190\ : std_logic;
signal \N__45187\ : std_logic;
signal \N__45186\ : std_logic;
signal \N__45183\ : std_logic;
signal \N__45182\ : std_logic;
signal \N__45179\ : std_logic;
signal \N__45172\ : std_logic;
signal \N__45167\ : std_logic;
signal \N__45166\ : std_logic;
signal \N__45163\ : std_logic;
signal \N__45158\ : std_logic;
signal \N__45157\ : std_logic;
signal \N__45154\ : std_logic;
signal \N__45151\ : std_logic;
signal \N__45150\ : std_logic;
signal \N__45147\ : std_logic;
signal \N__45144\ : std_logic;
signal \N__45141\ : std_logic;
signal \N__45136\ : std_logic;
signal \N__45131\ : std_logic;
signal \N__45128\ : std_logic;
signal \N__45125\ : std_logic;
signal \N__45122\ : std_logic;
signal \N__45119\ : std_logic;
signal \N__45116\ : std_logic;
signal \N__45113\ : std_logic;
signal \N__45110\ : std_logic;
signal \N__45107\ : std_logic;
signal \N__45104\ : std_logic;
signal \N__45101\ : std_logic;
signal \N__45100\ : std_logic;
signal \N__45095\ : std_logic;
signal \N__45092\ : std_logic;
signal \N__45089\ : std_logic;
signal \N__45088\ : std_logic;
signal \N__45083\ : std_logic;
signal \N__45080\ : std_logic;
signal \N__45079\ : std_logic;
signal \N__45076\ : std_logic;
signal \N__45073\ : std_logic;
signal \N__45072\ : std_logic;
signal \N__45071\ : std_logic;
signal \N__45066\ : std_logic;
signal \N__45061\ : std_logic;
signal \N__45056\ : std_logic;
signal \N__45055\ : std_logic;
signal \N__45054\ : std_logic;
signal \N__45053\ : std_logic;
signal \N__45052\ : std_logic;
signal \N__45051\ : std_logic;
signal \N__45050\ : std_logic;
signal \N__45047\ : std_logic;
signal \N__45046\ : std_logic;
signal \N__45045\ : std_logic;
signal \N__45044\ : std_logic;
signal \N__45043\ : std_logic;
signal \N__45040\ : std_logic;
signal \N__45039\ : std_logic;
signal \N__45038\ : std_logic;
signal \N__45037\ : std_logic;
signal \N__45036\ : std_logic;
signal \N__45035\ : std_logic;
signal \N__45034\ : std_logic;
signal \N__45033\ : std_logic;
signal \N__45032\ : std_logic;
signal \N__45031\ : std_logic;
signal \N__45030\ : std_logic;
signal \N__45029\ : std_logic;
signal \N__45028\ : std_logic;
signal \N__45027\ : std_logic;
signal \N__45024\ : std_logic;
signal \N__45023\ : std_logic;
signal \N__45020\ : std_logic;
signal \N__45019\ : std_logic;
signal \N__45016\ : std_logic;
signal \N__45015\ : std_logic;
signal \N__45014\ : std_logic;
signal \N__45013\ : std_logic;
signal \N__45012\ : std_logic;
signal \N__45011\ : std_logic;
signal \N__45010\ : std_logic;
signal \N__45009\ : std_logic;
signal \N__45008\ : std_logic;
signal \N__45007\ : std_logic;
signal \N__45006\ : std_logic;
signal \N__45005\ : std_logic;
signal \N__45004\ : std_logic;
signal \N__45003\ : std_logic;
signal \N__45000\ : std_logic;
signal \N__44999\ : std_logic;
signal \N__44998\ : std_logic;
signal \N__44997\ : std_logic;
signal \N__44996\ : std_logic;
signal \N__44995\ : std_logic;
signal \N__44994\ : std_logic;
signal \N__44989\ : std_logic;
signal \N__44986\ : std_logic;
signal \N__44983\ : std_logic;
signal \N__44980\ : std_logic;
signal \N__44979\ : std_logic;
signal \N__44976\ : std_logic;
signal \N__44975\ : std_logic;
signal \N__44974\ : std_logic;
signal \N__44973\ : std_logic;
signal \N__44972\ : std_logic;
signal \N__44971\ : std_logic;
signal \N__44970\ : std_logic;
signal \N__44969\ : std_logic;
signal \N__44966\ : std_logic;
signal \N__44965\ : std_logic;
signal \N__44962\ : std_logic;
signal \N__44961\ : std_logic;
signal \N__44958\ : std_logic;
signal \N__44955\ : std_logic;
signal \N__44954\ : std_logic;
signal \N__44949\ : std_logic;
signal \N__44948\ : std_logic;
signal \N__44939\ : std_logic;
signal \N__44938\ : std_logic;
signal \N__44937\ : std_logic;
signal \N__44936\ : std_logic;
signal \N__44935\ : std_logic;
signal \N__44934\ : std_logic;
signal \N__44933\ : std_logic;
signal \N__44932\ : std_logic;
signal \N__44931\ : std_logic;
signal \N__44928\ : std_logic;
signal \N__44927\ : std_logic;
signal \N__44926\ : std_logic;
signal \N__44925\ : std_logic;
signal \N__44924\ : std_logic;
signal \N__44923\ : std_logic;
signal \N__44920\ : std_logic;
signal \N__44919\ : std_logic;
signal \N__44902\ : std_logic;
signal \N__44899\ : std_logic;
signal \N__44898\ : std_logic;
signal \N__44895\ : std_logic;
signal \N__44894\ : std_logic;
signal \N__44891\ : std_logic;
signal \N__44890\ : std_logic;
signal \N__44887\ : std_logic;
signal \N__44886\ : std_logic;
signal \N__44883\ : std_logic;
signal \N__44882\ : std_logic;
signal \N__44879\ : std_logic;
signal \N__44878\ : std_logic;
signal \N__44875\ : std_logic;
signal \N__44874\ : std_logic;
signal \N__44871\ : std_logic;
signal \N__44870\ : std_logic;
signal \N__44867\ : std_logic;
signal \N__44866\ : std_logic;
signal \N__44863\ : std_logic;
signal \N__44862\ : std_logic;
signal \N__44859\ : std_logic;
signal \N__44858\ : std_logic;
signal \N__44853\ : std_logic;
signal \N__44852\ : std_logic;
signal \N__44851\ : std_logic;
signal \N__44850\ : std_logic;
signal \N__44847\ : std_logic;
signal \N__44844\ : std_logic;
signal \N__44841\ : std_logic;
signal \N__44838\ : std_logic;
signal \N__44835\ : std_logic;
signal \N__44834\ : std_logic;
signal \N__44833\ : std_logic;
signal \N__44830\ : std_logic;
signal \N__44829\ : std_logic;
signal \N__44828\ : std_logic;
signal \N__44827\ : std_logic;
signal \N__44824\ : std_logic;
signal \N__44821\ : std_logic;
signal \N__44818\ : std_logic;
signal \N__44811\ : std_logic;
signal \N__44810\ : std_logic;
signal \N__44807\ : std_logic;
signal \N__44806\ : std_logic;
signal \N__44803\ : std_logic;
signal \N__44802\ : std_logic;
signal \N__44799\ : std_logic;
signal \N__44798\ : std_logic;
signal \N__44795\ : std_logic;
signal \N__44794\ : std_logic;
signal \N__44791\ : std_logic;
signal \N__44790\ : std_logic;
signal \N__44787\ : std_logic;
signal \N__44786\ : std_logic;
signal \N__44783\ : std_logic;
signal \N__44782\ : std_logic;
signal \N__44781\ : std_logic;
signal \N__44780\ : std_logic;
signal \N__44779\ : std_logic;
signal \N__44778\ : std_logic;
signal \N__44777\ : std_logic;
signal \N__44776\ : std_logic;
signal \N__44775\ : std_logic;
signal \N__44772\ : std_logic;
signal \N__44769\ : std_logic;
signal \N__44764\ : std_logic;
signal \N__44761\ : std_logic;
signal \N__44756\ : std_logic;
signal \N__44753\ : std_logic;
signal \N__44750\ : std_logic;
signal \N__44747\ : std_logic;
signal \N__44732\ : std_logic;
signal \N__44717\ : std_logic;
signal \N__44712\ : std_logic;
signal \N__44709\ : std_logic;
signal \N__44692\ : std_logic;
signal \N__44675\ : std_logic;
signal \N__44662\ : std_logic;
signal \N__44659\ : std_logic;
signal \N__44652\ : std_logic;
signal \N__44645\ : std_logic;
signal \N__44628\ : std_logic;
signal \N__44627\ : std_logic;
signal \N__44626\ : std_logic;
signal \N__44625\ : std_logic;
signal \N__44624\ : std_logic;
signal \N__44623\ : std_logic;
signal \N__44622\ : std_logic;
signal \N__44619\ : std_logic;
signal \N__44612\ : std_logic;
signal \N__44597\ : std_logic;
signal \N__44580\ : std_logic;
signal \N__44577\ : std_logic;
signal \N__44576\ : std_logic;
signal \N__44573\ : std_logic;
signal \N__44572\ : std_logic;
signal \N__44569\ : std_logic;
signal \N__44568\ : std_logic;
signal \N__44565\ : std_logic;
signal \N__44564\ : std_logic;
signal \N__44561\ : std_logic;
signal \N__44560\ : std_logic;
signal \N__44557\ : std_logic;
signal \N__44556\ : std_logic;
signal \N__44553\ : std_logic;
signal \N__44552\ : std_logic;
signal \N__44545\ : std_logic;
signal \N__44542\ : std_logic;
signal \N__44539\ : std_logic;
signal \N__44518\ : std_logic;
signal \N__44515\ : std_logic;
signal \N__44508\ : std_logic;
signal \N__44505\ : std_logic;
signal \N__44494\ : std_logic;
signal \N__44485\ : std_logic;
signal \N__44468\ : std_logic;
signal \N__44455\ : std_logic;
signal \N__44446\ : std_logic;
signal \N__44429\ : std_logic;
signal \N__44428\ : std_logic;
signal \N__44427\ : std_logic;
signal \N__44426\ : std_logic;
signal \N__44425\ : std_logic;
signal \N__44424\ : std_logic;
signal \N__44423\ : std_logic;
signal \N__44422\ : std_logic;
signal \N__44421\ : std_logic;
signal \N__44420\ : std_logic;
signal \N__44419\ : std_logic;
signal \N__44418\ : std_logic;
signal \N__44417\ : std_logic;
signal \N__44416\ : std_logic;
signal \N__44415\ : std_logic;
signal \N__44414\ : std_logic;
signal \N__44411\ : std_logic;
signal \N__44408\ : std_logic;
signal \N__44407\ : std_logic;
signal \N__44406\ : std_logic;
signal \N__44405\ : std_logic;
signal \N__44404\ : std_logic;
signal \N__44403\ : std_logic;
signal \N__44402\ : std_logic;
signal \N__44401\ : std_logic;
signal \N__44400\ : std_logic;
signal \N__44399\ : std_logic;
signal \N__44398\ : std_logic;
signal \N__44397\ : std_logic;
signal \N__44396\ : std_logic;
signal \N__44395\ : std_logic;
signal \N__44394\ : std_logic;
signal \N__44393\ : std_logic;
signal \N__44392\ : std_logic;
signal \N__44391\ : std_logic;
signal \N__44390\ : std_logic;
signal \N__44389\ : std_logic;
signal \N__44388\ : std_logic;
signal \N__44385\ : std_logic;
signal \N__44382\ : std_logic;
signal \N__44369\ : std_logic;
signal \N__44366\ : std_logic;
signal \N__44365\ : std_logic;
signal \N__44364\ : std_logic;
signal \N__44363\ : std_logic;
signal \N__44362\ : std_logic;
signal \N__44361\ : std_logic;
signal \N__44360\ : std_logic;
signal \N__44359\ : std_logic;
signal \N__44356\ : std_logic;
signal \N__44355\ : std_logic;
signal \N__44352\ : std_logic;
signal \N__44349\ : std_logic;
signal \N__44344\ : std_logic;
signal \N__44339\ : std_logic;
signal \N__44336\ : std_logic;
signal \N__44323\ : std_logic;
signal \N__44316\ : std_logic;
signal \N__44311\ : std_logic;
signal \N__44302\ : std_logic;
signal \N__44299\ : std_logic;
signal \N__44298\ : std_logic;
signal \N__44297\ : std_logic;
signal \N__44296\ : std_logic;
signal \N__44295\ : std_logic;
signal \N__44294\ : std_logic;
signal \N__44293\ : std_logic;
signal \N__44292\ : std_logic;
signal \N__44291\ : std_logic;
signal \N__44288\ : std_logic;
signal \N__44283\ : std_logic;
signal \N__44282\ : std_logic;
signal \N__44281\ : std_logic;
signal \N__44280\ : std_logic;
signal \N__44279\ : std_logic;
signal \N__44278\ : std_logic;
signal \N__44277\ : std_logic;
signal \N__44272\ : std_logic;
signal \N__44269\ : std_logic;
signal \N__44252\ : std_logic;
signal \N__44249\ : std_logic;
signal \N__44246\ : std_logic;
signal \N__44243\ : std_logic;
signal \N__44240\ : std_logic;
signal \N__44239\ : std_logic;
signal \N__44236\ : std_logic;
signal \N__44227\ : std_logic;
signal \N__44222\ : std_logic;
signal \N__44219\ : std_logic;
signal \N__44216\ : std_logic;
signal \N__44201\ : std_logic;
signal \N__44200\ : std_logic;
signal \N__44199\ : std_logic;
signal \N__44198\ : std_logic;
signal \N__44197\ : std_logic;
signal \N__44196\ : std_logic;
signal \N__44195\ : std_logic;
signal \N__44194\ : std_logic;
signal \N__44193\ : std_logic;
signal \N__44192\ : std_logic;
signal \N__44191\ : std_logic;
signal \N__44190\ : std_logic;
signal \N__44189\ : std_logic;
signal \N__44184\ : std_logic;
signal \N__44171\ : std_logic;
signal \N__44162\ : std_logic;
signal \N__44155\ : std_logic;
signal \N__44152\ : std_logic;
signal \N__44145\ : std_logic;
signal \N__44138\ : std_logic;
signal \N__44123\ : std_logic;
signal \N__44118\ : std_logic;
signal \N__44115\ : std_logic;
signal \N__44110\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44102\ : std_logic;
signal \N__44095\ : std_logic;
signal \N__44078\ : std_logic;
signal \N__44075\ : std_logic;
signal \N__44072\ : std_logic;
signal \N__44069\ : std_logic;
signal \N__44066\ : std_logic;
signal \N__44063\ : std_logic;
signal \N__44062\ : std_logic;
signal \N__44061\ : std_logic;
signal \N__44058\ : std_logic;
signal \N__44055\ : std_logic;
signal \N__44052\ : std_logic;
signal \N__44047\ : std_logic;
signal \N__44046\ : std_logic;
signal \N__44043\ : std_logic;
signal \N__44040\ : std_logic;
signal \N__44037\ : std_logic;
signal \N__44034\ : std_logic;
signal \N__44029\ : std_logic;
signal \N__44024\ : std_logic;
signal \N__44021\ : std_logic;
signal \N__44018\ : std_logic;
signal \N__44015\ : std_logic;
signal \N__44012\ : std_logic;
signal \N__44009\ : std_logic;
signal \N__44008\ : std_logic;
signal \N__44007\ : std_logic;
signal \N__44004\ : std_logic;
signal \N__44001\ : std_logic;
signal \N__43998\ : std_logic;
signal \N__43997\ : std_logic;
signal \N__43990\ : std_logic;
signal \N__43987\ : std_logic;
signal \N__43982\ : std_logic;
signal \N__43979\ : std_logic;
signal \N__43976\ : std_logic;
signal \N__43973\ : std_logic;
signal \N__43970\ : std_logic;
signal \N__43967\ : std_logic;
signal \N__43966\ : std_logic;
signal \N__43963\ : std_logic;
signal \N__43960\ : std_logic;
signal \N__43959\ : std_logic;
signal \N__43956\ : std_logic;
signal \N__43953\ : std_logic;
signal \N__43950\ : std_logic;
signal \N__43949\ : std_logic;
signal \N__43946\ : std_logic;
signal \N__43943\ : std_logic;
signal \N__43940\ : std_logic;
signal \N__43937\ : std_logic;
signal \N__43934\ : std_logic;
signal \N__43931\ : std_logic;
signal \N__43928\ : std_logic;
signal \N__43925\ : std_logic;
signal \N__43916\ : std_logic;
signal \N__43913\ : std_logic;
signal \N__43910\ : std_logic;
signal \N__43907\ : std_logic;
signal \N__43904\ : std_logic;
signal \N__43901\ : std_logic;
signal \N__43900\ : std_logic;
signal \N__43899\ : std_logic;
signal \N__43896\ : std_logic;
signal \N__43891\ : std_logic;
signal \N__43890\ : std_logic;
signal \N__43885\ : std_logic;
signal \N__43882\ : std_logic;
signal \N__43879\ : std_logic;
signal \N__43876\ : std_logic;
signal \N__43871\ : std_logic;
signal \N__43868\ : std_logic;
signal \N__43865\ : std_logic;
signal \N__43862\ : std_logic;
signal \N__43859\ : std_logic;
signal \N__43856\ : std_logic;
signal \N__43855\ : std_logic;
signal \N__43852\ : std_logic;
signal \N__43851\ : std_logic;
signal \N__43848\ : std_logic;
signal \N__43847\ : std_logic;
signal \N__43846\ : std_logic;
signal \N__43845\ : std_logic;
signal \N__43844\ : std_logic;
signal \N__43843\ : std_logic;
signal \N__43840\ : std_logic;
signal \N__43837\ : std_logic;
signal \N__43830\ : std_logic;
signal \N__43827\ : std_logic;
signal \N__43822\ : std_logic;
signal \N__43821\ : std_logic;
signal \N__43818\ : std_logic;
signal \N__43811\ : std_logic;
signal \N__43808\ : std_logic;
signal \N__43805\ : std_logic;
signal \N__43804\ : std_logic;
signal \N__43799\ : std_logic;
signal \N__43796\ : std_logic;
signal \N__43793\ : std_logic;
signal \N__43790\ : std_logic;
signal \N__43781\ : std_logic;
signal \N__43778\ : std_logic;
signal \N__43775\ : std_logic;
signal \N__43772\ : std_logic;
signal \N__43769\ : std_logic;
signal \N__43766\ : std_logic;
signal \N__43763\ : std_logic;
signal \N__43760\ : std_logic;
signal \N__43757\ : std_logic;
signal \N__43754\ : std_logic;
signal \N__43751\ : std_logic;
signal \N__43750\ : std_logic;
signal \N__43747\ : std_logic;
signal \N__43744\ : std_logic;
signal \N__43743\ : std_logic;
signal \N__43740\ : std_logic;
signal \N__43735\ : std_logic;
signal \N__43730\ : std_logic;
signal \N__43727\ : std_logic;
signal \N__43726\ : std_logic;
signal \N__43723\ : std_logic;
signal \N__43720\ : std_logic;
signal \N__43717\ : std_logic;
signal \N__43716\ : std_logic;
signal \N__43711\ : std_logic;
signal \N__43708\ : std_logic;
signal \N__43703\ : std_logic;
signal \N__43700\ : std_logic;
signal \N__43697\ : std_logic;
signal \N__43694\ : std_logic;
signal \N__43691\ : std_logic;
signal \N__43688\ : std_logic;
signal \N__43685\ : std_logic;
signal \N__43684\ : std_logic;
signal \N__43681\ : std_logic;
signal \N__43680\ : std_logic;
signal \N__43679\ : std_logic;
signal \N__43676\ : std_logic;
signal \N__43673\ : std_logic;
signal \N__43668\ : std_logic;
signal \N__43665\ : std_logic;
signal \N__43660\ : std_logic;
signal \N__43657\ : std_logic;
signal \N__43654\ : std_logic;
signal \N__43649\ : std_logic;
signal \N__43646\ : std_logic;
signal \N__43645\ : std_logic;
signal \N__43644\ : std_logic;
signal \N__43641\ : std_logic;
signal \N__43638\ : std_logic;
signal \N__43635\ : std_logic;
signal \N__43628\ : std_logic;
signal \N__43625\ : std_logic;
signal \N__43622\ : std_logic;
signal \N__43619\ : std_logic;
signal \N__43616\ : std_logic;
signal \N__43613\ : std_logic;
signal \N__43610\ : std_logic;
signal \N__43607\ : std_logic;
signal \N__43604\ : std_logic;
signal \N__43601\ : std_logic;
signal \N__43598\ : std_logic;
signal \N__43595\ : std_logic;
signal \N__43594\ : std_logic;
signal \N__43593\ : std_logic;
signal \N__43590\ : std_logic;
signal \N__43587\ : std_logic;
signal \N__43584\ : std_logic;
signal \N__43581\ : std_logic;
signal \N__43574\ : std_logic;
signal \N__43573\ : std_logic;
signal \N__43572\ : std_logic;
signal \N__43571\ : std_logic;
signal \N__43570\ : std_logic;
signal \N__43569\ : std_logic;
signal \N__43568\ : std_logic;
signal \N__43567\ : std_logic;
signal \N__43550\ : std_logic;
signal \N__43547\ : std_logic;
signal \N__43544\ : std_logic;
signal \N__43541\ : std_logic;
signal \N__43538\ : std_logic;
signal \N__43535\ : std_logic;
signal \N__43532\ : std_logic;
signal \N__43529\ : std_logic;
signal \N__43526\ : std_logic;
signal \N__43523\ : std_logic;
signal \N__43520\ : std_logic;
signal \N__43517\ : std_logic;
signal \N__43516\ : std_logic;
signal \N__43513\ : std_logic;
signal \N__43510\ : std_logic;
signal \N__43507\ : std_logic;
signal \N__43506\ : std_logic;
signal \N__43501\ : std_logic;
signal \N__43498\ : std_logic;
signal \N__43493\ : std_logic;
signal \N__43490\ : std_logic;
signal \N__43487\ : std_logic;
signal \N__43484\ : std_logic;
signal \N__43481\ : std_logic;
signal \N__43478\ : std_logic;
signal \N__43475\ : std_logic;
signal \N__43474\ : std_logic;
signal \N__43473\ : std_logic;
signal \N__43470\ : std_logic;
signal \N__43467\ : std_logic;
signal \N__43464\ : std_logic;
signal \N__43457\ : std_logic;
signal \N__43454\ : std_logic;
signal \N__43451\ : std_logic;
signal \N__43448\ : std_logic;
signal \N__43445\ : std_logic;
signal \N__43442\ : std_logic;
signal \N__43441\ : std_logic;
signal \N__43438\ : std_logic;
signal \N__43435\ : std_logic;
signal \N__43432\ : std_logic;
signal \N__43429\ : std_logic;
signal \N__43424\ : std_logic;
signal \N__43423\ : std_logic;
signal \N__43420\ : std_logic;
signal \N__43417\ : std_logic;
signal \N__43412\ : std_logic;
signal \N__43409\ : std_logic;
signal \N__43406\ : std_logic;
signal \N__43403\ : std_logic;
signal \N__43400\ : std_logic;
signal \N__43397\ : std_logic;
signal \N__43396\ : std_logic;
signal \N__43393\ : std_logic;
signal \N__43392\ : std_logic;
signal \N__43389\ : std_logic;
signal \N__43386\ : std_logic;
signal \N__43383\ : std_logic;
signal \N__43378\ : std_logic;
signal \N__43375\ : std_logic;
signal \N__43370\ : std_logic;
signal \N__43367\ : std_logic;
signal \N__43364\ : std_logic;
signal \N__43361\ : std_logic;
signal \N__43358\ : std_logic;
signal \N__43355\ : std_logic;
signal \N__43352\ : std_logic;
signal \N__43349\ : std_logic;
signal \N__43348\ : std_logic;
signal \N__43345\ : std_logic;
signal \N__43342\ : std_logic;
signal \N__43341\ : std_logic;
signal \N__43338\ : std_logic;
signal \N__43335\ : std_logic;
signal \N__43332\ : std_logic;
signal \N__43325\ : std_logic;
signal \N__43322\ : std_logic;
signal \N__43319\ : std_logic;
signal \N__43316\ : std_logic;
signal \N__43313\ : std_logic;
signal \N__43310\ : std_logic;
signal \N__43309\ : std_logic;
signal \N__43306\ : std_logic;
signal \N__43303\ : std_logic;
signal \N__43300\ : std_logic;
signal \N__43297\ : std_logic;
signal \N__43294\ : std_logic;
signal \N__43291\ : std_logic;
signal \N__43290\ : std_logic;
signal \N__43285\ : std_logic;
signal \N__43282\ : std_logic;
signal \N__43277\ : std_logic;
signal \N__43274\ : std_logic;
signal \N__43271\ : std_logic;
signal \N__43268\ : std_logic;
signal \N__43265\ : std_logic;
signal \N__43262\ : std_logic;
signal \N__43261\ : std_logic;
signal \N__43258\ : std_logic;
signal \N__43255\ : std_logic;
signal \N__43252\ : std_logic;
signal \N__43249\ : std_logic;
signal \N__43248\ : std_logic;
signal \N__43245\ : std_logic;
signal \N__43242\ : std_logic;
signal \N__43239\ : std_logic;
signal \N__43232\ : std_logic;
signal \N__43229\ : std_logic;
signal \N__43226\ : std_logic;
signal \N__43223\ : std_logic;
signal \N__43220\ : std_logic;
signal \N__43217\ : std_logic;
signal \N__43216\ : std_logic;
signal \N__43211\ : std_logic;
signal \N__43210\ : std_logic;
signal \N__43207\ : std_logic;
signal \N__43204\ : std_logic;
signal \N__43199\ : std_logic;
signal \N__43196\ : std_logic;
signal \N__43193\ : std_logic;
signal \N__43190\ : std_logic;
signal \N__43187\ : std_logic;
signal \N__43184\ : std_logic;
signal \N__43183\ : std_logic;
signal \N__43178\ : std_logic;
signal \N__43177\ : std_logic;
signal \N__43174\ : std_logic;
signal \N__43171\ : std_logic;
signal \N__43166\ : std_logic;
signal \N__43163\ : std_logic;
signal \N__43160\ : std_logic;
signal \N__43157\ : std_logic;
signal \N__43154\ : std_logic;
signal \N__43151\ : std_logic;
signal \N__43148\ : std_logic;
signal \N__43147\ : std_logic;
signal \N__43144\ : std_logic;
signal \N__43141\ : std_logic;
signal \N__43140\ : std_logic;
signal \N__43137\ : std_logic;
signal \N__43134\ : std_logic;
signal \N__43131\ : std_logic;
signal \N__43124\ : std_logic;
signal \N__43121\ : std_logic;
signal \N__43118\ : std_logic;
signal \N__43117\ : std_logic;
signal \N__43114\ : std_logic;
signal \N__43111\ : std_logic;
signal \N__43108\ : std_logic;
signal \N__43105\ : std_logic;
signal \N__43102\ : std_logic;
signal \N__43101\ : std_logic;
signal \N__43098\ : std_logic;
signal \N__43095\ : std_logic;
signal \N__43092\ : std_logic;
signal \N__43085\ : std_logic;
signal \N__43082\ : std_logic;
signal \N__43079\ : std_logic;
signal \N__43076\ : std_logic;
signal \N__43073\ : std_logic;
signal \N__43070\ : std_logic;
signal \N__43069\ : std_logic;
signal \N__43066\ : std_logic;
signal \N__43063\ : std_logic;
signal \N__43062\ : std_logic;
signal \N__43059\ : std_logic;
signal \N__43056\ : std_logic;
signal \N__43053\ : std_logic;
signal \N__43046\ : std_logic;
signal \N__43043\ : std_logic;
signal \N__43040\ : std_logic;
signal \N__43037\ : std_logic;
signal \N__43034\ : std_logic;
signal \N__43031\ : std_logic;
signal \N__43028\ : std_logic;
signal \N__43027\ : std_logic;
signal \N__43024\ : std_logic;
signal \N__43021\ : std_logic;
signal \N__43018\ : std_logic;
signal \N__43017\ : std_logic;
signal \N__43014\ : std_logic;
signal \N__43011\ : std_logic;
signal \N__43008\ : std_logic;
signal \N__43001\ : std_logic;
signal \N__42998\ : std_logic;
signal \N__42995\ : std_logic;
signal \N__42994\ : std_logic;
signal \N__42993\ : std_logic;
signal \N__42990\ : std_logic;
signal \N__42987\ : std_logic;
signal \N__42984\ : std_logic;
signal \N__42981\ : std_logic;
signal \N__42978\ : std_logic;
signal \N__42971\ : std_logic;
signal \N__42968\ : std_logic;
signal \N__42965\ : std_logic;
signal \N__42962\ : std_logic;
signal \N__42959\ : std_logic;
signal \N__42956\ : std_logic;
signal \N__42955\ : std_logic;
signal \N__42952\ : std_logic;
signal \N__42949\ : std_logic;
signal \N__42948\ : std_logic;
signal \N__42943\ : std_logic;
signal \N__42940\ : std_logic;
signal \N__42935\ : std_logic;
signal \N__42932\ : std_logic;
signal \N__42931\ : std_logic;
signal \N__42928\ : std_logic;
signal \N__42927\ : std_logic;
signal \N__42924\ : std_logic;
signal \N__42921\ : std_logic;
signal \N__42918\ : std_logic;
signal \N__42915\ : std_logic;
signal \N__42910\ : std_logic;
signal \N__42905\ : std_logic;
signal \N__42902\ : std_logic;
signal \N__42899\ : std_logic;
signal \N__42896\ : std_logic;
signal \N__42893\ : std_logic;
signal \N__42890\ : std_logic;
signal \N__42889\ : std_logic;
signal \N__42886\ : std_logic;
signal \N__42883\ : std_logic;
signal \N__42880\ : std_logic;
signal \N__42877\ : std_logic;
signal \N__42876\ : std_logic;
signal \N__42871\ : std_logic;
signal \N__42868\ : std_logic;
signal \N__42863\ : std_logic;
signal \N__42860\ : std_logic;
signal \N__42857\ : std_logic;
signal \N__42854\ : std_logic;
signal \N__42851\ : std_logic;
signal \N__42848\ : std_logic;
signal \N__42845\ : std_logic;
signal \N__42844\ : std_logic;
signal \N__42839\ : std_logic;
signal \N__42838\ : std_logic;
signal \N__42835\ : std_logic;
signal \N__42832\ : std_logic;
signal \N__42827\ : std_logic;
signal \N__42824\ : std_logic;
signal \N__42821\ : std_logic;
signal \N__42818\ : std_logic;
signal \N__42815\ : std_logic;
signal \N__42812\ : std_logic;
signal \N__42809\ : std_logic;
signal \N__42806\ : std_logic;
signal \N__42803\ : std_logic;
signal \N__42800\ : std_logic;
signal \N__42799\ : std_logic;
signal \N__42796\ : std_logic;
signal \N__42793\ : std_logic;
signal \N__42792\ : std_logic;
signal \N__42789\ : std_logic;
signal \N__42786\ : std_logic;
signal \N__42783\ : std_logic;
signal \N__42776\ : std_logic;
signal \N__42773\ : std_logic;
signal \N__42770\ : std_logic;
signal \N__42767\ : std_logic;
signal \N__42764\ : std_logic;
signal \N__42761\ : std_logic;
signal \N__42760\ : std_logic;
signal \N__42757\ : std_logic;
signal \N__42754\ : std_logic;
signal \N__42751\ : std_logic;
signal \N__42748\ : std_logic;
signal \N__42747\ : std_logic;
signal \N__42742\ : std_logic;
signal \N__42739\ : std_logic;
signal \N__42734\ : std_logic;
signal \N__42731\ : std_logic;
signal \N__42728\ : std_logic;
signal \N__42725\ : std_logic;
signal \N__42722\ : std_logic;
signal \N__42719\ : std_logic;
signal \N__42716\ : std_logic;
signal \N__42715\ : std_logic;
signal \N__42712\ : std_logic;
signal \N__42709\ : std_logic;
signal \N__42706\ : std_logic;
signal \N__42703\ : std_logic;
signal \N__42702\ : std_logic;
signal \N__42697\ : std_logic;
signal \N__42694\ : std_logic;
signal \N__42689\ : std_logic;
signal \N__42686\ : std_logic;
signal \N__42683\ : std_logic;
signal \N__42680\ : std_logic;
signal \N__42677\ : std_logic;
signal \N__42674\ : std_logic;
signal \N__42671\ : std_logic;
signal \N__42670\ : std_logic;
signal \N__42667\ : std_logic;
signal \N__42664\ : std_logic;
signal \N__42661\ : std_logic;
signal \N__42660\ : std_logic;
signal \N__42655\ : std_logic;
signal \N__42652\ : std_logic;
signal \N__42647\ : std_logic;
signal \N__42644\ : std_logic;
signal \N__42641\ : std_logic;
signal \N__42638\ : std_logic;
signal \N__42635\ : std_logic;
signal \N__42632\ : std_logic;
signal \N__42631\ : std_logic;
signal \N__42628\ : std_logic;
signal \N__42625\ : std_logic;
signal \N__42622\ : std_logic;
signal \N__42621\ : std_logic;
signal \N__42618\ : std_logic;
signal \N__42615\ : std_logic;
signal \N__42612\ : std_logic;
signal \N__42605\ : std_logic;
signal \N__42602\ : std_logic;
signal \N__42599\ : std_logic;
signal \N__42598\ : std_logic;
signal \N__42597\ : std_logic;
signal \N__42596\ : std_logic;
signal \N__42593\ : std_logic;
signal \N__42588\ : std_logic;
signal \N__42585\ : std_logic;
signal \N__42582\ : std_logic;
signal \N__42579\ : std_logic;
signal \N__42576\ : std_logic;
signal \N__42573\ : std_logic;
signal \N__42570\ : std_logic;
signal \N__42567\ : std_logic;
signal \N__42560\ : std_logic;
signal \N__42559\ : std_logic;
signal \N__42554\ : std_logic;
signal \N__42551\ : std_logic;
signal \N__42548\ : std_logic;
signal \N__42547\ : std_logic;
signal \N__42546\ : std_logic;
signal \N__42545\ : std_logic;
signal \N__42542\ : std_logic;
signal \N__42537\ : std_logic;
signal \N__42534\ : std_logic;
signal \N__42529\ : std_logic;
signal \N__42526\ : std_logic;
signal \N__42523\ : std_logic;
signal \N__42518\ : std_logic;
signal \N__42517\ : std_logic;
signal \N__42514\ : std_logic;
signal \N__42511\ : std_logic;
signal \N__42510\ : std_logic;
signal \N__42507\ : std_logic;
signal \N__42504\ : std_logic;
signal \N__42501\ : std_logic;
signal \N__42498\ : std_logic;
signal \N__42495\ : std_logic;
signal \N__42488\ : std_logic;
signal \N__42485\ : std_logic;
signal \N__42482\ : std_logic;
signal \N__42479\ : std_logic;
signal \N__42476\ : std_logic;
signal \N__42473\ : std_logic;
signal \N__42470\ : std_logic;
signal \N__42467\ : std_logic;
signal \N__42466\ : std_logic;
signal \N__42463\ : std_logic;
signal \N__42462\ : std_logic;
signal \N__42459\ : std_logic;
signal \N__42456\ : std_logic;
signal \N__42453\ : std_logic;
signal \N__42450\ : std_logic;
signal \N__42445\ : std_logic;
signal \N__42444\ : std_logic;
signal \N__42441\ : std_logic;
signal \N__42438\ : std_logic;
signal \N__42435\ : std_logic;
signal \N__42428\ : std_logic;
signal \N__42425\ : std_logic;
signal \N__42422\ : std_logic;
signal \N__42419\ : std_logic;
signal \N__42416\ : std_logic;
signal \N__42415\ : std_logic;
signal \N__42414\ : std_logic;
signal \N__42411\ : std_logic;
signal \N__42408\ : std_logic;
signal \N__42405\ : std_logic;
signal \N__42400\ : std_logic;
signal \N__42397\ : std_logic;
signal \N__42394\ : std_logic;
signal \N__42391\ : std_logic;
signal \N__42388\ : std_logic;
signal \N__42383\ : std_logic;
signal \N__42382\ : std_logic;
signal \N__42381\ : std_logic;
signal \N__42380\ : std_logic;
signal \N__42377\ : std_logic;
signal \N__42374\ : std_logic;
signal \N__42371\ : std_logic;
signal \N__42370\ : std_logic;
signal \N__42369\ : std_logic;
signal \N__42368\ : std_logic;
signal \N__42367\ : std_logic;
signal \N__42366\ : std_logic;
signal \N__42365\ : std_logic;
signal \N__42364\ : std_logic;
signal \N__42363\ : std_logic;
signal \N__42362\ : std_logic;
signal \N__42361\ : std_logic;
signal \N__42360\ : std_logic;
signal \N__42359\ : std_logic;
signal \N__42358\ : std_logic;
signal \N__42355\ : std_logic;
signal \N__42352\ : std_logic;
signal \N__42349\ : std_logic;
signal \N__42346\ : std_logic;
signal \N__42331\ : std_logic;
signal \N__42318\ : std_logic;
signal \N__42317\ : std_logic;
signal \N__42316\ : std_logic;
signal \N__42315\ : std_logic;
signal \N__42314\ : std_logic;
signal \N__42313\ : std_logic;
signal \N__42312\ : std_logic;
signal \N__42311\ : std_logic;
signal \N__42310\ : std_logic;
signal \N__42305\ : std_logic;
signal \N__42296\ : std_logic;
signal \N__42287\ : std_logic;
signal \N__42278\ : std_logic;
signal \N__42275\ : std_logic;
signal \N__42266\ : std_logic;
signal \N__42265\ : std_logic;
signal \N__42262\ : std_logic;
signal \N__42261\ : std_logic;
signal \N__42258\ : std_logic;
signal \N__42255\ : std_logic;
signal \N__42252\ : std_logic;
signal \N__42247\ : std_logic;
signal \N__42242\ : std_logic;
signal \N__42239\ : std_logic;
signal \N__42236\ : std_logic;
signal \N__42233\ : std_logic;
signal \N__42230\ : std_logic;
signal \N__42227\ : std_logic;
signal \N__42226\ : std_logic;
signal \N__42221\ : std_logic;
signal \N__42218\ : std_logic;
signal \N__42217\ : std_logic;
signal \N__42214\ : std_logic;
signal \N__42211\ : std_logic;
signal \N__42206\ : std_logic;
signal \N__42203\ : std_logic;
signal \N__42200\ : std_logic;
signal \N__42197\ : std_logic;
signal \N__42194\ : std_logic;
signal \N__42191\ : std_logic;
signal \N__42190\ : std_logic;
signal \N__42187\ : std_logic;
signal \N__42184\ : std_logic;
signal \N__42181\ : std_logic;
signal \N__42178\ : std_logic;
signal \N__42177\ : std_logic;
signal \N__42172\ : std_logic;
signal \N__42169\ : std_logic;
signal \N__42164\ : std_logic;
signal \N__42161\ : std_logic;
signal \N__42158\ : std_logic;
signal \N__42155\ : std_logic;
signal \N__42152\ : std_logic;
signal \N__42149\ : std_logic;
signal \N__42146\ : std_logic;
signal \N__42145\ : std_logic;
signal \N__42142\ : std_logic;
signal \N__42139\ : std_logic;
signal \N__42136\ : std_logic;
signal \N__42133\ : std_logic;
signal \N__42130\ : std_logic;
signal \N__42127\ : std_logic;
signal \N__42122\ : std_logic;
signal \N__42121\ : std_logic;
signal \N__42118\ : std_logic;
signal \N__42115\ : std_logic;
signal \N__42110\ : std_logic;
signal \N__42109\ : std_logic;
signal \N__42106\ : std_logic;
signal \N__42103\ : std_logic;
signal \N__42100\ : std_logic;
signal \N__42097\ : std_logic;
signal \N__42094\ : std_logic;
signal \N__42091\ : std_logic;
signal \N__42086\ : std_logic;
signal \N__42083\ : std_logic;
signal \N__42080\ : std_logic;
signal \N__42077\ : std_logic;
signal \N__42074\ : std_logic;
signal \N__42071\ : std_logic;
signal \N__42068\ : std_logic;
signal \N__42065\ : std_logic;
signal \N__42062\ : std_logic;
signal \N__42059\ : std_logic;
signal \N__42058\ : std_logic;
signal \N__42055\ : std_logic;
signal \N__42052\ : std_logic;
signal \N__42047\ : std_logic;
signal \N__42044\ : std_logic;
signal \N__42041\ : std_logic;
signal \N__42040\ : std_logic;
signal \N__42037\ : std_logic;
signal \N__42034\ : std_logic;
signal \N__42031\ : std_logic;
signal \N__42028\ : std_logic;
signal \N__42025\ : std_logic;
signal \N__42022\ : std_logic;
signal \N__42021\ : std_logic;
signal \N__42020\ : std_logic;
signal \N__42017\ : std_logic;
signal \N__42014\ : std_logic;
signal \N__42009\ : std_logic;
signal \N__42002\ : std_logic;
signal \N__41999\ : std_logic;
signal \N__41996\ : std_logic;
signal \N__41993\ : std_logic;
signal \N__41990\ : std_logic;
signal \N__41987\ : std_logic;
signal \N__41984\ : std_logic;
signal \N__41983\ : std_logic;
signal \N__41982\ : std_logic;
signal \N__41979\ : std_logic;
signal \N__41974\ : std_logic;
signal \N__41969\ : std_logic;
signal \N__41968\ : std_logic;
signal \N__41965\ : std_logic;
signal \N__41964\ : std_logic;
signal \N__41961\ : std_logic;
signal \N__41956\ : std_logic;
signal \N__41951\ : std_logic;
signal \N__41948\ : std_logic;
signal \N__41945\ : std_logic;
signal \N__41942\ : std_logic;
signal \N__41939\ : std_logic;
signal \N__41936\ : std_logic;
signal \N__41935\ : std_logic;
signal \N__41932\ : std_logic;
signal \N__41929\ : std_logic;
signal \N__41926\ : std_logic;
signal \N__41925\ : std_logic;
signal \N__41922\ : std_logic;
signal \N__41919\ : std_logic;
signal \N__41916\ : std_logic;
signal \N__41911\ : std_logic;
signal \N__41906\ : std_logic;
signal \N__41905\ : std_logic;
signal \N__41904\ : std_logic;
signal \N__41901\ : std_logic;
signal \N__41900\ : std_logic;
signal \N__41897\ : std_logic;
signal \N__41894\ : std_logic;
signal \N__41891\ : std_logic;
signal \N__41888\ : std_logic;
signal \N__41885\ : std_logic;
signal \N__41880\ : std_logic;
signal \N__41877\ : std_logic;
signal \N__41872\ : std_logic;
signal \N__41867\ : std_logic;
signal \N__41864\ : std_logic;
signal \N__41863\ : std_logic;
signal \N__41858\ : std_logic;
signal \N__41855\ : std_logic;
signal \N__41852\ : std_logic;
signal \N__41849\ : std_logic;
signal \N__41846\ : std_logic;
signal \N__41845\ : std_logic;
signal \N__41842\ : std_logic;
signal \N__41839\ : std_logic;
signal \N__41834\ : std_logic;
signal \N__41833\ : std_logic;
signal \N__41830\ : std_logic;
signal \N__41829\ : std_logic;
signal \N__41826\ : std_logic;
signal \N__41823\ : std_logic;
signal \N__41820\ : std_logic;
signal \N__41813\ : std_logic;
signal \N__41810\ : std_logic;
signal \N__41809\ : std_logic;
signal \N__41808\ : std_logic;
signal \N__41805\ : std_logic;
signal \N__41802\ : std_logic;
signal \N__41799\ : std_logic;
signal \N__41792\ : std_logic;
signal \N__41791\ : std_logic;
signal \N__41788\ : std_logic;
signal \N__41785\ : std_logic;
signal \N__41780\ : std_logic;
signal \N__41777\ : std_logic;
signal \N__41774\ : std_logic;
signal \N__41771\ : std_logic;
signal \N__41768\ : std_logic;
signal \N__41765\ : std_logic;
signal \N__41764\ : std_logic;
signal \N__41761\ : std_logic;
signal \N__41758\ : std_logic;
signal \N__41755\ : std_logic;
signal \N__41754\ : std_logic;
signal \N__41749\ : std_logic;
signal \N__41746\ : std_logic;
signal \N__41741\ : std_logic;
signal \N__41740\ : std_logic;
signal \N__41739\ : std_logic;
signal \N__41738\ : std_logic;
signal \N__41735\ : std_logic;
signal \N__41732\ : std_logic;
signal \N__41729\ : std_logic;
signal \N__41726\ : std_logic;
signal \N__41723\ : std_logic;
signal \N__41720\ : std_logic;
signal \N__41717\ : std_logic;
signal \N__41712\ : std_logic;
signal \N__41707\ : std_logic;
signal \N__41704\ : std_logic;
signal \N__41701\ : std_logic;
signal \N__41698\ : std_logic;
signal \N__41693\ : std_logic;
signal \N__41692\ : std_logic;
signal \N__41691\ : std_logic;
signal \N__41688\ : std_logic;
signal \N__41685\ : std_logic;
signal \N__41682\ : std_logic;
signal \N__41675\ : std_logic;
signal \N__41674\ : std_logic;
signal \N__41673\ : std_logic;
signal \N__41672\ : std_logic;
signal \N__41669\ : std_logic;
signal \N__41666\ : std_logic;
signal \N__41663\ : std_logic;
signal \N__41660\ : std_logic;
signal \N__41657\ : std_logic;
signal \N__41652\ : std_logic;
signal \N__41649\ : std_logic;
signal \N__41644\ : std_logic;
signal \N__41641\ : std_logic;
signal \N__41638\ : std_logic;
signal \N__41635\ : std_logic;
signal \N__41630\ : std_logic;
signal \N__41629\ : std_logic;
signal \N__41626\ : std_logic;
signal \N__41623\ : std_logic;
signal \N__41618\ : std_logic;
signal \N__41615\ : std_logic;
signal \N__41612\ : std_logic;
signal \N__41609\ : std_logic;
signal \N__41606\ : std_logic;
signal \N__41603\ : std_logic;
signal \N__41602\ : std_logic;
signal \N__41597\ : std_logic;
signal \N__41594\ : std_logic;
signal \N__41593\ : std_logic;
signal \N__41588\ : std_logic;
signal \N__41587\ : std_logic;
signal \N__41584\ : std_logic;
signal \N__41581\ : std_logic;
signal \N__41578\ : std_logic;
signal \N__41573\ : std_logic;
signal \N__41572\ : std_logic;
signal \N__41569\ : std_logic;
signal \N__41568\ : std_logic;
signal \N__41563\ : std_logic;
signal \N__41560\ : std_logic;
signal \N__41557\ : std_logic;
signal \N__41552\ : std_logic;
signal \N__41551\ : std_logic;
signal \N__41548\ : std_logic;
signal \N__41543\ : std_logic;
signal \N__41540\ : std_logic;
signal \N__41537\ : std_logic;
signal \N__41534\ : std_logic;
signal \N__41531\ : std_logic;
signal \N__41528\ : std_logic;
signal \N__41525\ : std_logic;
signal \N__41524\ : std_logic;
signal \N__41521\ : std_logic;
signal \N__41520\ : std_logic;
signal \N__41517\ : std_logic;
signal \N__41514\ : std_logic;
signal \N__41511\ : std_logic;
signal \N__41504\ : std_logic;
signal \N__41503\ : std_logic;
signal \N__41502\ : std_logic;
signal \N__41501\ : std_logic;
signal \N__41498\ : std_logic;
signal \N__41495\ : std_logic;
signal \N__41492\ : std_logic;
signal \N__41489\ : std_logic;
signal \N__41484\ : std_logic;
signal \N__41479\ : std_logic;
signal \N__41474\ : std_logic;
signal \N__41471\ : std_logic;
signal \N__41468\ : std_logic;
signal \N__41465\ : std_logic;
signal \N__41462\ : std_logic;
signal \N__41459\ : std_logic;
signal \N__41456\ : std_logic;
signal \N__41455\ : std_logic;
signal \N__41454\ : std_logic;
signal \N__41451\ : std_logic;
signal \N__41448\ : std_logic;
signal \N__41447\ : std_logic;
signal \N__41444\ : std_logic;
signal \N__41439\ : std_logic;
signal \N__41436\ : std_logic;
signal \N__41433\ : std_logic;
signal \N__41428\ : std_logic;
signal \N__41423\ : std_logic;
signal \N__41420\ : std_logic;
signal \N__41417\ : std_logic;
signal \N__41416\ : std_logic;
signal \N__41415\ : std_logic;
signal \N__41412\ : std_logic;
signal \N__41409\ : std_logic;
signal \N__41406\ : std_logic;
signal \N__41401\ : std_logic;
signal \N__41396\ : std_logic;
signal \N__41395\ : std_logic;
signal \N__41394\ : std_logic;
signal \N__41389\ : std_logic;
signal \N__41386\ : std_logic;
signal \N__41383\ : std_logic;
signal \N__41378\ : std_logic;
signal \N__41375\ : std_logic;
signal \N__41372\ : std_logic;
signal \N__41371\ : std_logic;
signal \N__41368\ : std_logic;
signal \N__41365\ : std_logic;
signal \N__41362\ : std_logic;
signal \N__41357\ : std_logic;
signal \N__41354\ : std_logic;
signal \N__41353\ : std_logic;
signal \N__41352\ : std_logic;
signal \N__41351\ : std_logic;
signal \N__41350\ : std_logic;
signal \N__41349\ : std_logic;
signal \N__41348\ : std_logic;
signal \N__41347\ : std_logic;
signal \N__41346\ : std_logic;
signal \N__41345\ : std_logic;
signal \N__41344\ : std_logic;
signal \N__41343\ : std_logic;
signal \N__41342\ : std_logic;
signal \N__41341\ : std_logic;
signal \N__41340\ : std_logic;
signal \N__41339\ : std_logic;
signal \N__41338\ : std_logic;
signal \N__41337\ : std_logic;
signal \N__41336\ : std_logic;
signal \N__41335\ : std_logic;
signal \N__41334\ : std_logic;
signal \N__41333\ : std_logic;
signal \N__41332\ : std_logic;
signal \N__41331\ : std_logic;
signal \N__41330\ : std_logic;
signal \N__41329\ : std_logic;
signal \N__41328\ : std_logic;
signal \N__41327\ : std_logic;
signal \N__41326\ : std_logic;
signal \N__41325\ : std_logic;
signal \N__41316\ : std_logic;
signal \N__41307\ : std_logic;
signal \N__41302\ : std_logic;
signal \N__41293\ : std_logic;
signal \N__41284\ : std_logic;
signal \N__41275\ : std_logic;
signal \N__41266\ : std_logic;
signal \N__41257\ : std_logic;
signal \N__41254\ : std_logic;
signal \N__41247\ : std_logic;
signal \N__41240\ : std_logic;
signal \N__41237\ : std_logic;
signal \N__41234\ : std_logic;
signal \N__41229\ : std_logic;
signal \N__41224\ : std_logic;
signal \N__41219\ : std_logic;
signal \N__41216\ : std_logic;
signal \N__41213\ : std_logic;
signal \N__41212\ : std_logic;
signal \N__41209\ : std_logic;
signal \N__41206\ : std_logic;
signal \N__41203\ : std_logic;
signal \N__41198\ : std_logic;
signal \N__41197\ : std_logic;
signal \N__41194\ : std_logic;
signal \N__41193\ : std_logic;
signal \N__41190\ : std_logic;
signal \N__41187\ : std_logic;
signal \N__41186\ : std_logic;
signal \N__41183\ : std_logic;
signal \N__41180\ : std_logic;
signal \N__41177\ : std_logic;
signal \N__41174\ : std_logic;
signal \N__41171\ : std_logic;
signal \N__41168\ : std_logic;
signal \N__41163\ : std_logic;
signal \N__41160\ : std_logic;
signal \N__41155\ : std_logic;
signal \N__41150\ : std_logic;
signal \N__41149\ : std_logic;
signal \N__41148\ : std_logic;
signal \N__41147\ : std_logic;
signal \N__41144\ : std_logic;
signal \N__41141\ : std_logic;
signal \N__41136\ : std_logic;
signal \N__41133\ : std_logic;
signal \N__41128\ : std_logic;
signal \N__41125\ : std_logic;
signal \N__41122\ : std_logic;
signal \N__41119\ : std_logic;
signal \N__41114\ : std_logic;
signal \N__41113\ : std_logic;
signal \N__41112\ : std_logic;
signal \N__41111\ : std_logic;
signal \N__41106\ : std_logic;
signal \N__41103\ : std_logic;
signal \N__41100\ : std_logic;
signal \N__41097\ : std_logic;
signal \N__41094\ : std_logic;
signal \N__41091\ : std_logic;
signal \N__41088\ : std_logic;
signal \N__41085\ : std_logic;
signal \N__41082\ : std_logic;
signal \N__41079\ : std_logic;
signal \N__41076\ : std_logic;
signal \N__41069\ : std_logic;
signal \N__41066\ : std_logic;
signal \N__41063\ : std_logic;
signal \N__41062\ : std_logic;
signal \N__41059\ : std_logic;
signal \N__41056\ : std_logic;
signal \N__41053\ : std_logic;
signal \N__41050\ : std_logic;
signal \N__41047\ : std_logic;
signal \N__41046\ : std_logic;
signal \N__41045\ : std_logic;
signal \N__41042\ : std_logic;
signal \N__41039\ : std_logic;
signal \N__41034\ : std_logic;
signal \N__41031\ : std_logic;
signal \N__41024\ : std_logic;
signal \N__41021\ : std_logic;
signal \N__41018\ : std_logic;
signal \N__41017\ : std_logic;
signal \N__41016\ : std_logic;
signal \N__41011\ : std_logic;
signal \N__41008\ : std_logic;
signal \N__41005\ : std_logic;
signal \N__41000\ : std_logic;
signal \N__40997\ : std_logic;
signal \N__40994\ : std_logic;
signal \N__40993\ : std_logic;
signal \N__40992\ : std_logic;
signal \N__40989\ : std_logic;
signal \N__40986\ : std_logic;
signal \N__40983\ : std_logic;
signal \N__40978\ : std_logic;
signal \N__40973\ : std_logic;
signal \N__40970\ : std_logic;
signal \N__40969\ : std_logic;
signal \N__40966\ : std_logic;
signal \N__40963\ : std_logic;
signal \N__40962\ : std_logic;
signal \N__40957\ : std_logic;
signal \N__40954\ : std_logic;
signal \N__40951\ : std_logic;
signal \N__40946\ : std_logic;
signal \N__40943\ : std_logic;
signal \N__40942\ : std_logic;
signal \N__40941\ : std_logic;
signal \N__40936\ : std_logic;
signal \N__40933\ : std_logic;
signal \N__40930\ : std_logic;
signal \N__40925\ : std_logic;
signal \N__40922\ : std_logic;
signal \N__40921\ : std_logic;
signal \N__40920\ : std_logic;
signal \N__40915\ : std_logic;
signal \N__40912\ : std_logic;
signal \N__40909\ : std_logic;
signal \N__40904\ : std_logic;
signal \N__40901\ : std_logic;
signal \N__40900\ : std_logic;
signal \N__40897\ : std_logic;
signal \N__40894\ : std_logic;
signal \N__40893\ : std_logic;
signal \N__40888\ : std_logic;
signal \N__40885\ : std_logic;
signal \N__40882\ : std_logic;
signal \N__40877\ : std_logic;
signal \N__40874\ : std_logic;
signal \N__40873\ : std_logic;
signal \N__40870\ : std_logic;
signal \N__40867\ : std_logic;
signal \N__40864\ : std_logic;
signal \N__40863\ : std_logic;
signal \N__40860\ : std_logic;
signal \N__40857\ : std_logic;
signal \N__40854\ : std_logic;
signal \N__40851\ : std_logic;
signal \N__40848\ : std_logic;
signal \N__40841\ : std_logic;
signal \N__40838\ : std_logic;
signal \N__40837\ : std_logic;
signal \N__40834\ : std_logic;
signal \N__40831\ : std_logic;
signal \N__40830\ : std_logic;
signal \N__40827\ : std_logic;
signal \N__40824\ : std_logic;
signal \N__40821\ : std_logic;
signal \N__40818\ : std_logic;
signal \N__40815\ : std_logic;
signal \N__40808\ : std_logic;
signal \N__40805\ : std_logic;
signal \N__40804\ : std_logic;
signal \N__40803\ : std_logic;
signal \N__40798\ : std_logic;
signal \N__40795\ : std_logic;
signal \N__40792\ : std_logic;
signal \N__40787\ : std_logic;
signal \N__40784\ : std_logic;
signal \N__40783\ : std_logic;
signal \N__40782\ : std_logic;
signal \N__40777\ : std_logic;
signal \N__40774\ : std_logic;
signal \N__40771\ : std_logic;
signal \N__40766\ : std_logic;
signal \N__40763\ : std_logic;
signal \N__40762\ : std_logic;
signal \N__40761\ : std_logic;
signal \N__40756\ : std_logic;
signal \N__40753\ : std_logic;
signal \N__40750\ : std_logic;
signal \N__40745\ : std_logic;
signal \N__40742\ : std_logic;
signal \N__40741\ : std_logic;
signal \N__40738\ : std_logic;
signal \N__40737\ : std_logic;
signal \N__40734\ : std_logic;
signal \N__40731\ : std_logic;
signal \N__40728\ : std_logic;
signal \N__40723\ : std_logic;
signal \N__40718\ : std_logic;
signal \N__40715\ : std_logic;
signal \N__40714\ : std_logic;
signal \N__40711\ : std_logic;
signal \N__40710\ : std_logic;
signal \N__40707\ : std_logic;
signal \N__40704\ : std_logic;
signal \N__40701\ : std_logic;
signal \N__40696\ : std_logic;
signal \N__40691\ : std_logic;
signal \N__40688\ : std_logic;
signal \N__40687\ : std_logic;
signal \N__40684\ : std_logic;
signal \N__40681\ : std_logic;
signal \N__40680\ : std_logic;
signal \N__40675\ : std_logic;
signal \N__40672\ : std_logic;
signal \N__40669\ : std_logic;
signal \N__40664\ : std_logic;
signal \N__40661\ : std_logic;
signal \N__40660\ : std_logic;
signal \N__40657\ : std_logic;
signal \N__40654\ : std_logic;
signal \N__40653\ : std_logic;
signal \N__40648\ : std_logic;
signal \N__40645\ : std_logic;
signal \N__40642\ : std_logic;
signal \N__40637\ : std_logic;
signal \N__40634\ : std_logic;
signal \N__40633\ : std_logic;
signal \N__40630\ : std_logic;
signal \N__40627\ : std_logic;
signal \N__40626\ : std_logic;
signal \N__40623\ : std_logic;
signal \N__40620\ : std_logic;
signal \N__40617\ : std_logic;
signal \N__40614\ : std_logic;
signal \N__40611\ : std_logic;
signal \N__40604\ : std_logic;
signal \N__40601\ : std_logic;
signal \N__40600\ : std_logic;
signal \N__40597\ : std_logic;
signal \N__40594\ : std_logic;
signal \N__40591\ : std_logic;
signal \N__40588\ : std_logic;
signal \N__40587\ : std_logic;
signal \N__40582\ : std_logic;
signal \N__40579\ : std_logic;
signal \N__40576\ : std_logic;
signal \N__40571\ : std_logic;
signal \N__40568\ : std_logic;
signal \N__40567\ : std_logic;
signal \N__40566\ : std_logic;
signal \N__40561\ : std_logic;
signal \N__40558\ : std_logic;
signal \N__40555\ : std_logic;
signal \N__40550\ : std_logic;
signal \N__40547\ : std_logic;
signal \N__40546\ : std_logic;
signal \N__40543\ : std_logic;
signal \N__40540\ : std_logic;
signal \N__40537\ : std_logic;
signal \N__40536\ : std_logic;
signal \N__40531\ : std_logic;
signal \N__40528\ : std_logic;
signal \N__40525\ : std_logic;
signal \N__40520\ : std_logic;
signal \N__40517\ : std_logic;
signal \N__40516\ : std_logic;
signal \N__40513\ : std_logic;
signal \N__40510\ : std_logic;
signal \N__40509\ : std_logic;
signal \N__40504\ : std_logic;
signal \N__40501\ : std_logic;
signal \N__40498\ : std_logic;
signal \N__40493\ : std_logic;
signal \N__40490\ : std_logic;
signal \N__40489\ : std_logic;
signal \N__40486\ : std_logic;
signal \N__40483\ : std_logic;
signal \N__40482\ : std_logic;
signal \N__40477\ : std_logic;
signal \N__40474\ : std_logic;
signal \N__40471\ : std_logic;
signal \N__40466\ : std_logic;
signal \N__40463\ : std_logic;
signal \N__40462\ : std_logic;
signal \N__40461\ : std_logic;
signal \N__40456\ : std_logic;
signal \N__40453\ : std_logic;
signal \N__40450\ : std_logic;
signal \N__40445\ : std_logic;
signal \N__40442\ : std_logic;
signal \N__40441\ : std_logic;
signal \N__40440\ : std_logic;
signal \N__40435\ : std_logic;
signal \N__40432\ : std_logic;
signal \N__40429\ : std_logic;
signal \N__40424\ : std_logic;
signal \N__40421\ : std_logic;
signal \N__40420\ : std_logic;
signal \N__40417\ : std_logic;
signal \N__40414\ : std_logic;
signal \N__40413\ : std_logic;
signal \N__40410\ : std_logic;
signal \N__40407\ : std_logic;
signal \N__40404\ : std_logic;
signal \N__40399\ : std_logic;
signal \N__40394\ : std_logic;
signal \N__40391\ : std_logic;
signal \N__40388\ : std_logic;
signal \N__40387\ : std_logic;
signal \N__40384\ : std_logic;
signal \N__40381\ : std_logic;
signal \N__40378\ : std_logic;
signal \N__40375\ : std_logic;
signal \N__40374\ : std_logic;
signal \N__40371\ : std_logic;
signal \N__40368\ : std_logic;
signal \N__40365\ : std_logic;
signal \N__40360\ : std_logic;
signal \N__40355\ : std_logic;
signal \N__40352\ : std_logic;
signal \N__40349\ : std_logic;
signal \N__40348\ : std_logic;
signal \N__40347\ : std_logic;
signal \N__40344\ : std_logic;
signal \N__40341\ : std_logic;
signal \N__40338\ : std_logic;
signal \N__40335\ : std_logic;
signal \N__40332\ : std_logic;
signal \N__40329\ : std_logic;
signal \N__40328\ : std_logic;
signal \N__40323\ : std_logic;
signal \N__40320\ : std_logic;
signal \N__40317\ : std_logic;
signal \N__40310\ : std_logic;
signal \N__40307\ : std_logic;
signal \N__40304\ : std_logic;
signal \N__40303\ : std_logic;
signal \N__40302\ : std_logic;
signal \N__40297\ : std_logic;
signal \N__40294\ : std_logic;
signal \N__40289\ : std_logic;
signal \N__40288\ : std_logic;
signal \N__40285\ : std_logic;
signal \N__40282\ : std_logic;
signal \N__40277\ : std_logic;
signal \N__40274\ : std_logic;
signal \N__40271\ : std_logic;
signal \N__40268\ : std_logic;
signal \N__40265\ : std_logic;
signal \N__40262\ : std_logic;
signal \N__40261\ : std_logic;
signal \N__40260\ : std_logic;
signal \N__40255\ : std_logic;
signal \N__40252\ : std_logic;
signal \N__40249\ : std_logic;
signal \N__40248\ : std_logic;
signal \N__40245\ : std_logic;
signal \N__40242\ : std_logic;
signal \N__40239\ : std_logic;
signal \N__40232\ : std_logic;
signal \N__40229\ : std_logic;
signal \N__40226\ : std_logic;
signal \N__40223\ : std_logic;
signal \N__40220\ : std_logic;
signal \N__40217\ : std_logic;
signal \N__40214\ : std_logic;
signal \N__40211\ : std_logic;
signal \N__40208\ : std_logic;
signal \N__40205\ : std_logic;
signal \N__40202\ : std_logic;
signal \N__40199\ : std_logic;
signal \N__40196\ : std_logic;
signal \N__40193\ : std_logic;
signal \N__40192\ : std_logic;
signal \N__40191\ : std_logic;
signal \N__40188\ : std_logic;
signal \N__40185\ : std_logic;
signal \N__40182\ : std_logic;
signal \N__40179\ : std_logic;
signal \N__40178\ : std_logic;
signal \N__40175\ : std_logic;
signal \N__40170\ : std_logic;
signal \N__40167\ : std_logic;
signal \N__40160\ : std_logic;
signal \N__40157\ : std_logic;
signal \N__40154\ : std_logic;
signal \N__40153\ : std_logic;
signal \N__40150\ : std_logic;
signal \N__40147\ : std_logic;
signal \N__40146\ : std_logic;
signal \N__40143\ : std_logic;
signal \N__40140\ : std_logic;
signal \N__40137\ : std_logic;
signal \N__40132\ : std_logic;
signal \N__40127\ : std_logic;
signal \N__40124\ : std_logic;
signal \N__40121\ : std_logic;
signal \N__40120\ : std_logic;
signal \N__40117\ : std_logic;
signal \N__40114\ : std_logic;
signal \N__40113\ : std_logic;
signal \N__40110\ : std_logic;
signal \N__40107\ : std_logic;
signal \N__40104\ : std_logic;
signal \N__40101\ : std_logic;
signal \N__40096\ : std_logic;
signal \N__40095\ : std_logic;
signal \N__40090\ : std_logic;
signal \N__40087\ : std_logic;
signal \N__40082\ : std_logic;
signal \N__40079\ : std_logic;
signal \N__40076\ : std_logic;
signal \N__40073\ : std_logic;
signal \N__40072\ : std_logic;
signal \N__40069\ : std_logic;
signal \N__40066\ : std_logic;
signal \N__40065\ : std_logic;
signal \N__40062\ : std_logic;
signal \N__40059\ : std_logic;
signal \N__40056\ : std_logic;
signal \N__40053\ : std_logic;
signal \N__40052\ : std_logic;
signal \N__40049\ : std_logic;
signal \N__40046\ : std_logic;
signal \N__40043\ : std_logic;
signal \N__40040\ : std_logic;
signal \N__40031\ : std_logic;
signal \N__40028\ : std_logic;
signal \N__40025\ : std_logic;
signal \N__40022\ : std_logic;
signal \N__40019\ : std_logic;
signal \N__40018\ : std_logic;
signal \N__40017\ : std_logic;
signal \N__40014\ : std_logic;
signal \N__40011\ : std_logic;
signal \N__40008\ : std_logic;
signal \N__40003\ : std_logic;
signal \N__40000\ : std_logic;
signal \N__39999\ : std_logic;
signal \N__39994\ : std_logic;
signal \N__39991\ : std_logic;
signal \N__39986\ : std_logic;
signal \N__39983\ : std_logic;
signal \N__39980\ : std_logic;
signal \N__39977\ : std_logic;
signal \N__39974\ : std_logic;
signal \N__39971\ : std_logic;
signal \N__39970\ : std_logic;
signal \N__39969\ : std_logic;
signal \N__39966\ : std_logic;
signal \N__39963\ : std_logic;
signal \N__39960\ : std_logic;
signal \N__39957\ : std_logic;
signal \N__39952\ : std_logic;
signal \N__39951\ : std_logic;
signal \N__39946\ : std_logic;
signal \N__39943\ : std_logic;
signal \N__39938\ : std_logic;
signal \N__39935\ : std_logic;
signal \N__39932\ : std_logic;
signal \N__39929\ : std_logic;
signal \N__39926\ : std_logic;
signal \N__39925\ : std_logic;
signal \N__39922\ : std_logic;
signal \N__39919\ : std_logic;
signal \N__39918\ : std_logic;
signal \N__39915\ : std_logic;
signal \N__39912\ : std_logic;
signal \N__39909\ : std_logic;
signal \N__39904\ : std_logic;
signal \N__39901\ : std_logic;
signal \N__39900\ : std_logic;
signal \N__39895\ : std_logic;
signal \N__39892\ : std_logic;
signal \N__39887\ : std_logic;
signal \N__39884\ : std_logic;
signal \N__39881\ : std_logic;
signal \N__39878\ : std_logic;
signal \N__39877\ : std_logic;
signal \N__39876\ : std_logic;
signal \N__39873\ : std_logic;
signal \N__39870\ : std_logic;
signal \N__39867\ : std_logic;
signal \N__39864\ : std_logic;
signal \N__39861\ : std_logic;
signal \N__39860\ : std_logic;
signal \N__39857\ : std_logic;
signal \N__39852\ : std_logic;
signal \N__39849\ : std_logic;
signal \N__39842\ : std_logic;
signal \N__39839\ : std_logic;
signal \N__39836\ : std_logic;
signal \N__39833\ : std_logic;
signal \N__39830\ : std_logic;
signal \N__39827\ : std_logic;
signal \N__39824\ : std_logic;
signal \N__39823\ : std_logic;
signal \N__39822\ : std_logic;
signal \N__39819\ : std_logic;
signal \N__39816\ : std_logic;
signal \N__39813\ : std_logic;
signal \N__39808\ : std_logic;
signal \N__39805\ : std_logic;
signal \N__39804\ : std_logic;
signal \N__39801\ : std_logic;
signal \N__39798\ : std_logic;
signal \N__39795\ : std_logic;
signal \N__39788\ : std_logic;
signal \N__39785\ : std_logic;
signal \N__39782\ : std_logic;
signal \N__39779\ : std_logic;
signal \N__39776\ : std_logic;
signal \N__39773\ : std_logic;
signal \N__39770\ : std_logic;
signal \N__39767\ : std_logic;
signal \N__39764\ : std_logic;
signal \N__39761\ : std_logic;
signal \N__39758\ : std_logic;
signal \N__39757\ : std_logic;
signal \N__39754\ : std_logic;
signal \N__39751\ : std_logic;
signal \N__39750\ : std_logic;
signal \N__39747\ : std_logic;
signal \N__39744\ : std_logic;
signal \N__39741\ : std_logic;
signal \N__39736\ : std_logic;
signal \N__39733\ : std_logic;
signal \N__39728\ : std_logic;
signal \N__39727\ : std_logic;
signal \N__39724\ : std_logic;
signal \N__39721\ : std_logic;
signal \N__39716\ : std_logic;
signal \N__39713\ : std_logic;
signal \N__39710\ : std_logic;
signal \N__39709\ : std_logic;
signal \N__39706\ : std_logic;
signal \N__39703\ : std_logic;
signal \N__39702\ : std_logic;
signal \N__39697\ : std_logic;
signal \N__39694\ : std_logic;
signal \N__39691\ : std_logic;
signal \N__39688\ : std_logic;
signal \N__39687\ : std_logic;
signal \N__39682\ : std_logic;
signal \N__39679\ : std_logic;
signal \N__39674\ : std_logic;
signal \N__39671\ : std_logic;
signal \N__39668\ : std_logic;
signal \N__39665\ : std_logic;
signal \N__39664\ : std_logic;
signal \N__39661\ : std_logic;
signal \N__39660\ : std_logic;
signal \N__39657\ : std_logic;
signal \N__39654\ : std_logic;
signal \N__39651\ : std_logic;
signal \N__39648\ : std_logic;
signal \N__39643\ : std_logic;
signal \N__39642\ : std_logic;
signal \N__39637\ : std_logic;
signal \N__39634\ : std_logic;
signal \N__39629\ : std_logic;
signal \N__39626\ : std_logic;
signal \N__39623\ : std_logic;
signal \N__39620\ : std_logic;
signal \N__39619\ : std_logic;
signal \N__39616\ : std_logic;
signal \N__39615\ : std_logic;
signal \N__39612\ : std_logic;
signal \N__39609\ : std_logic;
signal \N__39606\ : std_logic;
signal \N__39603\ : std_logic;
signal \N__39600\ : std_logic;
signal \N__39597\ : std_logic;
signal \N__39596\ : std_logic;
signal \N__39593\ : std_logic;
signal \N__39588\ : std_logic;
signal \N__39585\ : std_logic;
signal \N__39578\ : std_logic;
signal \N__39575\ : std_logic;
signal \N__39572\ : std_logic;
signal \N__39571\ : std_logic;
signal \N__39568\ : std_logic;
signal \N__39567\ : std_logic;
signal \N__39564\ : std_logic;
signal \N__39561\ : std_logic;
signal \N__39558\ : std_logic;
signal \N__39553\ : std_logic;
signal \N__39552\ : std_logic;
signal \N__39549\ : std_logic;
signal \N__39546\ : std_logic;
signal \N__39543\ : std_logic;
signal \N__39536\ : std_logic;
signal \N__39533\ : std_logic;
signal \N__39530\ : std_logic;
signal \N__39527\ : std_logic;
signal \N__39526\ : std_logic;
signal \N__39525\ : std_logic;
signal \N__39522\ : std_logic;
signal \N__39517\ : std_logic;
signal \N__39516\ : std_logic;
signal \N__39513\ : std_logic;
signal \N__39510\ : std_logic;
signal \N__39507\ : std_logic;
signal \N__39504\ : std_logic;
signal \N__39501\ : std_logic;
signal \N__39494\ : std_logic;
signal \N__39493\ : std_logic;
signal \N__39490\ : std_logic;
signal \N__39489\ : std_logic;
signal \N__39486\ : std_logic;
signal \N__39483\ : std_logic;
signal \N__39480\ : std_logic;
signal \N__39475\ : std_logic;
signal \N__39474\ : std_logic;
signal \N__39471\ : std_logic;
signal \N__39468\ : std_logic;
signal \N__39465\ : std_logic;
signal \N__39458\ : std_logic;
signal \N__39455\ : std_logic;
signal \N__39452\ : std_logic;
signal \N__39449\ : std_logic;
signal \N__39448\ : std_logic;
signal \N__39447\ : std_logic;
signal \N__39444\ : std_logic;
signal \N__39441\ : std_logic;
signal \N__39438\ : std_logic;
signal \N__39435\ : std_logic;
signal \N__39434\ : std_logic;
signal \N__39429\ : std_logic;
signal \N__39426\ : std_logic;
signal \N__39423\ : std_logic;
signal \N__39416\ : std_logic;
signal \N__39413\ : std_logic;
signal \N__39410\ : std_logic;
signal \N__39407\ : std_logic;
signal \N__39406\ : std_logic;
signal \N__39405\ : std_logic;
signal \N__39400\ : std_logic;
signal \N__39397\ : std_logic;
signal \N__39392\ : std_logic;
signal \N__39391\ : std_logic;
signal \N__39388\ : std_logic;
signal \N__39385\ : std_logic;
signal \N__39380\ : std_logic;
signal \N__39377\ : std_logic;
signal \N__39374\ : std_logic;
signal \N__39373\ : std_logic;
signal \N__39370\ : std_logic;
signal \N__39369\ : std_logic;
signal \N__39366\ : std_logic;
signal \N__39363\ : std_logic;
signal \N__39360\ : std_logic;
signal \N__39357\ : std_logic;
signal \N__39354\ : std_logic;
signal \N__39351\ : std_logic;
signal \N__39350\ : std_logic;
signal \N__39343\ : std_logic;
signal \N__39340\ : std_logic;
signal \N__39335\ : std_logic;
signal \N__39332\ : std_logic;
signal \N__39329\ : std_logic;
signal \N__39326\ : std_logic;
signal \N__39325\ : std_logic;
signal \N__39322\ : std_logic;
signal \N__39321\ : std_logic;
signal \N__39316\ : std_logic;
signal \N__39313\ : std_logic;
signal \N__39310\ : std_logic;
signal \N__39307\ : std_logic;
signal \N__39306\ : std_logic;
signal \N__39301\ : std_logic;
signal \N__39298\ : std_logic;
signal \N__39293\ : std_logic;
signal \N__39290\ : std_logic;
signal \N__39287\ : std_logic;
signal \N__39284\ : std_logic;
signal \N__39281\ : std_logic;
signal \N__39280\ : std_logic;
signal \N__39277\ : std_logic;
signal \N__39274\ : std_logic;
signal \N__39273\ : std_logic;
signal \N__39270\ : std_logic;
signal \N__39267\ : std_logic;
signal \N__39266\ : std_logic;
signal \N__39263\ : std_logic;
signal \N__39258\ : std_logic;
signal \N__39255\ : std_logic;
signal \N__39248\ : std_logic;
signal \N__39245\ : std_logic;
signal \N__39242\ : std_logic;
signal \N__39239\ : std_logic;
signal \N__39236\ : std_logic;
signal \N__39235\ : std_logic;
signal \N__39234\ : std_logic;
signal \N__39231\ : std_logic;
signal \N__39228\ : std_logic;
signal \N__39225\ : std_logic;
signal \N__39220\ : std_logic;
signal \N__39215\ : std_logic;
signal \N__39212\ : std_logic;
signal \N__39209\ : std_logic;
signal \N__39208\ : std_logic;
signal \N__39207\ : std_logic;
signal \N__39202\ : std_logic;
signal \N__39199\ : std_logic;
signal \N__39196\ : std_logic;
signal \N__39191\ : std_logic;
signal \N__39188\ : std_logic;
signal \N__39185\ : std_logic;
signal \N__39182\ : std_logic;
signal \N__39179\ : std_logic;
signal \N__39176\ : std_logic;
signal \N__39173\ : std_logic;
signal \N__39170\ : std_logic;
signal \N__39169\ : std_logic;
signal \N__39166\ : std_logic;
signal \N__39165\ : std_logic;
signal \N__39160\ : std_logic;
signal \N__39159\ : std_logic;
signal \N__39156\ : std_logic;
signal \N__39153\ : std_logic;
signal \N__39150\ : std_logic;
signal \N__39147\ : std_logic;
signal \N__39144\ : std_logic;
signal \N__39137\ : std_logic;
signal \N__39134\ : std_logic;
signal \N__39133\ : std_logic;
signal \N__39130\ : std_logic;
signal \N__39127\ : std_logic;
signal \N__39122\ : std_logic;
signal \N__39119\ : std_logic;
signal \N__39118\ : std_logic;
signal \N__39115\ : std_logic;
signal \N__39112\ : std_logic;
signal \N__39107\ : std_logic;
signal \N__39104\ : std_logic;
signal \N__39103\ : std_logic;
signal \N__39100\ : std_logic;
signal \N__39097\ : std_logic;
signal \N__39092\ : std_logic;
signal \N__39089\ : std_logic;
signal \N__39086\ : std_logic;
signal \N__39083\ : std_logic;
signal \N__39080\ : std_logic;
signal \N__39077\ : std_logic;
signal \N__39076\ : std_logic;
signal \N__39073\ : std_logic;
signal \N__39072\ : std_logic;
signal \N__39067\ : std_logic;
signal \N__39064\ : std_logic;
signal \N__39061\ : std_logic;
signal \N__39056\ : std_logic;
signal \N__39053\ : std_logic;
signal \N__39052\ : std_logic;
signal \N__39051\ : std_logic;
signal \N__39046\ : std_logic;
signal \N__39043\ : std_logic;
signal \N__39040\ : std_logic;
signal \N__39035\ : std_logic;
signal \N__39032\ : std_logic;
signal \N__39031\ : std_logic;
signal \N__39028\ : std_logic;
signal \N__39025\ : std_logic;
signal \N__39020\ : std_logic;
signal \N__39017\ : std_logic;
signal \N__39016\ : std_logic;
signal \N__39013\ : std_logic;
signal \N__39010\ : std_logic;
signal \N__39005\ : std_logic;
signal \N__39002\ : std_logic;
signal \N__39001\ : std_logic;
signal \N__38998\ : std_logic;
signal \N__38995\ : std_logic;
signal \N__38990\ : std_logic;
signal \N__38987\ : std_logic;
signal \N__38986\ : std_logic;
signal \N__38983\ : std_logic;
signal \N__38980\ : std_logic;
signal \N__38975\ : std_logic;
signal \N__38972\ : std_logic;
signal \N__38971\ : std_logic;
signal \N__38968\ : std_logic;
signal \N__38965\ : std_logic;
signal \N__38960\ : std_logic;
signal \N__38957\ : std_logic;
signal \N__38956\ : std_logic;
signal \N__38953\ : std_logic;
signal \N__38950\ : std_logic;
signal \N__38945\ : std_logic;
signal \N__38942\ : std_logic;
signal \N__38941\ : std_logic;
signal \N__38938\ : std_logic;
signal \N__38935\ : std_logic;
signal \N__38930\ : std_logic;
signal \N__38927\ : std_logic;
signal \N__38926\ : std_logic;
signal \N__38923\ : std_logic;
signal \N__38920\ : std_logic;
signal \N__38915\ : std_logic;
signal \N__38912\ : std_logic;
signal \N__38911\ : std_logic;
signal \N__38910\ : std_logic;
signal \N__38907\ : std_logic;
signal \N__38904\ : std_logic;
signal \N__38903\ : std_logic;
signal \N__38900\ : std_logic;
signal \N__38897\ : std_logic;
signal \N__38894\ : std_logic;
signal \N__38891\ : std_logic;
signal \N__38888\ : std_logic;
signal \N__38885\ : std_logic;
signal \N__38880\ : std_logic;
signal \N__38877\ : std_logic;
signal \N__38874\ : std_logic;
signal \N__38867\ : std_logic;
signal \N__38866\ : std_logic;
signal \N__38865\ : std_logic;
signal \N__38862\ : std_logic;
signal \N__38859\ : std_logic;
signal \N__38856\ : std_logic;
signal \N__38851\ : std_logic;
signal \N__38846\ : std_logic;
signal \N__38843\ : std_logic;
signal \N__38842\ : std_logic;
signal \N__38841\ : std_logic;
signal \N__38838\ : std_logic;
signal \N__38833\ : std_logic;
signal \N__38830\ : std_logic;
signal \N__38825\ : std_logic;
signal \N__38824\ : std_logic;
signal \N__38821\ : std_logic;
signal \N__38818\ : std_logic;
signal \N__38817\ : std_logic;
signal \N__38814\ : std_logic;
signal \N__38809\ : std_logic;
signal \N__38806\ : std_logic;
signal \N__38801\ : std_logic;
signal \N__38798\ : std_logic;
signal \N__38797\ : std_logic;
signal \N__38796\ : std_logic;
signal \N__38795\ : std_logic;
signal \N__38792\ : std_logic;
signal \N__38789\ : std_logic;
signal \N__38786\ : std_logic;
signal \N__38783\ : std_logic;
signal \N__38780\ : std_logic;
signal \N__38773\ : std_logic;
signal \N__38770\ : std_logic;
signal \N__38767\ : std_logic;
signal \N__38762\ : std_logic;
signal \N__38759\ : std_logic;
signal \N__38758\ : std_logic;
signal \N__38755\ : std_logic;
signal \N__38754\ : std_logic;
signal \N__38751\ : std_logic;
signal \N__38748\ : std_logic;
signal \N__38745\ : std_logic;
signal \N__38738\ : std_logic;
signal \N__38737\ : std_logic;
signal \N__38736\ : std_logic;
signal \N__38735\ : std_logic;
signal \N__38732\ : std_logic;
signal \N__38729\ : std_logic;
signal \N__38726\ : std_logic;
signal \N__38723\ : std_logic;
signal \N__38718\ : std_logic;
signal \N__38715\ : std_logic;
signal \N__38712\ : std_logic;
signal \N__38709\ : std_logic;
signal \N__38706\ : std_logic;
signal \N__38699\ : std_logic;
signal \N__38698\ : std_logic;
signal \N__38697\ : std_logic;
signal \N__38694\ : std_logic;
signal \N__38691\ : std_logic;
signal \N__38688\ : std_logic;
signal \N__38681\ : std_logic;
signal \N__38678\ : std_logic;
signal \N__38675\ : std_logic;
signal \N__38674\ : std_logic;
signal \N__38671\ : std_logic;
signal \N__38670\ : std_logic;
signal \N__38667\ : std_logic;
signal \N__38664\ : std_logic;
signal \N__38661\ : std_logic;
signal \N__38658\ : std_logic;
signal \N__38653\ : std_logic;
signal \N__38648\ : std_logic;
signal \N__38647\ : std_logic;
signal \N__38644\ : std_logic;
signal \N__38641\ : std_logic;
signal \N__38636\ : std_logic;
signal \N__38633\ : std_logic;
signal \N__38632\ : std_logic;
signal \N__38629\ : std_logic;
signal \N__38626\ : std_logic;
signal \N__38621\ : std_logic;
signal \N__38618\ : std_logic;
signal \N__38617\ : std_logic;
signal \N__38614\ : std_logic;
signal \N__38611\ : std_logic;
signal \N__38606\ : std_logic;
signal \N__38603\ : std_logic;
signal \N__38600\ : std_logic;
signal \N__38597\ : std_logic;
signal \N__38594\ : std_logic;
signal \N__38591\ : std_logic;
signal \N__38588\ : std_logic;
signal \N__38585\ : std_logic;
signal \N__38582\ : std_logic;
signal \N__38579\ : std_logic;
signal \N__38576\ : std_logic;
signal \N__38573\ : std_logic;
signal \N__38570\ : std_logic;
signal \N__38567\ : std_logic;
signal \N__38564\ : std_logic;
signal \N__38561\ : std_logic;
signal \N__38558\ : std_logic;
signal \N__38557\ : std_logic;
signal \N__38554\ : std_logic;
signal \N__38551\ : std_logic;
signal \N__38546\ : std_logic;
signal \N__38543\ : std_logic;
signal \N__38542\ : std_logic;
signal \N__38537\ : std_logic;
signal \N__38534\ : std_logic;
signal \N__38531\ : std_logic;
signal \N__38528\ : std_logic;
signal \N__38525\ : std_logic;
signal \N__38522\ : std_logic;
signal \N__38521\ : std_logic;
signal \N__38520\ : std_logic;
signal \N__38517\ : std_logic;
signal \N__38514\ : std_logic;
signal \N__38511\ : std_logic;
signal \N__38508\ : std_logic;
signal \N__38501\ : std_logic;
signal \N__38500\ : std_logic;
signal \N__38499\ : std_logic;
signal \N__38498\ : std_logic;
signal \N__38495\ : std_logic;
signal \N__38490\ : std_logic;
signal \N__38487\ : std_logic;
signal \N__38482\ : std_logic;
signal \N__38479\ : std_logic;
signal \N__38476\ : std_logic;
signal \N__38471\ : std_logic;
signal \N__38468\ : std_logic;
signal \N__38465\ : std_logic;
signal \N__38462\ : std_logic;
signal \N__38459\ : std_logic;
signal \N__38458\ : std_logic;
signal \N__38457\ : std_logic;
signal \N__38454\ : std_logic;
signal \N__38451\ : std_logic;
signal \N__38448\ : std_logic;
signal \N__38445\ : std_logic;
signal \N__38444\ : std_logic;
signal \N__38439\ : std_logic;
signal \N__38436\ : std_logic;
signal \N__38433\ : std_logic;
signal \N__38428\ : std_logic;
signal \N__38423\ : std_logic;
signal \N__38420\ : std_logic;
signal \N__38417\ : std_logic;
signal \N__38414\ : std_logic;
signal \N__38413\ : std_logic;
signal \N__38410\ : std_logic;
signal \N__38407\ : std_logic;
signal \N__38402\ : std_logic;
signal \N__38399\ : std_logic;
signal \N__38396\ : std_logic;
signal \N__38395\ : std_logic;
signal \N__38390\ : std_logic;
signal \N__38387\ : std_logic;
signal \N__38384\ : std_logic;
signal \N__38381\ : std_logic;
signal \N__38378\ : std_logic;
signal \N__38375\ : std_logic;
signal \N__38372\ : std_logic;
signal \N__38369\ : std_logic;
signal \N__38366\ : std_logic;
signal \N__38363\ : std_logic;
signal \N__38360\ : std_logic;
signal \N__38357\ : std_logic;
signal \N__38356\ : std_logic;
signal \N__38353\ : std_logic;
signal \N__38350\ : std_logic;
signal \N__38347\ : std_logic;
signal \N__38344\ : std_logic;
signal \N__38343\ : std_logic;
signal \N__38342\ : std_logic;
signal \N__38339\ : std_logic;
signal \N__38336\ : std_logic;
signal \N__38331\ : std_logic;
signal \N__38328\ : std_logic;
signal \N__38321\ : std_logic;
signal \N__38318\ : std_logic;
signal \N__38315\ : std_logic;
signal \N__38312\ : std_logic;
signal \N__38309\ : std_logic;
signal \N__38308\ : std_logic;
signal \N__38305\ : std_logic;
signal \N__38302\ : std_logic;
signal \N__38301\ : std_logic;
signal \N__38300\ : std_logic;
signal \N__38295\ : std_logic;
signal \N__38292\ : std_logic;
signal \N__38289\ : std_logic;
signal \N__38286\ : std_logic;
signal \N__38283\ : std_logic;
signal \N__38280\ : std_logic;
signal \N__38277\ : std_logic;
signal \N__38272\ : std_logic;
signal \N__38267\ : std_logic;
signal \N__38266\ : std_logic;
signal \N__38265\ : std_logic;
signal \N__38264\ : std_logic;
signal \N__38259\ : std_logic;
signal \N__38256\ : std_logic;
signal \N__38253\ : std_logic;
signal \N__38250\ : std_logic;
signal \N__38247\ : std_logic;
signal \N__38244\ : std_logic;
signal \N__38241\ : std_logic;
signal \N__38236\ : std_logic;
signal \N__38231\ : std_logic;
signal \N__38228\ : std_logic;
signal \N__38227\ : std_logic;
signal \N__38224\ : std_logic;
signal \N__38221\ : std_logic;
signal \N__38218\ : std_logic;
signal \N__38217\ : std_logic;
signal \N__38214\ : std_logic;
signal \N__38213\ : std_logic;
signal \N__38210\ : std_logic;
signal \N__38207\ : std_logic;
signal \N__38204\ : std_logic;
signal \N__38201\ : std_logic;
signal \N__38192\ : std_logic;
signal \N__38191\ : std_logic;
signal \N__38188\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38184\ : std_logic;
signal \N__38181\ : std_logic;
signal \N__38178\ : std_logic;
signal \N__38175\ : std_logic;
signal \N__38170\ : std_logic;
signal \N__38165\ : std_logic;
signal \N__38162\ : std_logic;
signal \N__38161\ : std_logic;
signal \N__38160\ : std_logic;
signal \N__38159\ : std_logic;
signal \N__38156\ : std_logic;
signal \N__38153\ : std_logic;
signal \N__38150\ : std_logic;
signal \N__38147\ : std_logic;
signal \N__38144\ : std_logic;
signal \N__38141\ : std_logic;
signal \N__38138\ : std_logic;
signal \N__38135\ : std_logic;
signal \N__38132\ : std_logic;
signal \N__38127\ : std_logic;
signal \N__38120\ : std_logic;
signal \N__38119\ : std_logic;
signal \N__38118\ : std_logic;
signal \N__38115\ : std_logic;
signal \N__38112\ : std_logic;
signal \N__38109\ : std_logic;
signal \N__38106\ : std_logic;
signal \N__38099\ : std_logic;
signal \N__38098\ : std_logic;
signal \N__38097\ : std_logic;
signal \N__38094\ : std_logic;
signal \N__38091\ : std_logic;
signal \N__38088\ : std_logic;
signal \N__38081\ : std_logic;
signal \N__38080\ : std_logic;
signal \N__38079\ : std_logic;
signal \N__38076\ : std_logic;
signal \N__38073\ : std_logic;
signal \N__38070\ : std_logic;
signal \N__38067\ : std_logic;
signal \N__38060\ : std_logic;
signal \N__38057\ : std_logic;
signal \N__38056\ : std_logic;
signal \N__38055\ : std_logic;
signal \N__38050\ : std_logic;
signal \N__38047\ : std_logic;
signal \N__38046\ : std_logic;
signal \N__38043\ : std_logic;
signal \N__38040\ : std_logic;
signal \N__38037\ : std_logic;
signal \N__38034\ : std_logic;
signal \N__38031\ : std_logic;
signal \N__38024\ : std_logic;
signal \N__38021\ : std_logic;
signal \N__38020\ : std_logic;
signal \N__38017\ : std_logic;
signal \N__38014\ : std_logic;
signal \N__38011\ : std_logic;
signal \N__38008\ : std_logic;
signal \N__38003\ : std_logic;
signal \N__38002\ : std_logic;
signal \N__38001\ : std_logic;
signal \N__38000\ : std_logic;
signal \N__37999\ : std_logic;
signal \N__37998\ : std_logic;
signal \N__37997\ : std_logic;
signal \N__37996\ : std_logic;
signal \N__37995\ : std_logic;
signal \N__37994\ : std_logic;
signal \N__37993\ : std_logic;
signal \N__37992\ : std_logic;
signal \N__37991\ : std_logic;
signal \N__37990\ : std_logic;
signal \N__37987\ : std_logic;
signal \N__37984\ : std_logic;
signal \N__37981\ : std_logic;
signal \N__37980\ : std_logic;
signal \N__37979\ : std_logic;
signal \N__37978\ : std_logic;
signal \N__37977\ : std_logic;
signal \N__37976\ : std_logic;
signal \N__37975\ : std_logic;
signal \N__37972\ : std_logic;
signal \N__37971\ : std_logic;
signal \N__37968\ : std_logic;
signal \N__37967\ : std_logic;
signal \N__37964\ : std_logic;
signal \N__37963\ : std_logic;
signal \N__37960\ : std_logic;
signal \N__37959\ : std_logic;
signal \N__37956\ : std_logic;
signal \N__37955\ : std_logic;
signal \N__37952\ : std_logic;
signal \N__37951\ : std_logic;
signal \N__37948\ : std_logic;
signal \N__37947\ : std_logic;
signal \N__37944\ : std_logic;
signal \N__37943\ : std_logic;
signal \N__37940\ : std_logic;
signal \N__37939\ : std_logic;
signal \N__37936\ : std_logic;
signal \N__37935\ : std_logic;
signal \N__37932\ : std_logic;
signal \N__37931\ : std_logic;
signal \N__37930\ : std_logic;
signal \N__37929\ : std_logic;
signal \N__37928\ : std_logic;
signal \N__37921\ : std_logic;
signal \N__37918\ : std_logic;
signal \N__37917\ : std_logic;
signal \N__37914\ : std_logic;
signal \N__37909\ : std_logic;
signal \N__37906\ : std_logic;
signal \N__37905\ : std_logic;
signal \N__37904\ : std_logic;
signal \N__37903\ : std_logic;
signal \N__37902\ : std_logic;
signal \N__37901\ : std_logic;
signal \N__37900\ : std_logic;
signal \N__37899\ : std_logic;
signal \N__37898\ : std_logic;
signal \N__37897\ : std_logic;
signal \N__37894\ : std_logic;
signal \N__37879\ : std_logic;
signal \N__37864\ : std_logic;
signal \N__37847\ : std_logic;
signal \N__37846\ : std_logic;
signal \N__37845\ : std_logic;
signal \N__37844\ : std_logic;
signal \N__37843\ : std_logic;
signal \N__37840\ : std_logic;
signal \N__37835\ : std_logic;
signal \N__37830\ : std_logic;
signal \N__37829\ : std_logic;
signal \N__37828\ : std_logic;
signal \N__37827\ : std_logic;
signal \N__37826\ : std_logic;
signal \N__37825\ : std_logic;
signal \N__37824\ : std_logic;
signal \N__37823\ : std_logic;
signal \N__37822\ : std_logic;
signal \N__37819\ : std_logic;
signal \N__37818\ : std_logic;
signal \N__37815\ : std_logic;
signal \N__37810\ : std_logic;
signal \N__37807\ : std_logic;
signal \N__37804\ : std_logic;
signal \N__37797\ : std_logic;
signal \N__37788\ : std_logic;
signal \N__37785\ : std_logic;
signal \N__37782\ : std_logic;
signal \N__37777\ : std_logic;
signal \N__37774\ : std_logic;
signal \N__37773\ : std_logic;
signal \N__37770\ : std_logic;
signal \N__37769\ : std_logic;
signal \N__37766\ : std_logic;
signal \N__37765\ : std_logic;
signal \N__37762\ : std_logic;
signal \N__37761\ : std_logic;
signal \N__37760\ : std_logic;
signal \N__37759\ : std_logic;
signal \N__37756\ : std_logic;
signal \N__37753\ : std_logic;
signal \N__37750\ : std_logic;
signal \N__37743\ : std_logic;
signal \N__37734\ : std_logic;
signal \N__37727\ : std_logic;
signal \N__37720\ : std_logic;
signal \N__37711\ : std_logic;
signal \N__37706\ : std_logic;
signal \N__37689\ : std_logic;
signal \N__37684\ : std_logic;
signal \N__37679\ : std_logic;
signal \N__37670\ : std_logic;
signal \N__37667\ : std_logic;
signal \N__37660\ : std_logic;
signal \N__37657\ : std_logic;
signal \N__37654\ : std_logic;
signal \N__37651\ : std_logic;
signal \N__37644\ : std_logic;
signal \N__37637\ : std_logic;
signal \N__37634\ : std_logic;
signal \N__37633\ : std_logic;
signal \N__37632\ : std_logic;
signal \N__37631\ : std_logic;
signal \N__37628\ : std_logic;
signal \N__37625\ : std_logic;
signal \N__37624\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37622\ : std_logic;
signal \N__37621\ : std_logic;
signal \N__37616\ : std_logic;
signal \N__37613\ : std_logic;
signal \N__37610\ : std_logic;
signal \N__37607\ : std_logic;
signal \N__37602\ : std_logic;
signal \N__37601\ : std_logic;
signal \N__37600\ : std_logic;
signal \N__37599\ : std_logic;
signal \N__37598\ : std_logic;
signal \N__37595\ : std_logic;
signal \N__37594\ : std_logic;
signal \N__37593\ : std_logic;
signal \N__37590\ : std_logic;
signal \N__37589\ : std_logic;
signal \N__37586\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37578\ : std_logic;
signal \N__37563\ : std_logic;
signal \N__37560\ : std_logic;
signal \N__37557\ : std_logic;
signal \N__37552\ : std_logic;
signal \N__37547\ : std_logic;
signal \N__37544\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37532\ : std_logic;
signal \N__37529\ : std_logic;
signal \N__37526\ : std_logic;
signal \N__37523\ : std_logic;
signal \N__37520\ : std_logic;
signal \N__37517\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37511\ : std_logic;
signal \N__37508\ : std_logic;
signal \N__37505\ : std_logic;
signal \N__37502\ : std_logic;
signal \N__37501\ : std_logic;
signal \N__37498\ : std_logic;
signal \N__37495\ : std_logic;
signal \N__37492\ : std_logic;
signal \N__37487\ : std_logic;
signal \N__37484\ : std_logic;
signal \N__37481\ : std_logic;
signal \N__37478\ : std_logic;
signal \N__37475\ : std_logic;
signal \N__37472\ : std_logic;
signal \N__37469\ : std_logic;
signal \N__37466\ : std_logic;
signal \N__37463\ : std_logic;
signal \N__37460\ : std_logic;
signal \N__37457\ : std_logic;
signal \N__37454\ : std_logic;
signal \N__37451\ : std_logic;
signal \N__37448\ : std_logic;
signal \N__37445\ : std_logic;
signal \N__37442\ : std_logic;
signal \N__37439\ : std_logic;
signal \N__37436\ : std_logic;
signal \N__37433\ : std_logic;
signal \N__37430\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37421\ : std_logic;
signal \N__37418\ : std_logic;
signal \N__37415\ : std_logic;
signal \N__37412\ : std_logic;
signal \N__37409\ : std_logic;
signal \N__37406\ : std_logic;
signal \N__37403\ : std_logic;
signal \N__37400\ : std_logic;
signal \N__37397\ : std_logic;
signal \N__37394\ : std_logic;
signal \N__37391\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37385\ : std_logic;
signal \N__37382\ : std_logic;
signal \N__37379\ : std_logic;
signal \N__37376\ : std_logic;
signal \N__37373\ : std_logic;
signal \N__37370\ : std_logic;
signal \N__37367\ : std_logic;
signal \N__37364\ : std_logic;
signal \N__37361\ : std_logic;
signal \N__37358\ : std_logic;
signal \N__37355\ : std_logic;
signal \N__37352\ : std_logic;
signal \N__37349\ : std_logic;
signal \N__37346\ : std_logic;
signal \N__37343\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37334\ : std_logic;
signal \N__37331\ : std_logic;
signal \N__37328\ : std_logic;
signal \N__37325\ : std_logic;
signal \N__37322\ : std_logic;
signal \N__37321\ : std_logic;
signal \N__37316\ : std_logic;
signal \N__37313\ : std_logic;
signal \N__37310\ : std_logic;
signal \N__37309\ : std_logic;
signal \N__37306\ : std_logic;
signal \N__37305\ : std_logic;
signal \N__37302\ : std_logic;
signal \N__37299\ : std_logic;
signal \N__37296\ : std_logic;
signal \N__37289\ : std_logic;
signal \N__37286\ : std_logic;
signal \N__37283\ : std_logic;
signal \N__37282\ : std_logic;
signal \N__37281\ : std_logic;
signal \N__37280\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37274\ : std_logic;
signal \N__37269\ : std_logic;
signal \N__37262\ : std_logic;
signal \N__37261\ : std_logic;
signal \N__37260\ : std_logic;
signal \N__37257\ : std_logic;
signal \N__37254\ : std_logic;
signal \N__37251\ : std_logic;
signal \N__37248\ : std_logic;
signal \N__37247\ : std_logic;
signal \N__37244\ : std_logic;
signal \N__37241\ : std_logic;
signal \N__37238\ : std_logic;
signal \N__37235\ : std_logic;
signal \N__37230\ : std_logic;
signal \N__37227\ : std_logic;
signal \N__37220\ : std_logic;
signal \N__37217\ : std_logic;
signal \N__37216\ : std_logic;
signal \N__37213\ : std_logic;
signal \N__37212\ : std_logic;
signal \N__37209\ : std_logic;
signal \N__37206\ : std_logic;
signal \N__37203\ : std_logic;
signal \N__37198\ : std_logic;
signal \N__37193\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37184\ : std_logic;
signal \N__37181\ : std_logic;
signal \N__37178\ : std_logic;
signal \N__37175\ : std_logic;
signal \N__37172\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37166\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37157\ : std_logic;
signal \N__37154\ : std_logic;
signal \N__37151\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37145\ : std_logic;
signal \N__37142\ : std_logic;
signal \N__37139\ : std_logic;
signal \N__37136\ : std_logic;
signal \N__37133\ : std_logic;
signal \N__37130\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37121\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37115\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37109\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37103\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37097\ : std_logic;
signal \N__37096\ : std_logic;
signal \N__37093\ : std_logic;
signal \N__37090\ : std_logic;
signal \N__37085\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37078\ : std_logic;
signal \N__37075\ : std_logic;
signal \N__37072\ : std_logic;
signal \N__37067\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37061\ : std_logic;
signal \N__37060\ : std_logic;
signal \N__37059\ : std_logic;
signal \N__37058\ : std_logic;
signal \N__37055\ : std_logic;
signal \N__37048\ : std_logic;
signal \N__37043\ : std_logic;
signal \N__37040\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37034\ : std_logic;
signal \N__37033\ : std_logic;
signal \N__37032\ : std_logic;
signal \N__37031\ : std_logic;
signal \N__37028\ : std_logic;
signal \N__37021\ : std_logic;
signal \N__37016\ : std_logic;
signal \N__37015\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__37001\ : std_logic;
signal \N__36998\ : std_logic;
signal \N__36995\ : std_logic;
signal \N__36992\ : std_logic;
signal \N__36989\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36976\ : std_logic;
signal \N__36971\ : std_logic;
signal \N__36970\ : std_logic;
signal \N__36967\ : std_logic;
signal \N__36964\ : std_logic;
signal \N__36961\ : std_logic;
signal \N__36956\ : std_logic;
signal \N__36953\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36947\ : std_logic;
signal \N__36946\ : std_logic;
signal \N__36943\ : std_logic;
signal \N__36940\ : std_logic;
signal \N__36937\ : std_logic;
signal \N__36932\ : std_logic;
signal \N__36929\ : std_logic;
signal \N__36926\ : std_logic;
signal \N__36925\ : std_logic;
signal \N__36920\ : std_logic;
signal \N__36917\ : std_logic;
signal \N__36914\ : std_logic;
signal \N__36913\ : std_logic;
signal \N__36908\ : std_logic;
signal \N__36905\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36899\ : std_logic;
signal \N__36896\ : std_logic;
signal \N__36893\ : std_logic;
signal \N__36890\ : std_logic;
signal \N__36889\ : std_logic;
signal \N__36888\ : std_logic;
signal \N__36885\ : std_logic;
signal \N__36880\ : std_logic;
signal \N__36875\ : std_logic;
signal \N__36872\ : std_logic;
signal \N__36869\ : std_logic;
signal \N__36866\ : std_logic;
signal \N__36863\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36859\ : std_logic;
signal \N__36856\ : std_logic;
signal \N__36851\ : std_logic;
signal \N__36848\ : std_logic;
signal \N__36845\ : std_logic;
signal \N__36842\ : std_logic;
signal \N__36839\ : std_logic;
signal \N__36836\ : std_logic;
signal \N__36835\ : std_logic;
signal \N__36830\ : std_logic;
signal \N__36829\ : std_logic;
signal \N__36826\ : std_logic;
signal \N__36823\ : std_logic;
signal \N__36820\ : std_logic;
signal \N__36815\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36811\ : std_logic;
signal \N__36808\ : std_logic;
signal \N__36805\ : std_logic;
signal \N__36802\ : std_logic;
signal \N__36801\ : std_logic;
signal \N__36796\ : std_logic;
signal \N__36793\ : std_logic;
signal \N__36790\ : std_logic;
signal \N__36785\ : std_logic;
signal \N__36784\ : std_logic;
signal \N__36781\ : std_logic;
signal \N__36778\ : std_logic;
signal \N__36773\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36764\ : std_logic;
signal \N__36761\ : std_logic;
signal \N__36758\ : std_logic;
signal \N__36755\ : std_logic;
signal \N__36752\ : std_logic;
signal \N__36749\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36740\ : std_logic;
signal \N__36739\ : std_logic;
signal \N__36736\ : std_logic;
signal \N__36733\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36721\ : std_logic;
signal \N__36718\ : std_logic;
signal \N__36715\ : std_logic;
signal \N__36710\ : std_logic;
signal \N__36709\ : std_logic;
signal \N__36704\ : std_logic;
signal \N__36703\ : std_logic;
signal \N__36700\ : std_logic;
signal \N__36697\ : std_logic;
signal \N__36696\ : std_logic;
signal \N__36695\ : std_logic;
signal \N__36694\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36690\ : std_logic;
signal \N__36687\ : std_logic;
signal \N__36684\ : std_logic;
signal \N__36679\ : std_logic;
signal \N__36678\ : std_logic;
signal \N__36675\ : std_logic;
signal \N__36672\ : std_logic;
signal \N__36669\ : std_logic;
signal \N__36664\ : std_logic;
signal \N__36661\ : std_logic;
signal \N__36650\ : std_logic;
signal \N__36649\ : std_logic;
signal \N__36646\ : std_logic;
signal \N__36643\ : std_logic;
signal \N__36640\ : std_logic;
signal \N__36637\ : std_logic;
signal \N__36636\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36634\ : std_logic;
signal \N__36631\ : std_logic;
signal \N__36628\ : std_logic;
signal \N__36625\ : std_logic;
signal \N__36622\ : std_logic;
signal \N__36619\ : std_logic;
signal \N__36608\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36602\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36598\ : std_logic;
signal \N__36595\ : std_logic;
signal \N__36592\ : std_logic;
signal \N__36587\ : std_logic;
signal \N__36586\ : std_logic;
signal \N__36583\ : std_logic;
signal \N__36580\ : std_logic;
signal \N__36579\ : std_logic;
signal \N__36578\ : std_logic;
signal \N__36577\ : std_logic;
signal \N__36576\ : std_logic;
signal \N__36571\ : std_logic;
signal \N__36568\ : std_logic;
signal \N__36565\ : std_logic;
signal \N__36560\ : std_logic;
signal \N__36555\ : std_logic;
signal \N__36552\ : std_logic;
signal \N__36545\ : std_logic;
signal \N__36542\ : std_logic;
signal \N__36539\ : std_logic;
signal \N__36536\ : std_logic;
signal \N__36535\ : std_logic;
signal \N__36532\ : std_logic;
signal \N__36529\ : std_logic;
signal \N__36524\ : std_logic;
signal \N__36521\ : std_logic;
signal \N__36518\ : std_logic;
signal \N__36515\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36509\ : std_logic;
signal \N__36506\ : std_logic;
signal \N__36503\ : std_logic;
signal \N__36500\ : std_logic;
signal \N__36497\ : std_logic;
signal \N__36494\ : std_logic;
signal \N__36491\ : std_logic;
signal \N__36488\ : std_logic;
signal \N__36485\ : std_logic;
signal \N__36482\ : std_logic;
signal \N__36479\ : std_logic;
signal \N__36476\ : std_logic;
signal \N__36473\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36467\ : std_logic;
signal \N__36464\ : std_logic;
signal \N__36461\ : std_logic;
signal \N__36458\ : std_logic;
signal \N__36455\ : std_logic;
signal \N__36452\ : std_logic;
signal \N__36449\ : std_logic;
signal \N__36446\ : std_logic;
signal \N__36443\ : std_logic;
signal \N__36440\ : std_logic;
signal \N__36437\ : std_logic;
signal \N__36434\ : std_logic;
signal \N__36431\ : std_logic;
signal \N__36428\ : std_logic;
signal \N__36425\ : std_logic;
signal \N__36422\ : std_logic;
signal \N__36419\ : std_logic;
signal \N__36416\ : std_logic;
signal \N__36413\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36404\ : std_logic;
signal \N__36401\ : std_logic;
signal \N__36398\ : std_logic;
signal \N__36395\ : std_logic;
signal \N__36392\ : std_logic;
signal \N__36389\ : std_logic;
signal \N__36386\ : std_logic;
signal \N__36383\ : std_logic;
signal \N__36380\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36374\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36368\ : std_logic;
signal \N__36365\ : std_logic;
signal \N__36362\ : std_logic;
signal \N__36359\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36353\ : std_logic;
signal \N__36350\ : std_logic;
signal \N__36347\ : std_logic;
signal \N__36344\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36335\ : std_logic;
signal \N__36332\ : std_logic;
signal \N__36329\ : std_logic;
signal \N__36326\ : std_logic;
signal \N__36323\ : std_logic;
signal \N__36320\ : std_logic;
signal \N__36317\ : std_logic;
signal \N__36314\ : std_logic;
signal \N__36311\ : std_logic;
signal \N__36308\ : std_logic;
signal \N__36305\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36299\ : std_logic;
signal \N__36296\ : std_logic;
signal \N__36293\ : std_logic;
signal \N__36290\ : std_logic;
signal \N__36287\ : std_logic;
signal \N__36286\ : std_logic;
signal \N__36283\ : std_logic;
signal \N__36280\ : std_logic;
signal \N__36279\ : std_logic;
signal \N__36276\ : std_logic;
signal \N__36273\ : std_logic;
signal \N__36270\ : std_logic;
signal \N__36267\ : std_logic;
signal \N__36264\ : std_logic;
signal \N__36257\ : std_logic;
signal \N__36254\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36250\ : std_logic;
signal \N__36247\ : std_logic;
signal \N__36244\ : std_logic;
signal \N__36239\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36234\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36228\ : std_logic;
signal \N__36225\ : std_logic;
signal \N__36218\ : std_logic;
signal \N__36215\ : std_logic;
signal \N__36212\ : std_logic;
signal \N__36211\ : std_logic;
signal \N__36208\ : std_logic;
signal \N__36205\ : std_logic;
signal \N__36202\ : std_logic;
signal \N__36197\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36192\ : std_logic;
signal \N__36189\ : std_logic;
signal \N__36186\ : std_logic;
signal \N__36183\ : std_logic;
signal \N__36178\ : std_logic;
signal \N__36173\ : std_logic;
signal \N__36170\ : std_logic;
signal \N__36167\ : std_logic;
signal \N__36166\ : std_logic;
signal \N__36163\ : std_logic;
signal \N__36160\ : std_logic;
signal \N__36159\ : std_logic;
signal \N__36158\ : std_logic;
signal \N__36157\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36148\ : std_logic;
signal \N__36145\ : std_logic;
signal \N__36142\ : std_logic;
signal \N__36139\ : std_logic;
signal \N__36136\ : std_logic;
signal \N__36133\ : std_logic;
signal \N__36130\ : std_logic;
signal \N__36127\ : std_logic;
signal \N__36124\ : std_logic;
signal \N__36119\ : std_logic;
signal \N__36116\ : std_logic;
signal \N__36113\ : std_logic;
signal \N__36108\ : std_logic;
signal \N__36103\ : std_logic;
signal \N__36098\ : std_logic;
signal \N__36095\ : std_logic;
signal \N__36092\ : std_logic;
signal \N__36089\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36083\ : std_logic;
signal \N__36080\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36074\ : std_logic;
signal \N__36071\ : std_logic;
signal \N__36068\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36056\ : std_logic;
signal \N__36053\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36040\ : std_logic;
signal \N__36037\ : std_logic;
signal \N__36034\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36030\ : std_logic;
signal \N__36027\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36021\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36008\ : std_logic;
signal \N__36005\ : std_logic;
signal \N__36002\ : std_logic;
signal \N__36001\ : std_logic;
signal \N__36000\ : std_logic;
signal \N__35997\ : std_logic;
signal \N__35994\ : std_logic;
signal \N__35991\ : std_logic;
signal \N__35984\ : std_logic;
signal \N__35981\ : std_logic;
signal \N__35978\ : std_logic;
signal \N__35977\ : std_logic;
signal \N__35976\ : std_logic;
signal \N__35971\ : std_logic;
signal \N__35968\ : std_logic;
signal \N__35965\ : std_logic;
signal \N__35960\ : std_logic;
signal \N__35957\ : std_logic;
signal \N__35956\ : std_logic;
signal \N__35955\ : std_logic;
signal \N__35950\ : std_logic;
signal \N__35947\ : std_logic;
signal \N__35944\ : std_logic;
signal \N__35939\ : std_logic;
signal \N__35936\ : std_logic;
signal \N__35935\ : std_logic;
signal \N__35932\ : std_logic;
signal \N__35931\ : std_logic;
signal \N__35928\ : std_logic;
signal \N__35925\ : std_logic;
signal \N__35922\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35912\ : std_logic;
signal \N__35909\ : std_logic;
signal \N__35908\ : std_logic;
signal \N__35905\ : std_logic;
signal \N__35902\ : std_logic;
signal \N__35901\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35893\ : std_logic;
signal \N__35890\ : std_logic;
signal \N__35885\ : std_logic;
signal \N__35882\ : std_logic;
signal \N__35881\ : std_logic;
signal \N__35878\ : std_logic;
signal \N__35875\ : std_logic;
signal \N__35874\ : std_logic;
signal \N__35869\ : std_logic;
signal \N__35866\ : std_logic;
signal \N__35863\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35852\ : std_logic;
signal \N__35851\ : std_logic;
signal \N__35848\ : std_logic;
signal \N__35845\ : std_logic;
signal \N__35844\ : std_logic;
signal \N__35839\ : std_logic;
signal \N__35836\ : std_logic;
signal \N__35833\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35825\ : std_logic;
signal \N__35824\ : std_logic;
signal \N__35823\ : std_logic;
signal \N__35820\ : std_logic;
signal \N__35817\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35808\ : std_logic;
signal \N__35801\ : std_logic;
signal \N__35798\ : std_logic;
signal \N__35795\ : std_logic;
signal \N__35794\ : std_logic;
signal \N__35793\ : std_logic;
signal \N__35788\ : std_logic;
signal \N__35785\ : std_logic;
signal \N__35782\ : std_logic;
signal \N__35777\ : std_logic;
signal \N__35774\ : std_logic;
signal \N__35771\ : std_logic;
signal \N__35770\ : std_logic;
signal \N__35769\ : std_logic;
signal \N__35766\ : std_logic;
signal \N__35763\ : std_logic;
signal \N__35760\ : std_logic;
signal \N__35755\ : std_logic;
signal \N__35750\ : std_logic;
signal \N__35747\ : std_logic;
signal \N__35746\ : std_logic;
signal \N__35743\ : std_logic;
signal \N__35740\ : std_logic;
signal \N__35739\ : std_logic;
signal \N__35734\ : std_logic;
signal \N__35731\ : std_logic;
signal \N__35728\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35715\ : std_logic;
signal \N__35712\ : std_logic;
signal \N__35709\ : std_logic;
signal \N__35706\ : std_logic;
signal \N__35701\ : std_logic;
signal \N__35696\ : std_logic;
signal \N__35693\ : std_logic;
signal \N__35690\ : std_logic;
signal \N__35689\ : std_logic;
signal \N__35688\ : std_logic;
signal \N__35685\ : std_logic;
signal \N__35682\ : std_logic;
signal \N__35679\ : std_logic;
signal \N__35674\ : std_logic;
signal \N__35669\ : std_logic;
signal \N__35666\ : std_logic;
signal \N__35665\ : std_logic;
signal \N__35664\ : std_logic;
signal \N__35661\ : std_logic;
signal \N__35656\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35648\ : std_logic;
signal \N__35645\ : std_logic;
signal \N__35644\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35638\ : std_logic;
signal \N__35637\ : std_logic;
signal \N__35634\ : std_logic;
signal \N__35631\ : std_logic;
signal \N__35628\ : std_logic;
signal \N__35623\ : std_logic;
signal \N__35618\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35612\ : std_logic;
signal \N__35611\ : std_logic;
signal \N__35608\ : std_logic;
signal \N__35605\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35601\ : std_logic;
signal \N__35598\ : std_logic;
signal \N__35595\ : std_logic;
signal \N__35588\ : std_logic;
signal \N__35587\ : std_logic;
signal \N__35584\ : std_logic;
signal \N__35581\ : std_logic;
signal \N__35578\ : std_logic;
signal \N__35577\ : std_logic;
signal \N__35574\ : std_logic;
signal \N__35571\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35565\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35555\ : std_logic;
signal \N__35554\ : std_logic;
signal \N__35551\ : std_logic;
signal \N__35548\ : std_logic;
signal \N__35547\ : std_logic;
signal \N__35542\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35536\ : std_logic;
signal \N__35531\ : std_logic;
signal \N__35528\ : std_logic;
signal \N__35527\ : std_logic;
signal \N__35526\ : std_logic;
signal \N__35521\ : std_logic;
signal \N__35518\ : std_logic;
signal \N__35515\ : std_logic;
signal \N__35510\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35504\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35502\ : std_logic;
signal \N__35499\ : std_logic;
signal \N__35496\ : std_logic;
signal \N__35493\ : std_logic;
signal \N__35488\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35479\ : std_logic;
signal \N__35476\ : std_logic;
signal \N__35473\ : std_logic;
signal \N__35472\ : std_logic;
signal \N__35467\ : std_logic;
signal \N__35464\ : std_logic;
signal \N__35461\ : std_logic;
signal \N__35456\ : std_logic;
signal \N__35453\ : std_logic;
signal \N__35452\ : std_logic;
signal \N__35451\ : std_logic;
signal \N__35448\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35438\ : std_logic;
signal \N__35435\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35428\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35424\ : std_logic;
signal \N__35421\ : std_logic;
signal \N__35418\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35404\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35394\ : std_logic;
signal \N__35391\ : std_logic;
signal \N__35388\ : std_logic;
signal \N__35385\ : std_logic;
signal \N__35382\ : std_logic;
signal \N__35379\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35363\ : std_logic;
signal \N__35360\ : std_logic;
signal \N__35357\ : std_logic;
signal \N__35354\ : std_logic;
signal \N__35351\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35342\ : std_logic;
signal \N__35339\ : std_logic;
signal \N__35336\ : std_logic;
signal \N__35333\ : std_logic;
signal \N__35332\ : std_logic;
signal \N__35329\ : std_logic;
signal \N__35326\ : std_logic;
signal \N__35323\ : std_logic;
signal \N__35320\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35296\ : std_logic;
signal \N__35293\ : std_logic;
signal \N__35290\ : std_logic;
signal \N__35287\ : std_logic;
signal \N__35284\ : std_logic;
signal \N__35281\ : std_logic;
signal \N__35278\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35272\ : std_logic;
signal \N__35269\ : std_logic;
signal \N__35266\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35258\ : std_logic;
signal \N__35255\ : std_logic;
signal \N__35252\ : std_logic;
signal \N__35251\ : std_logic;
signal \N__35248\ : std_logic;
signal \N__35245\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35231\ : std_logic;
signal \N__35230\ : std_logic;
signal \N__35227\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35216\ : std_logic;
signal \N__35213\ : std_logic;
signal \N__35212\ : std_logic;
signal \N__35209\ : std_logic;
signal \N__35206\ : std_logic;
signal \N__35201\ : std_logic;
signal \N__35198\ : std_logic;
signal \N__35195\ : std_logic;
signal \N__35192\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35186\ : std_logic;
signal \N__35183\ : std_logic;
signal \N__35182\ : std_logic;
signal \N__35179\ : std_logic;
signal \N__35176\ : std_logic;
signal \N__35173\ : std_logic;
signal \N__35168\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35162\ : std_logic;
signal \N__35159\ : std_logic;
signal \N__35156\ : std_logic;
signal \N__35153\ : std_logic;
signal \N__35150\ : std_logic;
signal \N__35147\ : std_logic;
signal \N__35144\ : std_logic;
signal \N__35143\ : std_logic;
signal \N__35140\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35132\ : std_logic;
signal \N__35129\ : std_logic;
signal \N__35126\ : std_logic;
signal \N__35123\ : std_logic;
signal \N__35120\ : std_logic;
signal \N__35117\ : std_logic;
signal \N__35114\ : std_logic;
signal \N__35113\ : std_logic;
signal \N__35110\ : std_logic;
signal \N__35107\ : std_logic;
signal \N__35102\ : std_logic;
signal \N__35099\ : std_logic;
signal \N__35096\ : std_logic;
signal \N__35093\ : std_logic;
signal \N__35090\ : std_logic;
signal \N__35087\ : std_logic;
signal \N__35084\ : std_logic;
signal \N__35081\ : std_logic;
signal \N__35078\ : std_logic;
signal \N__35075\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35071\ : std_logic;
signal \N__35068\ : std_logic;
signal \N__35065\ : std_logic;
signal \N__35060\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35048\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35044\ : std_logic;
signal \N__35041\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35033\ : std_logic;
signal \N__35030\ : std_logic;
signal \N__35027\ : std_logic;
signal \N__35024\ : std_logic;
signal \N__35021\ : std_logic;
signal \N__35018\ : std_logic;
signal \N__35015\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35011\ : std_logic;
signal \N__35008\ : std_logic;
signal \N__35003\ : std_logic;
signal \N__35000\ : std_logic;
signal \N__34997\ : std_logic;
signal \N__34994\ : std_logic;
signal \N__34991\ : std_logic;
signal \N__34988\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34984\ : std_logic;
signal \N__34981\ : std_logic;
signal \N__34976\ : std_logic;
signal \N__34973\ : std_logic;
signal \N__34970\ : std_logic;
signal \N__34967\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34957\ : std_logic;
signal \N__34952\ : std_logic;
signal \N__34949\ : std_logic;
signal \N__34946\ : std_logic;
signal \N__34943\ : std_logic;
signal \N__34940\ : std_logic;
signal \N__34937\ : std_logic;
signal \N__34936\ : std_logic;
signal \N__34933\ : std_logic;
signal \N__34930\ : std_logic;
signal \N__34925\ : std_logic;
signal \N__34922\ : std_logic;
signal \N__34919\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34915\ : std_logic;
signal \N__34912\ : std_logic;
signal \N__34909\ : std_logic;
signal \N__34904\ : std_logic;
signal \N__34901\ : std_logic;
signal \N__34898\ : std_logic;
signal \N__34895\ : std_logic;
signal \N__34894\ : std_logic;
signal \N__34893\ : std_logic;
signal \N__34892\ : std_logic;
signal \N__34889\ : std_logic;
signal \N__34886\ : std_logic;
signal \N__34883\ : std_logic;
signal \N__34880\ : std_logic;
signal \N__34871\ : std_logic;
signal \N__34868\ : std_logic;
signal \N__34865\ : std_logic;
signal \N__34862\ : std_logic;
signal \N__34861\ : std_logic;
signal \N__34860\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34854\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34844\ : std_logic;
signal \N__34843\ : std_logic;
signal \N__34842\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34838\ : std_logic;
signal \N__34835\ : std_logic;
signal \N__34832\ : std_logic;
signal \N__34829\ : std_logic;
signal \N__34826\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34811\ : std_logic;
signal \N__34808\ : std_logic;
signal \N__34805\ : std_logic;
signal \N__34802\ : std_logic;
signal \N__34801\ : std_logic;
signal \N__34796\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34792\ : std_logic;
signal \N__34789\ : std_logic;
signal \N__34786\ : std_logic;
signal \N__34781\ : std_logic;
signal \N__34780\ : std_logic;
signal \N__34777\ : std_logic;
signal \N__34774\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34767\ : std_logic;
signal \N__34762\ : std_logic;
signal \N__34759\ : std_logic;
signal \N__34756\ : std_logic;
signal \N__34751\ : std_logic;
signal \N__34750\ : std_logic;
signal \N__34745\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34736\ : std_logic;
signal \N__34733\ : std_logic;
signal \N__34730\ : std_logic;
signal \N__34729\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34725\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34719\ : std_logic;
signal \N__34714\ : std_logic;
signal \N__34711\ : std_logic;
signal \N__34708\ : std_logic;
signal \N__34703\ : std_logic;
signal \N__34700\ : std_logic;
signal \N__34697\ : std_logic;
signal \N__34694\ : std_logic;
signal \N__34691\ : std_logic;
signal \N__34690\ : std_logic;
signal \N__34689\ : std_logic;
signal \N__34688\ : std_logic;
signal \N__34685\ : std_logic;
signal \N__34682\ : std_logic;
signal \N__34677\ : std_logic;
signal \N__34674\ : std_logic;
signal \N__34671\ : std_logic;
signal \N__34668\ : std_logic;
signal \N__34663\ : std_logic;
signal \N__34662\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34658\ : std_logic;
signal \N__34655\ : std_logic;
signal \N__34652\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34642\ : std_logic;
signal \N__34637\ : std_logic;
signal \N__34634\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34622\ : std_logic;
signal \N__34619\ : std_logic;
signal \N__34616\ : std_logic;
signal \N__34615\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34611\ : std_logic;
signal \N__34608\ : std_logic;
signal \N__34605\ : std_logic;
signal \N__34602\ : std_logic;
signal \N__34597\ : std_logic;
signal \N__34592\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34588\ : std_logic;
signal \N__34585\ : std_logic;
signal \N__34582\ : std_logic;
signal \N__34579\ : std_logic;
signal \N__34574\ : std_logic;
signal \N__34573\ : std_logic;
signal \N__34572\ : std_logic;
signal \N__34569\ : std_logic;
signal \N__34566\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34555\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34538\ : std_logic;
signal \N__34535\ : std_logic;
signal \N__34534\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34530\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34523\ : std_logic;
signal \N__34520\ : std_logic;
signal \N__34517\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34505\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34496\ : std_logic;
signal \N__34493\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34487\ : std_logic;
signal \N__34484\ : std_logic;
signal \N__34481\ : std_logic;
signal \N__34478\ : std_logic;
signal \N__34475\ : std_logic;
signal \N__34472\ : std_logic;
signal \N__34469\ : std_logic;
signal \N__34466\ : std_logic;
signal \N__34463\ : std_logic;
signal \N__34460\ : std_logic;
signal \N__34457\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34451\ : std_logic;
signal \N__34448\ : std_logic;
signal \N__34445\ : std_logic;
signal \N__34442\ : std_logic;
signal \N__34439\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34427\ : std_logic;
signal \N__34424\ : std_logic;
signal \N__34421\ : std_logic;
signal \N__34418\ : std_logic;
signal \N__34415\ : std_logic;
signal \N__34412\ : std_logic;
signal \N__34409\ : std_logic;
signal \N__34406\ : std_logic;
signal \N__34403\ : std_logic;
signal \N__34400\ : std_logic;
signal \N__34397\ : std_logic;
signal \N__34394\ : std_logic;
signal \N__34391\ : std_logic;
signal \N__34388\ : std_logic;
signal \N__34385\ : std_logic;
signal \N__34382\ : std_logic;
signal \N__34379\ : std_logic;
signal \N__34376\ : std_logic;
signal \N__34373\ : std_logic;
signal \N__34370\ : std_logic;
signal \N__34367\ : std_logic;
signal \N__34364\ : std_logic;
signal \N__34361\ : std_logic;
signal \N__34358\ : std_logic;
signal \N__34355\ : std_logic;
signal \N__34352\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34340\ : std_logic;
signal \N__34337\ : std_logic;
signal \N__34334\ : std_logic;
signal \N__34331\ : std_logic;
signal \N__34328\ : std_logic;
signal \N__34325\ : std_logic;
signal \N__34322\ : std_logic;
signal \N__34319\ : std_logic;
signal \N__34316\ : std_logic;
signal \N__34313\ : std_logic;
signal \N__34310\ : std_logic;
signal \N__34307\ : std_logic;
signal \N__34304\ : std_logic;
signal \N__34301\ : std_logic;
signal \N__34298\ : std_logic;
signal \N__34295\ : std_logic;
signal \N__34292\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34288\ : std_logic;
signal \N__34285\ : std_logic;
signal \N__34280\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34273\ : std_logic;
signal \N__34270\ : std_logic;
signal \N__34267\ : std_logic;
signal \N__34262\ : std_logic;
signal \N__34261\ : std_logic;
signal \N__34258\ : std_logic;
signal \N__34255\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34244\ : std_logic;
signal \N__34241\ : std_logic;
signal \N__34238\ : std_logic;
signal \N__34235\ : std_logic;
signal \N__34232\ : std_logic;
signal \N__34229\ : std_logic;
signal \N__34226\ : std_logic;
signal \N__34223\ : std_logic;
signal \N__34220\ : std_logic;
signal \N__34217\ : std_logic;
signal \N__34214\ : std_logic;
signal \N__34211\ : std_logic;
signal \N__34208\ : std_logic;
signal \N__34207\ : std_logic;
signal \N__34206\ : std_logic;
signal \N__34205\ : std_logic;
signal \N__34198\ : std_logic;
signal \N__34195\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34187\ : std_logic;
signal \N__34184\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34182\ : std_logic;
signal \N__34181\ : std_logic;
signal \N__34180\ : std_logic;
signal \N__34179\ : std_logic;
signal \N__34178\ : std_logic;
signal \N__34177\ : std_logic;
signal \N__34176\ : std_logic;
signal \N__34175\ : std_logic;
signal \N__34174\ : std_logic;
signal \N__34173\ : std_logic;
signal \N__34172\ : std_logic;
signal \N__34171\ : std_logic;
signal \N__34170\ : std_logic;
signal \N__34169\ : std_logic;
signal \N__34168\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34165\ : std_logic;
signal \N__34164\ : std_logic;
signal \N__34163\ : std_logic;
signal \N__34162\ : std_logic;
signal \N__34161\ : std_logic;
signal \N__34152\ : std_logic;
signal \N__34149\ : std_logic;
signal \N__34148\ : std_logic;
signal \N__34147\ : std_logic;
signal \N__34146\ : std_logic;
signal \N__34145\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34143\ : std_logic;
signal \N__34142\ : std_logic;
signal \N__34133\ : std_logic;
signal \N__34126\ : std_logic;
signal \N__34117\ : std_logic;
signal \N__34108\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34096\ : std_logic;
signal \N__34093\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34076\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34058\ : std_logic;
signal \N__34055\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34041\ : std_logic;
signal \N__34034\ : std_logic;
signal \N__34031\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34027\ : std_logic;
signal \N__34024\ : std_logic;
signal \N__34023\ : std_logic;
signal \N__34016\ : std_logic;
signal \N__34015\ : std_logic;
signal \N__34012\ : std_logic;
signal \N__34009\ : std_logic;
signal \N__34006\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__33998\ : std_logic;
signal \N__33997\ : std_logic;
signal \N__33994\ : std_logic;
signal \N__33991\ : std_logic;
signal \N__33986\ : std_logic;
signal \N__33983\ : std_logic;
signal \N__33980\ : std_logic;
signal \N__33979\ : std_logic;
signal \N__33978\ : std_logic;
signal \N__33973\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33967\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33959\ : std_logic;
signal \N__33956\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33954\ : std_logic;
signal \N__33949\ : std_logic;
signal \N__33946\ : std_logic;
signal \N__33943\ : std_logic;
signal \N__33938\ : std_logic;
signal \N__33935\ : std_logic;
signal \N__33932\ : std_logic;
signal \N__33929\ : std_logic;
signal \N__33926\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33920\ : std_logic;
signal \N__33917\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33908\ : std_logic;
signal \N__33905\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33896\ : std_logic;
signal \N__33893\ : std_logic;
signal \N__33890\ : std_logic;
signal \N__33889\ : std_logic;
signal \N__33884\ : std_logic;
signal \N__33881\ : std_logic;
signal \N__33878\ : std_logic;
signal \N__33875\ : std_logic;
signal \N__33872\ : std_logic;
signal \N__33869\ : std_logic;
signal \N__33866\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33857\ : std_logic;
signal \N__33854\ : std_logic;
signal \N__33851\ : std_logic;
signal \N__33848\ : std_logic;
signal \N__33847\ : std_logic;
signal \N__33842\ : std_logic;
signal \N__33839\ : std_logic;
signal \N__33836\ : std_logic;
signal \N__33833\ : std_logic;
signal \N__33830\ : std_logic;
signal \N__33827\ : std_logic;
signal \N__33824\ : std_logic;
signal \N__33821\ : std_logic;
signal \N__33818\ : std_logic;
signal \N__33815\ : std_logic;
signal \N__33812\ : std_logic;
signal \N__33809\ : std_logic;
signal \N__33806\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33800\ : std_logic;
signal \N__33797\ : std_logic;
signal \N__33794\ : std_logic;
signal \N__33791\ : std_logic;
signal \N__33788\ : std_logic;
signal \N__33787\ : std_logic;
signal \N__33784\ : std_logic;
signal \N__33781\ : std_logic;
signal \N__33778\ : std_logic;
signal \N__33775\ : std_logic;
signal \N__33772\ : std_logic;
signal \N__33769\ : std_logic;
signal \N__33764\ : std_logic;
signal \N__33763\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33757\ : std_logic;
signal \N__33754\ : std_logic;
signal \N__33751\ : std_logic;
signal \N__33748\ : std_logic;
signal \N__33745\ : std_logic;
signal \N__33742\ : std_logic;
signal \N__33741\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33735\ : std_logic;
signal \N__33732\ : std_logic;
signal \N__33729\ : std_logic;
signal \N__33722\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33708\ : std_logic;
signal \N__33705\ : std_logic;
signal \N__33702\ : std_logic;
signal \N__33699\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33677\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33665\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33653\ : std_logic;
signal \N__33650\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33638\ : std_logic;
signal \N__33635\ : std_logic;
signal \N__33632\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33623\ : std_logic;
signal \N__33620\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33614\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33599\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33593\ : std_logic;
signal \N__33590\ : std_logic;
signal \N__33587\ : std_logic;
signal \N__33584\ : std_logic;
signal \N__33581\ : std_logic;
signal \N__33578\ : std_logic;
signal \N__33575\ : std_logic;
signal \N__33572\ : std_logic;
signal \N__33569\ : std_logic;
signal \N__33566\ : std_logic;
signal \N__33563\ : std_logic;
signal \N__33560\ : std_logic;
signal \N__33557\ : std_logic;
signal \N__33554\ : std_logic;
signal \N__33551\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33545\ : std_logic;
signal \N__33542\ : std_logic;
signal \N__33539\ : std_logic;
signal \N__33536\ : std_logic;
signal \N__33533\ : std_logic;
signal \N__33530\ : std_logic;
signal \N__33527\ : std_logic;
signal \N__33524\ : std_logic;
signal \N__33521\ : std_logic;
signal \N__33518\ : std_logic;
signal \N__33515\ : std_logic;
signal \N__33512\ : std_logic;
signal \N__33509\ : std_logic;
signal \N__33506\ : std_logic;
signal \N__33503\ : std_logic;
signal \N__33500\ : std_logic;
signal \N__33497\ : std_logic;
signal \N__33494\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33488\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33482\ : std_logic;
signal \N__33479\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33473\ : std_logic;
signal \N__33470\ : std_logic;
signal \N__33467\ : std_logic;
signal \N__33464\ : std_logic;
signal \N__33463\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33454\ : std_logic;
signal \N__33449\ : std_logic;
signal \N__33446\ : std_logic;
signal \N__33445\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33443\ : std_logic;
signal \N__33440\ : std_logic;
signal \N__33437\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33422\ : std_logic;
signal \N__33421\ : std_logic;
signal \N__33420\ : std_logic;
signal \N__33419\ : std_logic;
signal \N__33418\ : std_logic;
signal \N__33417\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33415\ : std_logic;
signal \N__33414\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33412\ : std_logic;
signal \N__33411\ : std_logic;
signal \N__33410\ : std_logic;
signal \N__33409\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33407\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33405\ : std_logic;
signal \N__33404\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33402\ : std_logic;
signal \N__33401\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33399\ : std_logic;
signal \N__33398\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33396\ : std_logic;
signal \N__33395\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33393\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33375\ : std_logic;
signal \N__33370\ : std_logic;
signal \N__33361\ : std_logic;
signal \N__33352\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33334\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33314\ : std_logic;
signal \N__33305\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33284\ : std_logic;
signal \N__33281\ : std_logic;
signal \N__33278\ : std_logic;
signal \N__33275\ : std_logic;
signal \N__33272\ : std_logic;
signal \N__33269\ : std_logic;
signal \N__33266\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33257\ : std_logic;
signal \N__33254\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33248\ : std_logic;
signal \N__33245\ : std_logic;
signal \N__33244\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33237\ : std_logic;
signal \N__33236\ : std_logic;
signal \N__33233\ : std_logic;
signal \N__33230\ : std_logic;
signal \N__33227\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33217\ : std_logic;
signal \N__33214\ : std_logic;
signal \N__33211\ : std_logic;
signal \N__33208\ : std_logic;
signal \N__33203\ : std_logic;
signal \N__33200\ : std_logic;
signal \N__33199\ : std_logic;
signal \N__33196\ : std_logic;
signal \N__33195\ : std_logic;
signal \N__33194\ : std_logic;
signal \N__33191\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33179\ : std_logic;
signal \N__33176\ : std_logic;
signal \N__33173\ : std_logic;
signal \N__33170\ : std_logic;
signal \N__33167\ : std_logic;
signal \N__33164\ : std_logic;
signal \N__33161\ : std_logic;
signal \N__33158\ : std_logic;
signal \N__33155\ : std_logic;
signal \N__33152\ : std_logic;
signal \N__33149\ : std_logic;
signal \N__33146\ : std_logic;
signal \N__33143\ : std_logic;
signal \N__33140\ : std_logic;
signal \N__33137\ : std_logic;
signal \N__33134\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33128\ : std_logic;
signal \N__33125\ : std_logic;
signal \N__33122\ : std_logic;
signal \N__33119\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33114\ : std_logic;
signal \N__33107\ : std_logic;
signal \N__33104\ : std_logic;
signal \N__33101\ : std_logic;
signal \N__33098\ : std_logic;
signal \N__33095\ : std_logic;
signal \N__33092\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33086\ : std_logic;
signal \N__33083\ : std_logic;
signal \N__33080\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33077\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33073\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33057\ : std_logic;
signal \N__33050\ : std_logic;
signal \N__33049\ : std_logic;
signal \N__33046\ : std_logic;
signal \N__33043\ : std_logic;
signal \N__33038\ : std_logic;
signal \N__33035\ : std_logic;
signal \N__33032\ : std_logic;
signal \N__33029\ : std_logic;
signal \N__33026\ : std_logic;
signal \N__33025\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33017\ : std_logic;
signal \N__33014\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33010\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33004\ : std_logic;
signal \N__33003\ : std_logic;
signal \N__33002\ : std_logic;
signal \N__32999\ : std_logic;
signal \N__32996\ : std_logic;
signal \N__32991\ : std_logic;
signal \N__32988\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32978\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32972\ : std_logic;
signal \N__32969\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32963\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32959\ : std_logic;
signal \N__32956\ : std_logic;
signal \N__32953\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32947\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32940\ : std_logic;
signal \N__32937\ : std_logic;
signal \N__32934\ : std_logic;
signal \N__32927\ : std_logic;
signal \N__32926\ : std_logic;
signal \N__32921\ : std_logic;
signal \N__32918\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32906\ : std_logic;
signal \N__32903\ : std_logic;
signal \N__32902\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32890\ : std_logic;
signal \N__32887\ : std_logic;
signal \N__32884\ : std_logic;
signal \N__32879\ : std_logic;
signal \N__32878\ : std_logic;
signal \N__32875\ : std_logic;
signal \N__32872\ : std_logic;
signal \N__32871\ : std_logic;
signal \N__32870\ : std_logic;
signal \N__32867\ : std_logic;
signal \N__32864\ : std_logic;
signal \N__32859\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32851\ : std_logic;
signal \N__32848\ : std_logic;
signal \N__32847\ : std_logic;
signal \N__32844\ : std_logic;
signal \N__32841\ : std_logic;
signal \N__32838\ : std_logic;
signal \N__32831\ : std_logic;
signal \N__32830\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32821\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32813\ : std_logic;
signal \N__32812\ : std_logic;
signal \N__32811\ : std_logic;
signal \N__32808\ : std_logic;
signal \N__32803\ : std_logic;
signal \N__32802\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32783\ : std_logic;
signal \N__32780\ : std_logic;
signal \N__32777\ : std_logic;
signal \N__32774\ : std_logic;
signal \N__32771\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32759\ : std_logic;
signal \N__32756\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32732\ : std_logic;
signal \N__32729\ : std_logic;
signal \N__32726\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32720\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32714\ : std_logic;
signal \N__32711\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32699\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32693\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32671\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32668\ : std_logic;
signal \N__32667\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32665\ : std_logic;
signal \N__32664\ : std_logic;
signal \N__32663\ : std_logic;
signal \N__32662\ : std_logic;
signal \N__32661\ : std_logic;
signal \N__32660\ : std_logic;
signal \N__32659\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32657\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32655\ : std_logic;
signal \N__32654\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32648\ : std_logic;
signal \N__32647\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32626\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32616\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32612\ : std_logic;
signal \N__32611\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32608\ : std_logic;
signal \N__32607\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32605\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32601\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32598\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32594\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32584\ : std_logic;
signal \N__32581\ : std_logic;
signal \N__32578\ : std_logic;
signal \N__32575\ : std_logic;
signal \N__32574\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32572\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32568\ : std_logic;
signal \N__32559\ : std_logic;
signal \N__32556\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32554\ : std_logic;
signal \N__32553\ : std_logic;
signal \N__32552\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32540\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32528\ : std_logic;
signal \N__32525\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32512\ : std_logic;
signal \N__32509\ : std_logic;
signal \N__32506\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32498\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32492\ : std_logic;
signal \N__32489\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32475\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32453\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32443\ : std_logic;
signal \N__32438\ : std_logic;
signal \N__32435\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32419\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32409\ : std_logic;
signal \N__32406\ : std_logic;
signal \N__32399\ : std_logic;
signal \N__32396\ : std_logic;
signal \N__32395\ : std_logic;
signal \N__32392\ : std_logic;
signal \N__32389\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32378\ : std_logic;
signal \N__32377\ : std_logic;
signal \N__32374\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32372\ : std_logic;
signal \N__32369\ : std_logic;
signal \N__32368\ : std_logic;
signal \N__32365\ : std_logic;
signal \N__32360\ : std_logic;
signal \N__32357\ : std_logic;
signal \N__32354\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32342\ : std_logic;
signal \N__32339\ : std_logic;
signal \N__32336\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32329\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32323\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32312\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32308\ : std_logic;
signal \N__32305\ : std_logic;
signal \N__32302\ : std_logic;
signal \N__32297\ : std_logic;
signal \N__32296\ : std_logic;
signal \N__32295\ : std_logic;
signal \N__32294\ : std_logic;
signal \N__32287\ : std_logic;
signal \N__32286\ : std_logic;
signal \N__32283\ : std_logic;
signal \N__32280\ : std_logic;
signal \N__32275\ : std_logic;
signal \N__32272\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32266\ : std_logic;
signal \N__32263\ : std_logic;
signal \N__32262\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32258\ : std_logic;
signal \N__32255\ : std_logic;
signal \N__32252\ : std_logic;
signal \N__32249\ : std_logic;
signal \N__32242\ : std_logic;
signal \N__32239\ : std_logic;
signal \N__32236\ : std_logic;
signal \N__32231\ : std_logic;
signal \N__32230\ : std_logic;
signal \N__32229\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32221\ : std_logic;
signal \N__32216\ : std_logic;
signal \N__32213\ : std_logic;
signal \N__32210\ : std_logic;
signal \N__32207\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32195\ : std_logic;
signal \N__32192\ : std_logic;
signal \N__32191\ : std_logic;
signal \N__32190\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32188\ : std_logic;
signal \N__32187\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32185\ : std_logic;
signal \N__32184\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32182\ : std_logic;
signal \N__32181\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32179\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32176\ : std_logic;
signal \N__32175\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32173\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32167\ : std_logic;
signal \N__32166\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32156\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32140\ : std_logic;
signal \N__32131\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32119\ : std_logic;
signal \N__32116\ : std_logic;
signal \N__32115\ : std_logic;
signal \N__32114\ : std_logic;
signal \N__32113\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32111\ : std_logic;
signal \N__32110\ : std_logic;
signal \N__32109\ : std_logic;
signal \N__32100\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32083\ : std_logic;
signal \N__32076\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32064\ : std_logic;
signal \N__32059\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32045\ : std_logic;
signal \N__32042\ : std_logic;
signal \N__32041\ : std_logic;
signal \N__32040\ : std_logic;
signal \N__32039\ : std_logic;
signal \N__32036\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32022\ : std_logic;
signal \N__32017\ : std_logic;
signal \N__32012\ : std_logic;
signal \N__32009\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32006\ : std_logic;
signal \N__32005\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32003\ : std_logic;
signal \N__32000\ : std_logic;
signal \N__31997\ : std_logic;
signal \N__31996\ : std_logic;
signal \N__31995\ : std_logic;
signal \N__31994\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31991\ : std_logic;
signal \N__31990\ : std_logic;
signal \N__31989\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31987\ : std_logic;
signal \N__31986\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31984\ : std_logic;
signal \N__31983\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31981\ : std_logic;
signal \N__31980\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31978\ : std_logic;
signal \N__31977\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31975\ : std_logic;
signal \N__31974\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31972\ : std_logic;
signal \N__31971\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31969\ : std_logic;
signal \N__31968\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31966\ : std_logic;
signal \N__31965\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31959\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31947\ : std_logic;
signal \N__31944\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31942\ : std_logic;
signal \N__31941\ : std_logic;
signal \N__31940\ : std_logic;
signal \N__31939\ : std_logic;
signal \N__31938\ : std_logic;
signal \N__31937\ : std_logic;
signal \N__31932\ : std_logic;
signal \N__31925\ : std_logic;
signal \N__31922\ : std_logic;
signal \N__31913\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31910\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31907\ : std_logic;
signal \N__31906\ : std_logic;
signal \N__31905\ : std_logic;
signal \N__31904\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31902\ : std_logic;
signal \N__31901\ : std_logic;
signal \N__31900\ : std_logic;
signal \N__31899\ : std_logic;
signal \N__31898\ : std_logic;
signal \N__31895\ : std_logic;
signal \N__31894\ : std_logic;
signal \N__31885\ : std_logic;
signal \N__31882\ : std_logic;
signal \N__31865\ : std_logic;
signal \N__31854\ : std_logic;
signal \N__31849\ : std_logic;
signal \N__31838\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31834\ : std_logic;
signal \N__31833\ : std_logic;
signal \N__31830\ : std_logic;
signal \N__31823\ : std_logic;
signal \N__31816\ : std_logic;
signal \N__31815\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31813\ : std_logic;
signal \N__31812\ : std_logic;
signal \N__31809\ : std_logic;
signal \N__31806\ : std_logic;
signal \N__31801\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31793\ : std_logic;
signal \N__31790\ : std_logic;
signal \N__31781\ : std_logic;
signal \N__31780\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31778\ : std_logic;
signal \N__31777\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31775\ : std_logic;
signal \N__31774\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31771\ : std_logic;
signal \N__31770\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31766\ : std_logic;
signal \N__31765\ : std_logic;
signal \N__31764\ : std_logic;
signal \N__31761\ : std_logic;
signal \N__31750\ : std_logic;
signal \N__31749\ : std_logic;
signal \N__31748\ : std_logic;
signal \N__31747\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31706\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31693\ : std_logic;
signal \N__31684\ : std_logic;
signal \N__31679\ : std_logic;
signal \N__31674\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31668\ : std_logic;
signal \N__31665\ : std_logic;
signal \N__31656\ : std_logic;
signal \N__31645\ : std_logic;
signal \N__31638\ : std_logic;
signal \N__31635\ : std_logic;
signal \N__31630\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31616\ : std_logic;
signal \N__31603\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31565\ : std_logic;
signal \N__31562\ : std_logic;
signal \N__31561\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31557\ : std_logic;
signal \N__31554\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31532\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31526\ : std_logic;
signal \N__31523\ : std_logic;
signal \N__31520\ : std_logic;
signal \N__31517\ : std_logic;
signal \N__31514\ : std_logic;
signal \N__31511\ : std_logic;
signal \N__31510\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31498\ : std_logic;
signal \N__31493\ : std_logic;
signal \N__31492\ : std_logic;
signal \N__31491\ : std_logic;
signal \N__31488\ : std_logic;
signal \N__31485\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31475\ : std_logic;
signal \N__31472\ : std_logic;
signal \N__31469\ : std_logic;
signal \N__31466\ : std_logic;
signal \N__31463\ : std_logic;
signal \N__31462\ : std_logic;
signal \N__31457\ : std_logic;
signal \N__31454\ : std_logic;
signal \N__31453\ : std_logic;
signal \N__31450\ : std_logic;
signal \N__31447\ : std_logic;
signal \N__31446\ : std_logic;
signal \N__31443\ : std_logic;
signal \N__31440\ : std_logic;
signal \N__31437\ : std_logic;
signal \N__31434\ : std_logic;
signal \N__31431\ : std_logic;
signal \N__31424\ : std_logic;
signal \N__31421\ : std_logic;
signal \N__31420\ : std_logic;
signal \N__31417\ : std_logic;
signal \N__31414\ : std_logic;
signal \N__31413\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31409\ : std_logic;
signal \N__31406\ : std_logic;
signal \N__31403\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31387\ : std_logic;
signal \N__31382\ : std_logic;
signal \N__31381\ : std_logic;
signal \N__31376\ : std_logic;
signal \N__31373\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31371\ : std_logic;
signal \N__31368\ : std_logic;
signal \N__31363\ : std_logic;
signal \N__31362\ : std_logic;
signal \N__31359\ : std_logic;
signal \N__31356\ : std_logic;
signal \N__31353\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31340\ : std_logic;
signal \N__31339\ : std_logic;
signal \N__31336\ : std_logic;
signal \N__31333\ : std_logic;
signal \N__31328\ : std_logic;
signal \N__31325\ : std_logic;
signal \N__31322\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31316\ : std_logic;
signal \N__31315\ : std_logic;
signal \N__31314\ : std_logic;
signal \N__31313\ : std_logic;
signal \N__31312\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31309\ : std_logic;
signal \N__31308\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31283\ : std_logic;
signal \N__31280\ : std_logic;
signal \N__31277\ : std_logic;
signal \N__31276\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31274\ : std_logic;
signal \N__31271\ : std_logic;
signal \N__31266\ : std_logic;
signal \N__31263\ : std_logic;
signal \N__31258\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31247\ : std_logic;
signal \N__31244\ : std_logic;
signal \N__31241\ : std_logic;
signal \N__31238\ : std_logic;
signal \N__31237\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31228\ : std_logic;
signal \N__31225\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31219\ : std_logic;
signal \N__31216\ : std_logic;
signal \N__31213\ : std_logic;
signal \N__31208\ : std_logic;
signal \N__31205\ : std_logic;
signal \N__31204\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31197\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31187\ : std_logic;
signal \N__31184\ : std_logic;
signal \N__31181\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31175\ : std_logic;
signal \N__31174\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31170\ : std_logic;
signal \N__31169\ : std_logic;
signal \N__31166\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31151\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31138\ : std_logic;
signal \N__31133\ : std_logic;
signal \N__31132\ : std_logic;
signal \N__31129\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31122\ : std_logic;
signal \N__31121\ : std_logic;
signal \N__31118\ : std_logic;
signal \N__31113\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31100\ : std_logic;
signal \N__31097\ : std_logic;
signal \N__31096\ : std_logic;
signal \N__31093\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31086\ : std_logic;
signal \N__31083\ : std_logic;
signal \N__31080\ : std_logic;
signal \N__31077\ : std_logic;
signal \N__31074\ : std_logic;
signal \N__31071\ : std_logic;
signal \N__31064\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31058\ : std_logic;
signal \N__31055\ : std_logic;
signal \N__31052\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31040\ : std_logic;
signal \N__31039\ : std_logic;
signal \N__31036\ : std_logic;
signal \N__31033\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31025\ : std_logic;
signal \N__31024\ : std_logic;
signal \N__31023\ : std_logic;
signal \N__31018\ : std_logic;
signal \N__31015\ : std_logic;
signal \N__31012\ : std_logic;
signal \N__31011\ : std_logic;
signal \N__31006\ : std_logic;
signal \N__31003\ : std_logic;
signal \N__31000\ : std_logic;
signal \N__30997\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30991\ : std_logic;
signal \N__30986\ : std_logic;
signal \N__30983\ : std_logic;
signal \N__30982\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30976\ : std_logic;
signal \N__30973\ : std_logic;
signal \N__30970\ : std_logic;
signal \N__30965\ : std_logic;
signal \N__30964\ : std_logic;
signal \N__30961\ : std_logic;
signal \N__30958\ : std_logic;
signal \N__30957\ : std_logic;
signal \N__30952\ : std_logic;
signal \N__30949\ : std_logic;
signal \N__30946\ : std_logic;
signal \N__30941\ : std_logic;
signal \N__30940\ : std_logic;
signal \N__30935\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30926\ : std_logic;
signal \N__30923\ : std_logic;
signal \N__30920\ : std_logic;
signal \N__30919\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30912\ : std_logic;
signal \N__30909\ : std_logic;
signal \N__30906\ : std_logic;
signal \N__30903\ : std_logic;
signal \N__30900\ : std_logic;
signal \N__30895\ : std_logic;
signal \N__30890\ : std_logic;
signal \N__30887\ : std_logic;
signal \N__30884\ : std_logic;
signal \N__30881\ : std_logic;
signal \N__30878\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30872\ : std_logic;
signal \N__30869\ : std_logic;
signal \N__30866\ : std_logic;
signal \N__30863\ : std_logic;
signal \N__30862\ : std_logic;
signal \N__30861\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30848\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30842\ : std_logic;
signal \N__30839\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30827\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30821\ : std_logic;
signal \N__30818\ : std_logic;
signal \N__30815\ : std_logic;
signal \N__30812\ : std_logic;
signal \N__30811\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30807\ : std_logic;
signal \N__30804\ : std_logic;
signal \N__30801\ : std_logic;
signal \N__30798\ : std_logic;
signal \N__30793\ : std_logic;
signal \N__30790\ : std_logic;
signal \N__30787\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30776\ : std_logic;
signal \N__30775\ : std_logic;
signal \N__30772\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30767\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30749\ : std_logic;
signal \N__30746\ : std_logic;
signal \N__30745\ : std_logic;
signal \N__30744\ : std_logic;
signal \N__30741\ : std_logic;
signal \N__30738\ : std_logic;
signal \N__30735\ : std_logic;
signal \N__30730\ : std_logic;
signal \N__30725\ : std_logic;
signal \N__30724\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30720\ : std_logic;
signal \N__30719\ : std_logic;
signal \N__30716\ : std_logic;
signal \N__30713\ : std_logic;
signal \N__30710\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30702\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30694\ : std_logic;
signal \N__30693\ : std_logic;
signal \N__30690\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30680\ : std_logic;
signal \N__30677\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30663\ : std_logic;
signal \N__30660\ : std_logic;
signal \N__30657\ : std_logic;
signal \N__30654\ : std_logic;
signal \N__30651\ : std_logic;
signal \N__30644\ : std_logic;
signal \N__30643\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30630\ : std_logic;
signal \N__30623\ : std_logic;
signal \N__30622\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30618\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30609\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30596\ : std_logic;
signal \N__30595\ : std_logic;
signal \N__30592\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30588\ : std_logic;
signal \N__30585\ : std_logic;
signal \N__30582\ : std_logic;
signal \N__30575\ : std_logic;
signal \N__30572\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30567\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30561\ : std_logic;
signal \N__30554\ : std_logic;
signal \N__30551\ : std_logic;
signal \N__30550\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30548\ : std_logic;
signal \N__30541\ : std_logic;
signal \N__30538\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30530\ : std_logic;
signal \N__30527\ : std_logic;
signal \N__30524\ : std_logic;
signal \N__30521\ : std_logic;
signal \N__30520\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30518\ : std_logic;
signal \N__30515\ : std_logic;
signal \N__30510\ : std_logic;
signal \N__30507\ : std_logic;
signal \N__30502\ : std_logic;
signal \N__30497\ : std_logic;
signal \N__30494\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30490\ : std_logic;
signal \N__30487\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30479\ : std_logic;
signal \N__30476\ : std_logic;
signal \N__30473\ : std_logic;
signal \N__30470\ : std_logic;
signal \N__30467\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30465\ : std_logic;
signal \N__30464\ : std_logic;
signal \N__30461\ : std_logic;
signal \N__30458\ : std_logic;
signal \N__30455\ : std_logic;
signal \N__30452\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30440\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30419\ : std_logic;
signal \N__30416\ : std_logic;
signal \N__30415\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30409\ : std_logic;
signal \N__30406\ : std_logic;
signal \N__30403\ : std_logic;
signal \N__30400\ : std_logic;
signal \N__30395\ : std_logic;
signal \N__30392\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30383\ : std_logic;
signal \N__30382\ : std_logic;
signal \N__30377\ : std_logic;
signal \N__30376\ : std_logic;
signal \N__30373\ : std_logic;
signal \N__30370\ : std_logic;
signal \N__30367\ : std_logic;
signal \N__30362\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30353\ : std_logic;
signal \N__30352\ : std_logic;
signal \N__30349\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30343\ : std_logic;
signal \N__30338\ : std_logic;
signal \N__30335\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30333\ : std_logic;
signal \N__30330\ : std_logic;
signal \N__30325\ : std_logic;
signal \N__30320\ : std_logic;
signal \N__30317\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30315\ : std_logic;
signal \N__30312\ : std_logic;
signal \N__30309\ : std_logic;
signal \N__30304\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30294\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30274\ : std_logic;
signal \N__30271\ : std_logic;
signal \N__30270\ : std_logic;
signal \N__30267\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30258\ : std_logic;
signal \N__30255\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30245\ : std_logic;
signal \N__30244\ : std_logic;
signal \N__30241\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30230\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30226\ : std_logic;
signal \N__30223\ : std_logic;
signal \N__30218\ : std_logic;
signal \N__30215\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30208\ : std_logic;
signal \N__30203\ : std_logic;
signal \N__30200\ : std_logic;
signal \N__30199\ : std_logic;
signal \N__30196\ : std_logic;
signal \N__30193\ : std_logic;
signal \N__30188\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30184\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30178\ : std_logic;
signal \N__30173\ : std_logic;
signal \N__30170\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30166\ : std_logic;
signal \N__30161\ : std_logic;
signal \N__30160\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30151\ : std_logic;
signal \N__30146\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30139\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30135\ : std_logic;
signal \N__30132\ : std_logic;
signal \N__30129\ : std_logic;
signal \N__30124\ : std_logic;
signal \N__30119\ : std_logic;
signal \N__30116\ : std_logic;
signal \N__30115\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30103\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30095\ : std_logic;
signal \N__30092\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30086\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30082\ : std_logic;
signal \N__30079\ : std_logic;
signal \N__30076\ : std_logic;
signal \N__30071\ : std_logic;
signal \N__30068\ : std_logic;
signal \N__30067\ : std_logic;
signal \N__30064\ : std_logic;
signal \N__30061\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30053\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30046\ : std_logic;
signal \N__30041\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30037\ : std_logic;
signal \N__30034\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30023\ : std_logic;
signal \N__30022\ : std_logic;
signal \N__30019\ : std_logic;
signal \N__30016\ : std_logic;
signal \N__30011\ : std_logic;
signal \N__30008\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30004\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__29996\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29986\ : std_logic;
signal \N__29983\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29974\ : std_logic;
signal \N__29971\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29963\ : std_logic;
signal \N__29960\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29954\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29935\ : std_logic;
signal \N__29932\ : std_logic;
signal \N__29929\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29920\ : std_logic;
signal \N__29919\ : std_logic;
signal \N__29916\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29908\ : std_logic;
signal \N__29905\ : std_logic;
signal \N__29902\ : std_logic;
signal \N__29899\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29893\ : std_logic;
signal \N__29890\ : std_logic;
signal \N__29889\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29867\ : std_logic;
signal \N__29864\ : std_logic;
signal \N__29861\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29845\ : std_logic;
signal \N__29842\ : std_logic;
signal \N__29839\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29829\ : std_logic;
signal \N__29822\ : std_logic;
signal \N__29821\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29810\ : std_logic;
signal \N__29807\ : std_logic;
signal \N__29806\ : std_logic;
signal \N__29805\ : std_logic;
signal \N__29802\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29786\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29779\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29776\ : std_logic;
signal \N__29775\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29773\ : std_logic;
signal \N__29772\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29766\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29748\ : std_logic;
signal \N__29745\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29734\ : std_logic;
signal \N__29731\ : std_logic;
signal \N__29730\ : std_logic;
signal \N__29727\ : std_logic;
signal \N__29724\ : std_logic;
signal \N__29721\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29713\ : std_logic;
signal \N__29710\ : std_logic;
signal \N__29707\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29703\ : std_logic;
signal \N__29700\ : std_logic;
signal \N__29697\ : std_logic;
signal \N__29696\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29685\ : std_logic;
signal \N__29682\ : std_logic;
signal \N__29679\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29669\ : std_logic;
signal \N__29666\ : std_logic;
signal \N__29663\ : std_logic;
signal \N__29660\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29654\ : std_logic;
signal \N__29653\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29645\ : std_logic;
signal \N__29644\ : std_logic;
signal \N__29641\ : std_logic;
signal \N__29638\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29627\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29621\ : std_logic;
signal \N__29620\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29611\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29605\ : std_logic;
signal \N__29604\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29595\ : std_logic;
signal \N__29588\ : std_logic;
signal \N__29585\ : std_logic;
signal \N__29584\ : std_logic;
signal \N__29581\ : std_logic;
signal \N__29578\ : std_logic;
signal \N__29573\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29567\ : std_logic;
signal \N__29564\ : std_logic;
signal \N__29561\ : std_logic;
signal \N__29558\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29540\ : std_logic;
signal \N__29537\ : std_logic;
signal \N__29536\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29526\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29515\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29498\ : std_logic;
signal \N__29495\ : std_logic;
signal \N__29494\ : std_logic;
signal \N__29493\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29487\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29477\ : std_logic;
signal \N__29474\ : std_logic;
signal \N__29473\ : std_logic;
signal \N__29472\ : std_logic;
signal \N__29469\ : std_logic;
signal \N__29466\ : std_logic;
signal \N__29463\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29452\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29435\ : std_logic;
signal \N__29432\ : std_logic;
signal \N__29429\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29421\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29408\ : std_logic;
signal \N__29407\ : std_logic;
signal \N__29404\ : std_logic;
signal \N__29401\ : std_logic;
signal \N__29400\ : std_logic;
signal \N__29397\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29379\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29366\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29360\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29350\ : std_logic;
signal \N__29349\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29342\ : std_logic;
signal \N__29339\ : std_logic;
signal \N__29336\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29321\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29312\ : std_logic;
signal \N__29309\ : std_logic;
signal \N__29306\ : std_logic;
signal \N__29303\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29296\ : std_logic;
signal \N__29293\ : std_logic;
signal \N__29290\ : std_logic;
signal \N__29287\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29276\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29255\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29252\ : std_logic;
signal \N__29251\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29249\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29237\ : std_logic;
signal \N__29236\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29234\ : std_logic;
signal \N__29233\ : std_logic;
signal \N__29232\ : std_logic;
signal \N__29231\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29229\ : std_logic;
signal \N__29228\ : std_logic;
signal \N__29227\ : std_logic;
signal \N__29226\ : std_logic;
signal \N__29225\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29222\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29219\ : std_logic;
signal \N__29218\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29205\ : std_logic;
signal \N__29196\ : std_logic;
signal \N__29191\ : std_logic;
signal \N__29182\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29164\ : std_logic;
signal \N__29155\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29132\ : std_logic;
signal \N__29129\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29119\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29112\ : std_logic;
signal \N__29109\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29099\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29095\ : std_logic;
signal \N__29094\ : std_logic;
signal \N__29091\ : std_logic;
signal \N__29088\ : std_logic;
signal \N__29085\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29075\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29055\ : std_logic;
signal \N__29052\ : std_logic;
signal \N__29049\ : std_logic;
signal \N__29046\ : std_logic;
signal \N__29039\ : std_logic;
signal \N__29036\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29032\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29026\ : std_logic;
signal \N__29025\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29017\ : std_logic;
signal \N__29014\ : std_logic;
signal \N__29009\ : std_logic;
signal \N__29008\ : std_logic;
signal \N__29007\ : std_logic;
signal \N__29004\ : std_logic;
signal \N__29001\ : std_logic;
signal \N__28998\ : std_logic;
signal \N__28995\ : std_logic;
signal \N__28992\ : std_logic;
signal \N__28989\ : std_logic;
signal \N__28984\ : std_logic;
signal \N__28983\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28970\ : std_logic;
signal \N__28967\ : std_logic;
signal \N__28964\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28940\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28923\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28914\ : std_logic;
signal \N__28911\ : std_logic;
signal \N__28904\ : std_logic;
signal \N__28903\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28901\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28890\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28882\ : std_logic;
signal \N__28879\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28871\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28864\ : std_logic;
signal \N__28863\ : std_logic;
signal \N__28860\ : std_logic;
signal \N__28857\ : std_logic;
signal \N__28854\ : std_logic;
signal \N__28851\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28840\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28823\ : std_logic;
signal \N__28820\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28813\ : std_logic;
signal \N__28810\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28799\ : std_logic;
signal \N__28798\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28782\ : std_logic;
signal \N__28779\ : std_logic;
signal \N__28776\ : std_logic;
signal \N__28773\ : std_logic;
signal \N__28768\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28760\ : std_logic;
signal \N__28759\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28755\ : std_logic;
signal \N__28752\ : std_logic;
signal \N__28749\ : std_logic;
signal \N__28746\ : std_logic;
signal \N__28743\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28739\ : std_logic;
signal \N__28732\ : std_logic;
signal \N__28729\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28718\ : std_logic;
signal \N__28717\ : std_logic;
signal \N__28714\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28710\ : std_logic;
signal \N__28709\ : std_logic;
signal \N__28706\ : std_logic;
signal \N__28703\ : std_logic;
signal \N__28698\ : std_logic;
signal \N__28695\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28684\ : std_logic;
signal \N__28683\ : std_logic;
signal \N__28680\ : std_logic;
signal \N__28677\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28671\ : std_logic;
signal \N__28668\ : std_logic;
signal \N__28665\ : std_logic;
signal \N__28662\ : std_logic;
signal \N__28659\ : std_logic;
signal \N__28656\ : std_logic;
signal \N__28653\ : std_logic;
signal \N__28650\ : std_logic;
signal \N__28645\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28630\ : std_logic;
signal \N__28625\ : std_logic;
signal \N__28624\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28617\ : std_logic;
signal \N__28612\ : std_logic;
signal \N__28609\ : std_logic;
signal \N__28606\ : std_logic;
signal \N__28601\ : std_logic;
signal \N__28598\ : std_logic;
signal \N__28595\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28591\ : std_logic;
signal \N__28588\ : std_logic;
signal \N__28587\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28576\ : std_logic;
signal \N__28571\ : std_logic;
signal \N__28570\ : std_logic;
signal \N__28569\ : std_logic;
signal \N__28566\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28552\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28546\ : std_logic;
signal \N__28543\ : std_logic;
signal \N__28540\ : std_logic;
signal \N__28535\ : std_logic;
signal \N__28532\ : std_logic;
signal \N__28529\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28516\ : std_logic;
signal \N__28513\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28505\ : std_logic;
signal \N__28504\ : std_logic;
signal \N__28503\ : std_logic;
signal \N__28500\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28484\ : std_logic;
signal \N__28483\ : std_logic;
signal \N__28480\ : std_logic;
signal \N__28477\ : std_logic;
signal \N__28472\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28466\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28459\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28452\ : std_logic;
signal \N__28449\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28443\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28435\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28427\ : std_logic;
signal \N__28424\ : std_logic;
signal \N__28421\ : std_logic;
signal \N__28418\ : std_logic;
signal \N__28415\ : std_logic;
signal \N__28412\ : std_logic;
signal \N__28409\ : std_logic;
signal \N__28404\ : std_logic;
signal \N__28401\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28388\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28381\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28377\ : std_logic;
signal \N__28374\ : std_logic;
signal \N__28371\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28362\ : std_logic;
signal \N__28355\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28351\ : std_logic;
signal \N__28350\ : std_logic;
signal \N__28345\ : std_logic;
signal \N__28342\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28334\ : std_logic;
signal \N__28331\ : std_logic;
signal \N__28330\ : std_logic;
signal \N__28327\ : std_logic;
signal \N__28324\ : std_logic;
signal \N__28323\ : std_logic;
signal \N__28318\ : std_logic;
signal \N__28315\ : std_logic;
signal \N__28312\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28305\ : std_logic;
signal \N__28302\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28288\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28277\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28273\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28267\ : std_logic;
signal \N__28266\ : std_logic;
signal \N__28261\ : std_logic;
signal \N__28258\ : std_logic;
signal \N__28255\ : std_logic;
signal \N__28250\ : std_logic;
signal \N__28249\ : std_logic;
signal \N__28248\ : std_logic;
signal \N__28245\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28233\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28227\ : std_logic;
signal \N__28224\ : std_logic;
signal \N__28217\ : std_logic;
signal \N__28214\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28201\ : std_logic;
signal \N__28198\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28187\ : std_logic;
signal \N__28184\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28177\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28165\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28157\ : std_logic;
signal \N__28156\ : std_logic;
signal \N__28155\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28144\ : std_logic;
signal \N__28139\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28132\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28120\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28112\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28107\ : std_logic;
signal \N__28106\ : std_logic;
signal \N__28103\ : std_logic;
signal \N__28100\ : std_logic;
signal \N__28093\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28085\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28078\ : std_logic;
signal \N__28075\ : std_logic;
signal \N__28072\ : std_logic;
signal \N__28071\ : std_logic;
signal \N__28068\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28062\ : std_logic;
signal \N__28059\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28049\ : std_logic;
signal \N__28046\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28044\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28022\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28018\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28012\ : std_logic;
signal \N__28009\ : std_logic;
signal \N__28006\ : std_logic;
signal \N__28005\ : std_logic;
signal \N__28002\ : std_logic;
signal \N__27999\ : std_logic;
signal \N__27996\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27983\ : std_logic;
signal \N__27982\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27980\ : std_logic;
signal \N__27977\ : std_logic;
signal \N__27974\ : std_logic;
signal \N__27971\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27961\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27953\ : std_logic;
signal \N__27952\ : std_logic;
signal \N__27951\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27935\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27922\ : std_logic;
signal \N__27919\ : std_logic;
signal \N__27916\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27910\ : std_logic;
signal \N__27909\ : std_logic;
signal \N__27906\ : std_logic;
signal \N__27903\ : std_logic;
signal \N__27900\ : std_logic;
signal \N__27895\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27889\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27881\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27877\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27851\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27845\ : std_logic;
signal \N__27842\ : std_logic;
signal \N__27839\ : std_logic;
signal \N__27836\ : std_logic;
signal \N__27833\ : std_logic;
signal \N__27830\ : std_logic;
signal \N__27827\ : std_logic;
signal \N__27826\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27818\ : std_logic;
signal \N__27817\ : std_logic;
signal \N__27814\ : std_logic;
signal \N__27811\ : std_logic;
signal \N__27810\ : std_logic;
signal \N__27807\ : std_logic;
signal \N__27804\ : std_logic;
signal \N__27801\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27791\ : std_logic;
signal \N__27790\ : std_logic;
signal \N__27789\ : std_logic;
signal \N__27786\ : std_logic;
signal \N__27783\ : std_logic;
signal \N__27780\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27772\ : std_logic;
signal \N__27769\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27765\ : std_logic;
signal \N__27762\ : std_logic;
signal \N__27759\ : std_logic;
signal \N__27752\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27750\ : std_logic;
signal \N__27747\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27736\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27732\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27726\ : std_logic;
signal \N__27723\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27717\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27702\ : std_logic;
signal \N__27699\ : std_logic;
signal \N__27696\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27683\ : std_logic;
signal \N__27682\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27671\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27665\ : std_logic;
signal \N__27662\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27656\ : std_logic;
signal \N__27653\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27627\ : std_logic;
signal \N__27624\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27618\ : std_logic;
signal \N__27613\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27606\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27598\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27594\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27585\ : std_logic;
signal \N__27580\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27572\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27570\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27550\ : std_logic;
signal \N__27549\ : std_logic;
signal \N__27548\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27524\ : std_logic;
signal \N__27521\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27508\ : std_logic;
signal \N__27505\ : std_logic;
signal \N__27502\ : std_logic;
signal \N__27497\ : std_logic;
signal \N__27494\ : std_logic;
signal \N__27491\ : std_logic;
signal \N__27488\ : std_logic;
signal \N__27485\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27481\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27470\ : std_logic;
signal \N__27469\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27458\ : std_logic;
signal \N__27455\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27446\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27441\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27413\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27407\ : std_logic;
signal \N__27404\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27398\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27392\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27385\ : std_logic;
signal \N__27380\ : std_logic;
signal \N__27379\ : std_logic;
signal \N__27376\ : std_logic;
signal \N__27373\ : std_logic;
signal \N__27368\ : std_logic;
signal \N__27365\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27344\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27332\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27320\ : std_logic;
signal \N__27317\ : std_logic;
signal \N__27314\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27308\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27287\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27281\ : std_logic;
signal \N__27278\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27269\ : std_logic;
signal \N__27266\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27257\ : std_logic;
signal \N__27254\ : std_logic;
signal \N__27251\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27233\ : std_logic;
signal \N__27230\ : std_logic;
signal \N__27227\ : std_logic;
signal \N__27224\ : std_logic;
signal \N__27221\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27208\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27204\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27198\ : std_logic;
signal \N__27195\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27185\ : std_logic;
signal \N__27182\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27173\ : std_logic;
signal \N__27170\ : std_logic;
signal \N__27167\ : std_logic;
signal \N__27164\ : std_logic;
signal \N__27161\ : std_logic;
signal \N__27158\ : std_logic;
signal \N__27155\ : std_logic;
signal \N__27152\ : std_logic;
signal \N__27149\ : std_logic;
signal \N__27146\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27140\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27125\ : std_logic;
signal \N__27122\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27101\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27095\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27089\ : std_logic;
signal \N__27086\ : std_logic;
signal \N__27083\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27079\ : std_logic;
signal \N__27076\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27072\ : std_logic;
signal \N__27069\ : std_logic;
signal \N__27066\ : std_logic;
signal \N__27059\ : std_logic;
signal \N__27058\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27020\ : std_logic;
signal \N__27019\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27013\ : std_logic;
signal \N__27010\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27004\ : std_logic;
signal \N__27001\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26993\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26987\ : std_logic;
signal \N__26984\ : std_logic;
signal \N__26981\ : std_logic;
signal \N__26980\ : std_logic;
signal \N__26977\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26973\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26967\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26959\ : std_logic;
signal \N__26958\ : std_logic;
signal \N__26955\ : std_logic;
signal \N__26952\ : std_logic;
signal \N__26949\ : std_logic;
signal \N__26946\ : std_logic;
signal \N__26945\ : std_logic;
signal \N__26942\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26926\ : std_logic;
signal \N__26921\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26913\ : std_logic;
signal \N__26910\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26897\ : std_logic;
signal \N__26896\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26892\ : std_logic;
signal \N__26889\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26876\ : std_logic;
signal \N__26873\ : std_logic;
signal \N__26872\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26868\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26862\ : std_logic;
signal \N__26859\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26847\ : std_logic;
signal \N__26844\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26825\ : std_logic;
signal \N__26822\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26816\ : std_logic;
signal \N__26813\ : std_logic;
signal \N__26810\ : std_logic;
signal \N__26807\ : std_logic;
signal \N__26804\ : std_logic;
signal \N__26801\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26795\ : std_logic;
signal \N__26792\ : std_logic;
signal \N__26789\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26756\ : std_logic;
signal \N__26753\ : std_logic;
signal \N__26750\ : std_logic;
signal \N__26747\ : std_logic;
signal \N__26744\ : std_logic;
signal \N__26741\ : std_logic;
signal \N__26738\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26729\ : std_logic;
signal \N__26726\ : std_logic;
signal \N__26723\ : std_logic;
signal \N__26720\ : std_logic;
signal \N__26717\ : std_logic;
signal \N__26714\ : std_logic;
signal \N__26711\ : std_logic;
signal \N__26708\ : std_logic;
signal \N__26705\ : std_logic;
signal \N__26702\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26687\ : std_logic;
signal \N__26686\ : std_logic;
signal \N__26683\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26675\ : std_logic;
signal \N__26672\ : std_logic;
signal \N__26669\ : std_logic;
signal \N__26666\ : std_logic;
signal \N__26663\ : std_logic;
signal \N__26660\ : std_logic;
signal \N__26657\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26645\ : std_logic;
signal \N__26642\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26636\ : std_logic;
signal \N__26633\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26621\ : std_logic;
signal \N__26618\ : std_logic;
signal \N__26615\ : std_logic;
signal \N__26612\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26597\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26588\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26582\ : std_logic;
signal \N__26579\ : std_logic;
signal \N__26576\ : std_logic;
signal \N__26573\ : std_logic;
signal \N__26570\ : std_logic;
signal \N__26567\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26546\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26534\ : std_logic;
signal \N__26531\ : std_logic;
signal \N__26528\ : std_logic;
signal \N__26525\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26516\ : std_logic;
signal \N__26513\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26507\ : std_logic;
signal \N__26504\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26495\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26480\ : std_logic;
signal \N__26477\ : std_logic;
signal \N__26474\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26468\ : std_logic;
signal \N__26465\ : std_logic;
signal \N__26462\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26453\ : std_logic;
signal \N__26450\ : std_logic;
signal \N__26447\ : std_logic;
signal \N__26444\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26411\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26359\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26352\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26344\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26331\ : std_logic;
signal \N__26324\ : std_logic;
signal \N__26321\ : std_logic;
signal \N__26318\ : std_logic;
signal \N__26315\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26308\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26297\ : std_logic;
signal \N__26294\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26228\ : std_logic;
signal \N__26225\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26209\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26186\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26181\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26170\ : std_logic;
signal \N__26165\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26158\ : std_logic;
signal \N__26155\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26146\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26137\ : std_logic;
signal \N__26134\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26123\ : std_logic;
signal \N__26122\ : std_logic;
signal \N__26117\ : std_logic;
signal \N__26114\ : std_logic;
signal \N__26111\ : std_logic;
signal \N__26110\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26101\ : std_logic;
signal \N__26100\ : std_logic;
signal \N__26097\ : std_logic;
signal \N__26094\ : std_logic;
signal \N__26091\ : std_logic;
signal \N__26088\ : std_logic;
signal \N__26085\ : std_logic;
signal \N__26078\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26064\ : std_logic;
signal \N__26061\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26053\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26041\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26037\ : std_logic;
signal \N__26034\ : std_logic;
signal \N__26031\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26014\ : std_logic;
signal \N__26011\ : std_logic;
signal \N__26008\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25997\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25987\ : std_logic;
signal \N__25986\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25965\ : std_logic;
signal \N__25960\ : std_logic;
signal \N__25955\ : std_logic;
signal \N__25954\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25950\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25941\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25928\ : std_logic;
signal \N__25927\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25923\ : std_logic;
signal \N__25920\ : std_logic;
signal \N__25917\ : std_logic;
signal \N__25914\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25903\ : std_logic;
signal \N__25900\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25889\ : std_logic;
signal \N__25888\ : std_logic;
signal \N__25885\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25865\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25859\ : std_logic;
signal \N__25856\ : std_logic;
signal \N__25853\ : std_logic;
signal \N__25850\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25846\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25833\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25823\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25821\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25769\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25742\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25719\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25717\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25702\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25694\ : std_logic;
signal \N__25691\ : std_logic;
signal \N__25690\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25688\ : std_logic;
signal \N__25687\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25684\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25671\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25649\ : std_logic;
signal \N__25646\ : std_logic;
signal \N__25643\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25631\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25627\ : std_logic;
signal \N__25624\ : std_logic;
signal \N__25621\ : std_logic;
signal \N__25618\ : std_logic;
signal \N__25615\ : std_logic;
signal \N__25612\ : std_logic;
signal \N__25609\ : std_logic;
signal \N__25606\ : std_logic;
signal \N__25601\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25591\ : std_logic;
signal \N__25588\ : std_logic;
signal \N__25585\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25579\ : std_logic;
signal \N__25576\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25567\ : std_logic;
signal \N__25564\ : std_logic;
signal \N__25561\ : std_logic;
signal \N__25558\ : std_logic;
signal \N__25555\ : std_logic;
signal \N__25552\ : std_logic;
signal \N__25549\ : std_logic;
signal \N__25546\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25532\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25528\ : std_logic;
signal \N__25525\ : std_logic;
signal \N__25522\ : std_logic;
signal \N__25519\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25513\ : std_logic;
signal \N__25510\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25498\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25495\ : std_logic;
signal \N__25494\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25492\ : std_logic;
signal \N__25491\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25488\ : std_logic;
signal \N__25487\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25485\ : std_logic;
signal \N__25484\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25435\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25429\ : std_logic;
signal \N__25426\ : std_logic;
signal \N__25423\ : std_logic;
signal \N__25420\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25412\ : std_logic;
signal \N__25409\ : std_logic;
signal \N__25406\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25397\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25384\ : std_logic;
signal \N__25381\ : std_logic;
signal \N__25378\ : std_logic;
signal \N__25375\ : std_logic;
signal \N__25372\ : std_logic;
signal \N__25369\ : std_logic;
signal \N__25366\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25354\ : std_logic;
signal \N__25351\ : std_logic;
signal \N__25348\ : std_logic;
signal \N__25345\ : std_logic;
signal \N__25342\ : std_logic;
signal \N__25339\ : std_logic;
signal \N__25336\ : std_logic;
signal \N__25333\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25324\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25318\ : std_logic;
signal \N__25315\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25309\ : std_logic;
signal \N__25306\ : std_logic;
signal \N__25303\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25294\ : std_logic;
signal \N__25291\ : std_logic;
signal \N__25288\ : std_logic;
signal \N__25285\ : std_logic;
signal \N__25282\ : std_logic;
signal \N__25279\ : std_logic;
signal \N__25276\ : std_logic;
signal \N__25273\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25265\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25249\ : std_logic;
signal \N__25246\ : std_logic;
signal \N__25243\ : std_logic;
signal \N__25240\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25228\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25192\ : std_logic;
signal \N__25189\ : std_logic;
signal \N__25186\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25177\ : std_logic;
signal \N__25174\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25159\ : std_logic;
signal \N__25156\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25150\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25142\ : std_logic;
signal \N__25139\ : std_logic;
signal \N__25136\ : std_logic;
signal \N__25133\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25114\ : std_logic;
signal \N__25111\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25105\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25097\ : std_logic;
signal \N__25094\ : std_logic;
signal \N__25093\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25087\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25075\ : std_logic;
signal \N__25072\ : std_logic;
signal \N__25071\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25060\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25049\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25043\ : std_logic;
signal \N__25040\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25022\ : std_logic;
signal \N__25019\ : std_logic;
signal \N__25016\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24997\ : std_logic;
signal \N__24994\ : std_logic;
signal \N__24991\ : std_logic;
signal \N__24988\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24971\ : std_logic;
signal \N__24968\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24953\ : std_logic;
signal \N__24950\ : std_logic;
signal \N__24947\ : std_logic;
signal \N__24944\ : std_logic;
signal \N__24941\ : std_logic;
signal \N__24938\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24931\ : std_logic;
signal \N__24926\ : std_logic;
signal \N__24923\ : std_logic;
signal \N__24920\ : std_logic;
signal \N__24917\ : std_logic;
signal \N__24914\ : std_logic;
signal \N__24913\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24907\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24898\ : std_logic;
signal \N__24895\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24881\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24877\ : std_logic;
signal \N__24874\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24860\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24844\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24823\ : std_logic;
signal \N__24820\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24799\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24793\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24781\ : std_logic;
signal \N__24778\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24761\ : std_logic;
signal \N__24758\ : std_logic;
signal \N__24755\ : std_logic;
signal \N__24752\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24724\ : std_logic;
signal \N__24721\ : std_logic;
signal \N__24718\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24686\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24667\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24656\ : std_logic;
signal \N__24653\ : std_logic;
signal \N__24650\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24625\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24619\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24598\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24592\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24571\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24563\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24554\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24541\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24532\ : std_logic;
signal \N__24529\ : std_logic;
signal \N__24526\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24499\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24482\ : std_logic;
signal \N__24479\ : std_logic;
signal \N__24476\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24455\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24439\ : std_logic;
signal \N__24436\ : std_logic;
signal \N__24433\ : std_logic;
signal \N__24430\ : std_logic;
signal \N__24425\ : std_logic;
signal \N__24422\ : std_logic;
signal \N__24419\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24403\ : std_logic;
signal \N__24402\ : std_logic;
signal \N__24397\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24391\ : std_logic;
signal \N__24386\ : std_logic;
signal \N__24383\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24374\ : std_logic;
signal \N__24373\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24356\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24346\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24331\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24316\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24296\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24281\ : std_logic;
signal \N__24278\ : std_logic;
signal \N__24275\ : std_logic;
signal \N__24272\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24245\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24200\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24182\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24161\ : std_logic;
signal \N__24158\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24146\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24134\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24125\ : std_logic;
signal \N__24122\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24116\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24110\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24090\ : std_logic;
signal \N__24087\ : std_logic;
signal \N__24080\ : std_logic;
signal \N__24079\ : std_logic;
signal \N__24076\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24070\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24064\ : std_logic;
signal \N__24061\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24053\ : std_logic;
signal \N__24050\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24031\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24015\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23995\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23947\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23937\ : std_logic;
signal \N__23934\ : std_logic;
signal \N__23931\ : std_logic;
signal \N__23924\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23916\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23904\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23896\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23884\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23817\ : std_logic;
signal \N__23814\ : std_logic;
signal \N__23811\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23791\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23781\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23754\ : std_logic;
signal \N__23751\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23725\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23710\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23700\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23672\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23569\ : std_logic;
signal \N__23566\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23562\ : std_logic;
signal \N__23559\ : std_logic;
signal \N__23556\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23530\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23505\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23443\ : std_logic;
signal \N__23440\ : std_logic;
signal \N__23437\ : std_logic;
signal \N__23434\ : std_logic;
signal \N__23431\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23416\ : std_logic;
signal \N__23413\ : std_logic;
signal \N__23410\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23291\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23287\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23256\ : std_logic;
signal \N__23255\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23235\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23223\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23190\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23187\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23181\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23165\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23082\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23076\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23050\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23044\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22990\ : std_logic;
signal \N__22977\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22955\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22931\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22905\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22873\ : std_logic;
signal \N__22870\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22851\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22837\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22811\ : std_logic;
signal \N__22808\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22791\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22782\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22767\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22732\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22728\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22718\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22658\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22629\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22626\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22602\ : std_logic;
signal \N__22599\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22566\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22515\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22485\ : std_logic;
signal \N__22482\ : std_logic;
signal \N__22479\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22417\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22381\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22211\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22148\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22130\ : std_logic;
signal \N__22127\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22029\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21597\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21590\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21575\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21567\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21536\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21515\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21492\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21480\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21435\ : std_logic;
signal \N__21432\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21393\ : std_logic;
signal \N__21390\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21364\ : std_logic;
signal \N__21363\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21333\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21314\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21309\ : std_logic;
signal \N__21306\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21285\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21272\ : std_logic;
signal \N__21269\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21241\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21188\ : std_logic;
signal \N__21187\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21068\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21027\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21010\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21006\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20973\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20884\ : std_logic;
signal \N__20881\ : std_logic;
signal \N__20880\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20871\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20835\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20821\ : std_logic;
signal \N__20818\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20791\ : std_logic;
signal \N__20788\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20784\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20747\ : std_logic;
signal \N__20744\ : std_logic;
signal \N__20741\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20729\ : std_logic;
signal \N__20726\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20683\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20645\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20575\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20567\ : std_logic;
signal \N__20564\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20511\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20478\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20451\ : std_logic;
signal \N__20448\ : std_logic;
signal \N__20445\ : std_logic;
signal \N__20442\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20383\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20376\ : std_logic;
signal \N__20373\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20353\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20347\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20308\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20290\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20251\ : std_logic;
signal \N__20248\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20233\ : std_logic;
signal \N__20230\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20017\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19993\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19804\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19800\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19699\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19675\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19654\ : std_logic;
signal \N__19653\ : std_logic;
signal \N__19650\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19636\ : std_logic;
signal \N__19635\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19617\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19611\ : std_logic;
signal \N__19608\ : std_logic;
signal \N__19605\ : std_logic;
signal \N__19602\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19584\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19485\ : std_logic;
signal \N__19482\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19464\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19166\ : std_logic;
signal \N__19163\ : std_logic;
signal \N__19160\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19091\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19079\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19052\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19034\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19028\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18974\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18956\ : std_logic;
signal \N__18953\ : std_logic;
signal \N__18950\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18866\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18752\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18734\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18729\ : std_logic;
signal \N__18722\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18686\ : std_logic;
signal \N__18683\ : std_logic;
signal \N__18680\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18661\ : std_logic;
signal \N__18660\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18657\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18652\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18631\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18625\ : std_logic;
signal \N__18622\ : std_logic;
signal \N__18621\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18609\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18580\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18542\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18458\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18350\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18311\ : std_logic;
signal delay_tr_input_ibuf_gb_io_gb_input : std_logic;
signal delay_hc_input_ibuf_gb_io_gb_input : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_15\ : std_logic;
signal \bfn_1_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_8\ : std_logic;
signal \bfn_1_14_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_97\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_91\ : std_logic;
signal \N_42_i_i\ : std_logic;
signal un7_start_stop_0_a2 : std_logic;
signal \bfn_2_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_9\ : std_logic;
signal \bfn_2_14_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_17\ : std_logic;
signal \bfn_2_15_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_25\ : std_logic;
signal \bfn_2_16_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_159\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_96\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_96_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_3\ : std_logic;
signal pwm_duty_input_0 : std_logic;
signal pwm_duty_input_1 : std_logic;
signal pwm_duty_input_2 : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\ : std_logic;
signal \pwm_generator_inst.un1_duty_inputlt3\ : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_\ : std_logic;
signal pwm_duty_input_9 : std_logic;
signal pwm_duty_input_7 : std_logic;
signal pwm_duty_input_6 : std_logic;
signal pwm_duty_input_8 : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\ : std_logic;
signal \bfn_3_17_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\ : std_logic;
signal \bfn_3_18_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\ : std_logic;
signal \bfn_3_19_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\ : std_logic;
signal \bfn_3_20_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto3\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_98\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_27\ : std_logic;
signal pwm_duty_input_3 : std_logic;
signal pwm_duty_input_4 : std_logic;
signal pwm_duty_input_5 : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\ : std_logic;
signal \bfn_3_24_0_\ : std_logic;
signal \pwm_generator_inst.O_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_0\ : std_logic;
signal \pwm_generator_inst.O_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_1\ : std_logic;
signal \pwm_generator_inst.O_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_2\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_3\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_4\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_5\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_6\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_7\ : std_logic;
signal \bfn_3_25_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_9\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_15\ : std_logic;
signal \bfn_3_26_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_16\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_17\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_77_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_43\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_axbZ0Z_4\ : std_logic;
signal \bfn_4_23_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_18\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_20\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_5\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_21\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_6\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_22\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_7\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_23\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0\ : std_logic;
signal \bfn_4_24_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_24\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\ : std_logic;
signal \bfn_4_25_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81_cascade_\ : std_logic;
signal \pwm_generator_inst.O_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_16_cascade_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.runningZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_47\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_44_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_46\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\ : std_logic;
signal \pwm_generator_inst.O_0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_0\ : std_logic;
signal \bfn_5_25_0_\ : std_logic;
signal \pwm_generator_inst.O_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_0\ : std_logic;
signal \pwm_generator_inst.O_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_1\ : std_logic;
signal \pwm_generator_inst.O_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_2\ : std_logic;
signal \pwm_generator_inst.O_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_3\ : std_logic;
signal \pwm_generator_inst.O_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_4\ : std_logic;
signal \pwm_generator_inst.O_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_5\ : std_logic;
signal \pwm_generator_inst.O_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_7\ : std_logic;
signal \pwm_generator_inst.O_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_8\ : std_logic;
signal \bfn_5_26_0_\ : std_logic;
signal \pwm_generator_inst.O_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un3_threshold\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_15\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\ : std_logic;
signal \bfn_5_27_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18\ : std_logic;
signal \elapsed_time_ns_1_RNIH33T9_0_5_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_df30_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latchedZ0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_0\ : std_logic;
signal \bfn_7_23_0_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_7\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_7\ : std_logic;
signal \bfn_7_24_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_8\ : std_logic;
signal il_max_comp1_c : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\ : std_logic;
signal \bfn_8_5_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3Z0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \bfn_8_6_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_8_7_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\ : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_8_9_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_8_10_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_16\ : std_logic;
signal \bfn_8_11_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\ : std_logic;
signal \elapsed_time_ns_1_RNI58DN9_0_27_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axb_0\ : std_logic;
signal \bfn_8_19_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_8\ : std_logic;
signal \bfn_8_20_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_14\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93\ : std_logic;
signal \pwm_generator_inst.N_17\ : std_logic;
signal \pwm_generator_inst.N_16\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt18\ : std_logic;
signal \elapsed_time_ns_1_RNI57CN9_0_18_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\ : std_logic;
signal \elapsed_time_ns_1_RNI24CN9_0_15_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \elapsed_time_ns_1_RNIE03T9_0_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\ : std_logic;
signal \elapsed_time_ns_1_RNIF13T9_0_3\ : std_logic;
signal \elapsed_time_ns_1_RNIH33T9_0_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22\ : std_logic;
signal \elapsed_time_ns_1_RNI14DN9_0_23_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_23\ : std_logic;
signal \elapsed_time_ns_1_RNI03DN9_0_22_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_22\ : std_logic;
signal \elapsed_time_ns_1_RNIG23T9_0_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \elapsed_time_ns_1_RNI03DN9_0_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_22\ : std_logic;
signal \elapsed_time_ns_1_RNI14DN9_0_23\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNITUBN9_0_10\ : std_logic;
signal \elapsed_time_ns_1_RNITUBN9_0_10_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3\ : std_logic;
signal \elapsed_time_ns_1_RNIL73T9_0_9_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\ : std_logic;
signal \elapsed_time_ns_1_RNIUVBN9_0_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\ : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_7\ : std_logic;
signal \bfn_9_16_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_15\ : std_logic;
signal \bfn_9_17_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_23\ : std_logic;
signal \bfn_9_18_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_28\ : std_logic;
signal \current_shift_inst.control_input_18\ : std_logic;
signal \bfn_9_19_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\ : std_logic;
signal \current_shift_inst.control_input_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\ : std_logic;
signal \current_shift_inst.control_input_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\ : std_logic;
signal \current_shift_inst.control_input_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\ : std_logic;
signal \current_shift_inst.control_input_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\ : std_logic;
signal \current_shift_inst.control_input_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\ : std_logic;
signal \current_shift_inst.control_input_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\ : std_logic;
signal \current_shift_inst.control_input_cry_6\ : std_logic;
signal \current_shift_inst.control_input_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\ : std_logic;
signal \bfn_9_20_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\ : std_logic;
signal \current_shift_inst.control_input_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\ : std_logic;
signal \current_shift_inst.control_input_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\ : std_logic;
signal \current_shift_inst.control_input_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\ : std_logic;
signal \current_shift_inst.control_input_cry_11\ : std_logic;
signal \current_shift_inst.control_input_cry_12\ : std_logic;
signal \current_shift_inst.control_input_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\ : std_logic;
signal \pwm_generator_inst.threshold_0\ : std_logic;
signal \pwm_generator_inst.counter_i_0\ : std_logic;
signal \bfn_9_24_0_\ : std_logic;
signal \pwm_generator_inst.un14_counter_1\ : std_logic;
signal \pwm_generator_inst.counter_i_1\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_0\ : std_logic;
signal \pwm_generator_inst.threshold_2\ : std_logic;
signal \pwm_generator_inst.counter_i_2\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_1\ : std_logic;
signal \pwm_generator_inst.threshold_3\ : std_logic;
signal \pwm_generator_inst.counter_i_3\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_2\ : std_logic;
signal \pwm_generator_inst.threshold_4\ : std_logic;
signal \pwm_generator_inst.counter_i_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_3\ : std_logic;
signal \pwm_generator_inst.threshold_5\ : std_logic;
signal \pwm_generator_inst.counter_i_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_6\ : std_logic;
signal \pwm_generator_inst.counter_i_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_7\ : std_logic;
signal \pwm_generator_inst.counter_i_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_8\ : std_logic;
signal \pwm_generator_inst.counter_i_8\ : std_logic;
signal \bfn_9_25_0_\ : std_logic;
signal \pwm_generator_inst.threshold_9\ : std_logic;
signal \pwm_generator_inst.counter_i_9\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_8\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_9\ : std_logic;
signal pwm_output_c : std_logic;
signal s3_phy_c : std_logic;
signal \elapsed_time_ns_1_RNI68CN9_0_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \elapsed_time_ns_1_RNIL73T9_0_9\ : std_logic;
signal \elapsed_time_ns_1_RNI57CN9_0_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \elapsed_time_ns_1_RNIDV2T9_0_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\ : std_logic;
signal \elapsed_time_ns_1_RNI25DN9_0_24\ : std_logic;
signal \elapsed_time_ns_1_RNI46CN9_0_17\ : std_logic;
signal \elapsed_time_ns_1_RNII43T9_0_6\ : std_logic;
signal \elapsed_time_ns_1_RNI13CN9_0_14\ : std_logic;
signal \elapsed_time_ns_1_RNI36DN9_0_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_10_7_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_10_8_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt18\ : std_logic;
signal \bfn_10_9_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24\ : std_logic;
signal \elapsed_time_ns_1_RNIV0CN9_0_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt26\ : std_logic;
signal \elapsed_time_ns_1_RNI58DN9_0_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_29\ : std_logic;
signal \elapsed_time_ns_1_RNI04EN9_0_31\ : std_logic;
signal \elapsed_time_ns_1_RNIV2EN9_0_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\ : std_logic;
signal \bfn_10_12_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\ : std_logic;
signal \bfn_10_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\ : std_logic;
signal \bfn_10_14_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\ : std_logic;
signal \bfn_10_15_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_202_i\ : std_logic;
signal \elapsed_time_ns_1_RNIK63T9_0_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_203_i\ : std_logic;
signal \il_max_comp1_D1\ : std_logic;
signal \current_shift_inst.control_input_axb_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.running_i\ : std_logic;
signal \current_shift_inst.control_input_axb_12\ : std_logic;
signal \current_shift_inst.N_1304_i\ : std_logic;
signal \pwm_generator_inst.un1_counterlto2_0_cascade_\ : std_logic;
signal \pwm_generator_inst.un1_counterlt9_cascade_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_0\ : std_logic;
signal \bfn_10_24_0_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_1\ : std_logic;
signal \pwm_generator_inst.counter_cry_0\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_3\ : std_logic;
signal \pwm_generator_inst.counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_5\ : std_logic;
signal \pwm_generator_inst.counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counter_cry_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_7\ : std_logic;
signal \bfn_10_25_0_\ : std_logic;
signal \pwm_generator_inst.un1_counter_0\ : std_logic;
signal \pwm_generator_inst.counter_cry_8\ : std_logic;
signal \elapsed_time_ns_1_RNI35CN9_0_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\ : std_logic;
signal \elapsed_time_ns_1_RNI24CN9_0_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_df30_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_11_8_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3Z0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \bfn_11_10_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\ : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\ : std_logic;
signal \elapsed_time_ns_1_RNI02CN9_0_13\ : std_logic;
signal start_stop_c : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\ : std_logic;
signal \elapsed_time_ns_1_RNI47DN9_0_26\ : std_logic;
signal \delay_measurement_inst.start_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_trZ0\ : std_logic;
signal delay_tr_input_c_g : std_logic;
signal \pwm_generator_inst.counterZ0Z_9\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_8\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_7\ : std_logic;
signal \pwm_generator_inst.un1_counterlto9_2\ : std_logic;
signal \delay_measurement_inst.stop_timer_hcZ0\ : std_logic;
signal clk_12mhz : std_logic;
signal \GB_BUFFER_clk_12mhz_THRU_CO\ : std_logic;
signal \phase_controller_inst2.start_timer_tr_RNO_0_0\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst2.start_timer_hc_0_sqmuxa\ : std_logic;
signal \phase_controller_inst2.state_RNIG7JFZ0Z_2\ : std_logic;
signal il_min_comp2_c : std_logic;
signal il_max_comp2_c : std_logic;
signal \phase_controller_inst2.stateZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\ : std_logic;
signal \elapsed_time_ns_1_RNI69DN9_0_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt28\ : std_logic;
signal \elapsed_time_ns_1_RNI7ADN9_0_29\ : std_logic;
signal \elapsed_time_ns_1_RNI7ADN9_0_29_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28\ : std_logic;
signal \elapsed_time_ns_1_RNIJ53T9_0_7_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_20\ : std_logic;
signal \elapsed_time_ns_1_RNIV1DN9_0_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\ : std_logic;
signal \elapsed_time_ns_1_RNIJ53T9_0_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_start_g\ : std_logic;
signal \phase_controller_inst2.hc_time_passed\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_start_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.runningZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un2_start_0\ : std_logic;
signal \phase_controller_inst2.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latchedZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3\ : std_logic;
signal \elapsed_time_ns_1_RNIU0DN9_0_20\ : std_logic;
signal \current_shift_inst.un4_control_input1_1_cascade_\ : std_logic;
signal \bfn_12_15_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s1\ : std_logic;
signal \bfn_12_16_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s1\ : std_logic;
signal \bfn_12_17_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s1\ : std_logic;
signal \bfn_12_18_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s1\ : std_logic;
signal il_min_comp1_c : std_logic;
signal \il_min_comp1_D1\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_1\ : std_logic;
signal s4_phy_c : std_logic;
signal \delay_measurement_inst.start_timer_hcZ0\ : std_logic;
signal delay_hc_input_c_g : std_logic;
signal \pll_inst.red_c_i\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_0\ : std_logic;
signal \phase_controller_inst2.state_RNI9M3OZ0Z_0\ : std_logic;
signal \phase_controller_inst2.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst2.tr_time_passed\ : std_logic;
signal \phase_controller_inst2.stoper_tr.runningZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latchedZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un2_start_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_df30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_30\ : std_logic;
signal \elapsed_time_ns_1_RNI0AOBB_0_13_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_31\ : std_logic;
signal \bfn_13_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_7\ : std_logic;
signal \bfn_13_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_15\ : std_logic;
signal \bfn_13_12_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_23\ : std_logic;
signal \bfn_13_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_205_i\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_fast_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.running_i\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_21\ : std_logic;
signal \current_shift_inst.control_input_axb_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_22\ : std_logic;
signal \current_shift_inst.control_input_axb_2\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_23\ : std_logic;
signal \current_shift_inst.control_input_axb_3\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_24\ : std_logic;
signal \current_shift_inst.control_input_axb_4\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_25\ : std_logic;
signal \current_shift_inst.control_input_axb_5\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_26\ : std_logic;
signal \current_shift_inst.control_input_axb_6\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_27\ : std_logic;
signal \current_shift_inst.control_input_axb_7\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_28\ : std_logic;
signal \current_shift_inst.control_input_axb_8\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_29\ : std_logic;
signal \current_shift_inst.control_input_axb_9\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_30\ : std_logic;
signal \current_shift_inst.control_input_axb_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\ : std_logic;
signal state_ns_i_a2_1 : std_logic;
signal \phase_controller_inst1.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst1.start_timer_hc_0_sqmuxa\ : std_logic;
signal \il_max_comp1_D2\ : std_logic;
signal \current_shift_inst.timer_s1.N_162_i\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\ : std_logic;
signal \bfn_14_8_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34Z0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \bfn_14_9_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_14_10_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\ : std_logic;
signal \bfn_14_11_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\ : std_logic;
signal \elapsed_time_ns_1_RNIVAQBB_0_30\ : std_logic;
signal \elapsed_time_ns_1_RNIVAQBB_0_30_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI0CQBB_0_31\ : std_logic;
signal \elapsed_time_ns_1_RNI0CQBB_0_31_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI0AOBB_0_13\ : std_logic;
signal \current_shift_inst.un38_control_input_5_0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0_sf\ : std_logic;
signal \bfn_14_13_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s0\ : std_logic;
signal \bfn_14_14_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s0\ : std_logic;
signal \bfn_14_15_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_24\ : std_logic;
signal \bfn_14_16_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_25\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_31\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s0\ : std_logic;
signal \current_shift_inst.control_input_axb_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\ : std_logic;
signal phase_controller_inst1_state_4 : std_logic;
signal \phase_controller_inst1.time_passed_RNIE87F\ : std_logic;
signal \phase_controller_inst1.hc_time_passed\ : std_logic;
signal \il_min_comp1_D2\ : std_logic;
signal \phase_controller_inst1.start_timer_tr_RNOZ0Z_0\ : std_logic;
signal \current_shift_inst.timer_s1.runningZ0\ : std_logic;
signal \current_shift_inst.start_timer_sZ0Z1\ : std_logic;
signal s1_phy_c : std_logic;
signal \current_shift_inst.stop_timer_sZ0Z1\ : std_logic;
signal s2_phy_c : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_15_7_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_15_8_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt18\ : std_logic;
signal \bfn_15_9_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\ : std_logic;
signal \bfn_15_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\ : std_logic;
signal \bfn_15_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\ : std_logic;
signal \bfn_15_12_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\ : std_logic;
signal \bfn_15_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_204_i\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\ : std_logic;
signal \bfn_15_18_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \bfn_15_19_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \bfn_15_20_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \bfn_15_21_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \T12_c\ : std_logic;
signal \T45_c\ : std_logic;
signal state_3 : std_logic;
signal \phase_controller_inst1.stateZ0Z_2\ : std_logic;
signal \T01_c\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_1\ : std_logic;
signal \T23_c\ : std_logic;
signal \elapsed_time_ns_1_RNIHG91B_0_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \elapsed_time_ns_1_RNIU7OBB_0_11\ : std_logic;
signal \elapsed_time_ns_1_RNIU7OBB_0_11_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIT6OBB_0_10\ : std_logic;
signal \elapsed_time_ns_1_RNIT6OBB_0_10_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_20\ : std_logic;
signal \elapsed_time_ns_1_RNIDC91B_0_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\ : std_logic;
signal \elapsed_time_ns_1_RNIGF91B_0_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_16_11_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_16_12_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_16\ : std_logic;
signal \bfn_16_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\ : std_logic;
signal \bfn_16_14_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7\ : std_logic;
signal \bfn_16_15_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15\ : std_logic;
signal \bfn_16_16_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23\ : std_logic;
signal \bfn_16_17_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\ : std_logic;
signal \phase_controller_inst1.tr_time_passed\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.time_passed_RNI7NN7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\ : std_logic;
signal \elapsed_time_ns_1_RNIED91B_0_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\ : std_logic;
signal \elapsed_time_ns_1_RNIFE91B_0_3\ : std_logic;
signal \elapsed_time_ns_1_RNIIH91B_0_6\ : std_logic;
signal \elapsed_time_ns_1_RNIV9PBB_0_21\ : std_logic;
signal \elapsed_time_ns_1_RNIV9PBB_0_21_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22\ : std_logic;
signal \elapsed_time_ns_1_RNI0BPBB_0_22\ : std_logic;
signal \elapsed_time_ns_1_RNI0BPBB_0_22_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \elapsed_time_ns_1_RNIKJ91B_0_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\ : std_logic;
signal \elapsed_time_ns_1_RNIU8PBB_0_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\ : std_logic;
signal \elapsed_time_ns_1_RNIJI91B_0_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\ : std_logic;
signal \elapsed_time_ns_1_RNIV8OBB_0_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_17_10_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_17_11_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_17_12_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\ : std_logic;
signal \bfn_17_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_10\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_9\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_5\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_8\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_3\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_4\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_6\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_14\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_13\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_11\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_12\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_16\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_17\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_26\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_23\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_24\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_19\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_25\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_28\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_27\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_0\ : std_logic;
signal \bfn_17_18_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_0\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_2\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_1\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_3\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_4\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_5\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_7\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_8\ : std_logic;
signal \bfn_17_19_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_10\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_11\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_12\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_13\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_15\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_16\ : std_logic;
signal \bfn_17_20_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_17\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_18\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_19\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_20\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_21\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_23\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_24\ : std_logic;
signal \bfn_17_21_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_25\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_26\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_27\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_28\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.running_i\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_29\ : std_logic;
signal \current_shift_inst.timer_s1.N_163_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21\ : std_logic;
signal \elapsed_time_ns_1_RNILK91B_0_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \elapsed_time_ns_1_RNI4EOBB_0_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\ : std_logic;
signal \elapsed_time_ns_1_RNI1CPBB_0_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\ : std_logic;
signal \elapsed_time_ns_1_RNI1BOBB_0_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\ : std_logic;
signal \elapsed_time_ns_1_RNI3DOBB_0_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_start_0_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4Z0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.runningZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_df30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_start_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\ : std_logic;
signal \elapsed_time_ns_1_RNI6GOBB_0_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \elapsed_time_ns_1_RNI5FOBB_0_18\ : std_logic;
signal \elapsed_time_ns_1_RNI5FOBB_0_18_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\ : std_logic;
signal \elapsed_time_ns_1_RNI2COBB_0_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \current_shift_inst.un38_control_input_axb_31_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31_rep1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1\ : std_logic;
signal \bfn_18_14_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.un4_control_input1_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_3\ : std_logic;
signal \current_shift_inst.un4_control_input1_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.un4_control_input1_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.un4_control_input1_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_7\ : std_logic;
signal \current_shift_inst.un4_control_input1_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.un4_control_input1_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_9\ : std_logic;
signal \current_shift_inst.un4_control_input1_10\ : std_logic;
signal \bfn_18_15_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_10\ : std_logic;
signal \current_shift_inst.un4_control_input1_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_11\ : std_logic;
signal \current_shift_inst.un4_control_input1_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_12\ : std_logic;
signal \current_shift_inst.un4_control_input1_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_13\ : std_logic;
signal \current_shift_inst.un4_control_input1_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_12\ : std_logic;
signal \current_shift_inst.un4_control_input1_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_15\ : std_logic;
signal \current_shift_inst.un4_control_input1_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_16\ : std_logic;
signal \current_shift_inst.un4_control_input1_17\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_16\ : std_logic;
signal \current_shift_inst.un4_control_input1_18\ : std_logic;
signal \bfn_18_16_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_18\ : std_logic;
signal \current_shift_inst.un4_control_input1_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_17\ : std_logic;
signal \current_shift_inst.un4_control_input1_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_20\ : std_logic;
signal \current_shift_inst.un4_control_input1_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_21\ : std_logic;
signal \current_shift_inst.un4_control_input1_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_22\ : std_logic;
signal \current_shift_inst.un4_control_input1_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_23\ : std_logic;
signal \current_shift_inst.un4_control_input1_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_24\ : std_logic;
signal \current_shift_inst.un4_control_input1_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_25\ : std_logic;
signal \current_shift_inst.un4_control_input1_26\ : std_logic;
signal \bfn_18_17_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_26\ : std_logic;
signal \current_shift_inst.un4_control_input1_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_27\ : std_logic;
signal \current_shift_inst.un4_control_input1_28\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_29\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_27\ : std_logic;
signal \current_shift_inst.un4_control_input1_30\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_31\ : std_logic;
signal \current_shift_inst.un4_control_input1_31_THRU_CO_cascade_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_7\ : std_logic;
signal \current_shift_inst.un4_control_input1_7\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_1\ : std_logic;
signal \current_shift_inst.timer_s1.N_162_i_g\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_2\ : std_logic;
signal \current_shift_inst.un38_control_input_5_1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_31_THRU_CO\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31\ : std_logic;
signal \current_shift_inst.un38_control_input_5_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_30\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un8_enablelto31\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\ : std_logic;
signal \elapsed_time_ns_1_RNI6HPBB_0_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt26\ : std_logic;
signal \phase_controller_inst1.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latchedZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_start_g\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\ : std_logic;
signal \elapsed_time_ns_1_RNI7IPBB_0_29\ : std_logic;
signal \elapsed_time_ns_1_RNI2DPBB_0_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\ : std_logic;
signal \elapsed_time_ns_1_RNI4FPBB_0_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\ : std_logic;
signal \elapsed_time_ns_1_RNI5GPBB_0_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\ : std_logic;
signal \elapsed_time_ns_1_RNI3EPBB_0_25\ : std_logic;
signal clk_100mhz_0 : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\ : std_logic;
signal red_c_g : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1_15\ : std_logic;
signal \N_19_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_25\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal reset_wire : std_logic;
signal \T01_wire\ : std_logic;
signal start_stop_wire : std_logic;
signal il_max_comp2_wire : std_logic;
signal \T23_wire\ : std_logic;
signal pwm_output_wire : std_logic;
signal il_max_comp1_wire : std_logic;
signal s2_phy_wire : std_logic;
signal \T12_wire\ : std_logic;
signal il_min_comp2_wire : std_logic;
signal s1_phy_wire : std_logic;
signal s4_phy_wire : std_logic;
signal il_min_comp1_wire : std_logic;
signal s3_phy_wire : std_logic;
signal \T45_wire\ : std_logic;
signal delay_hc_input_wire : std_logic;
signal delay_tr_input_wire : std_logic;
signal rgb_b_wire : std_logic;
signal rgb_g_wire : std_logic;
signal rgb_r_wire : std_logic;
signal \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\ : std_logic_vector(31 downto 0);

begin
    reset_wire <= reset;
    T01 <= \T01_wire\;
    start_stop_wire <= start_stop;
    il_max_comp2_wire <= il_max_comp2;
    T23 <= \T23_wire\;
    pwm_output <= pwm_output_wire;
    il_max_comp1_wire <= il_max_comp1;
    s2_phy <= s2_phy_wire;
    T12 <= \T12_wire\;
    il_min_comp2_wire <= il_min_comp2;
    s1_phy <= s1_phy_wire;
    s4_phy <= s4_phy_wire;
    il_min_comp1_wire <= il_min_comp1;
    s3_phy <= s3_phy_wire;
    T45 <= \T45_wire\;
    delay_hc_input_wire <= delay_hc_input;
    delay_tr_input_wire <= delay_tr_input;
    rgb_b <= rgb_b_wire;
    rgb_g <= rgb_g_wire;
    rgb_r <= rgb_r_wire;
    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\ <= \N__25490\&\N__25498\&\N__25489\&\N__25496\&\N__25488\&\N__25495\&\N__25487\&\N__25497\&\N__25484\&\N__25491\&\N__25483\&\N__25492\&\N__25486\&\N__25493\&\N__25485\&\N__25494\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__37929\&'0'&\N__37928\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(15);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_14\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(14);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_13\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(13);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_12\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(12);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_11\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(11);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_10\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(10);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_9\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(9);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_8\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(8);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_7\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(7);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_6\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(6);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_5\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(5);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_4\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(4);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_3\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(3);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_2\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(2);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_1\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(1);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_0\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\ <= '0'&\N__46183\&\N__46176\&\N__46181\&\N__46175\&\N__46182\&\N__46174\&\N__46184\&\N__46171\&\N__46177\&\N__46170\&\N__46178\&\N__46172\&\N__46179\&\N__46173\&\N__46180\;
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__37903\&\N__37900\&'0'&'0'&'0'&\N__37898\&\N__37902\&\N__37899\&\N__37901\;
    \pwm_generator_inst.un2_threshold_2_1_16\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_2_1_15\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.un2_threshold_2_14\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.un2_threshold_2_13\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.un2_threshold_2_12\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un2_threshold_2_11\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.un2_threshold_2_10\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.un2_threshold_2_9\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.un2_threshold_2_8\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.un2_threshold_2_7\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.un2_threshold_2_6\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.un2_threshold_2_5\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.un2_threshold_2_4\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.un2_threshold_2_3\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.un2_threshold_2_2\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.un2_threshold_2_1\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.un2_threshold_2_0\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\ <= '0'&\N__46231\&\N__46234\&\N__46232\&\N__46235\&\N__46233\&\N__19655\&\N__19593\&\N__19637\&\N__19618\&\N__20281\&\N__20309\&\N__20338\&\N__19685\&\N__19700\&\N__19718\;
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__37829\&\N__37826\&'0'&'0'&'0'&\N__37824\&\N__37828\&\N__37825\&\N__37827\;
    \pwm_generator_inst.un2_threshold_1_25\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(25);
    \pwm_generator_inst.un2_threshold_1_24\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(24);
    \pwm_generator_inst.un2_threshold_1_23\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(23);
    \pwm_generator_inst.un2_threshold_1_22\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(22);
    \pwm_generator_inst.un2_threshold_1_21\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(21);
    \pwm_generator_inst.un2_threshold_1_20\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(20);
    \pwm_generator_inst.un2_threshold_1_19\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(19);
    \pwm_generator_inst.un2_threshold_1_18\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(18);
    \pwm_generator_inst.un2_threshold_1_17\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(17);
    \pwm_generator_inst.un2_threshold_1_16\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_1_15\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.O_14\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.O_13\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.O_12\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un3_threshold\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.O_10\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.O_9\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.O_8\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.O_7\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.O_6\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.O_5\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.O_4\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.O_3\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.O_2\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.O_1\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.O_0\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(0);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\ <= '0'&\N__25499\&\N__25538\&\N__25568\&\N__25598\&\N__25631\&\N__25136\&\N__25166\&\N__25199\&\N__25232\&\N__25265\&\N__25295\&\N__25325\&\N__25355\&\N__25384\&\N__24998\;
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__37978\&'0'&\N__37977\;
    \current_shift_inst.PI_CTRL.integrator_1_0_1_19\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(19);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_18\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(18);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_17\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(17);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_16\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(16);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(15);
    \current_shift_inst.PI_CTRL.integrator_1_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(14);
    \current_shift_inst.PI_CTRL.integrator_1_14\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(13);
    \current_shift_inst.PI_CTRL.integrator_1_13\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(12);
    \current_shift_inst.PI_CTRL.integrator_1_12\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(11);
    \current_shift_inst.PI_CTRL.integrator_1_11\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(10);
    \current_shift_inst.PI_CTRL.integrator_1_10\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(9);
    \current_shift_inst.PI_CTRL.integrator_1_9\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(8);
    \current_shift_inst.PI_CTRL.integrator_1_8\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(7);
    \current_shift_inst.PI_CTRL.integrator_1_7\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(6);
    \current_shift_inst.PI_CTRL.integrator_1_6\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(5);
    \current_shift_inst.PI_CTRL.integrator_1_5\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(4);
    \current_shift_inst.PI_CTRL.integrator_1_4\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(3);
    \current_shift_inst.PI_CTRL.integrator_1_3\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(2);
    \current_shift_inst.PI_CTRL.integrator_1_2\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(1);
    \current_shift_inst.PI_CTRL.un1_integrator\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(0);

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__30875\,
            RESETB => \N__32915\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => clk_100mhz_0
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__37930\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__37905\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\,
            ADDSUBBOT => '0',
            A => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\,
            C => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\,
            B => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\,
            OHOLDTOP => '0',
            O => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__37904\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__37897\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__37980\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__37823\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__37979\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__37976\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\,
            ADDSUBBOT => '0',
            A => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\,
            C => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\,
            B => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\,
            OHOLDTOP => '0',
            O => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\
        );

    \reset_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__48450\,
            GLOBALBUFFEROUTPUT => red_c_g
        );

    \reset_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48452\,
            DIN => \N__48451\,
            DOUT => \N__48450\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48452\,
            PADOUT => \N__48451\,
            PADIN => \N__48450\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T01_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48441\,
            DIN => \N__48440\,
            DOUT => \N__48439\,
            PACKAGEPIN => \T01_wire\
        );

    \T01_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48441\,
            PADOUT => \N__48440\,
            PADIN => \N__48439\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__36608\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \start_stop_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48432\,
            DIN => \N__48431\,
            DOUT => \N__48430\,
            PACKAGEPIN => start_stop_wire
        );

    \start_stop_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48432\,
            PADOUT => \N__48431\,
            PADIN => \N__48430\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => start_stop_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48423\,
            DIN => \N__48422\,
            DOUT => \N__48421\,
            PACKAGEPIN => il_max_comp2_wire
        );

    \il_max_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48423\,
            PADOUT => \N__48422\,
            PADIN => \N__48421\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T23_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48414\,
            DIN => \N__48413\,
            DOUT => \N__48412\,
            PACKAGEPIN => \T23_wire\
        );

    \T23_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48414\,
            PADOUT => \N__48413\,
            PADIN => \N__48412\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__36545\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48405\,
            DIN => \N__48404\,
            DOUT => \N__48403\,
            PACKAGEPIN => pwm_output_wire
        );

    \pwm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48405\,
            PADOUT => \N__48404\,
            PADIN => \N__48403\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__26735\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48396\,
            DIN => \N__48395\,
            DOUT => \N__48394\,
            PACKAGEPIN => il_max_comp1_wire
        );

    \il_max_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48396\,
            PADOUT => \N__48395\,
            PADIN => \N__48394\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s2_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48387\,
            DIN => \N__48386\,
            DOUT => \N__48385\,
            PACKAGEPIN => s2_phy_wire
        );

    \s2_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48387\,
            PADOUT => \N__48386\,
            PADIN => \N__48385\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__34814\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T12_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48378\,
            DIN => \N__48377\,
            DOUT => \N__48376\,
            PACKAGEPIN => \T12_wire\
        );

    \T12_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48378\,
            PADOUT => \N__48377\,
            PADIN => \N__48376\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__36749\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48369\,
            DIN => \N__48368\,
            DOUT => \N__48367\,
            PACKAGEPIN => il_min_comp2_wire
        );

    \il_min_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48369\,
            PADOUT => \N__48368\,
            PADIN => \N__48367\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s1_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48360\,
            DIN => \N__48359\,
            DOUT => \N__48358\,
            PACKAGEPIN => s1_phy_wire
        );

    \s1_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48360\,
            PADOUT => \N__48359\,
            PADIN => \N__48358\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__34871\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s4_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48351\,
            DIN => \N__48350\,
            DOUT => \N__48349\,
            PACKAGEPIN => s4_phy_wire
        );

    \s4_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48351\,
            PADOUT => \N__48350\,
            PADIN => \N__48349\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__32978\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48342\,
            DIN => \N__48341\,
            DOUT => \N__48340\,
            PACKAGEPIN => il_min_comp1_wire
        );

    \il_min_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48342\,
            PADOUT => \N__48341\,
            PADIN => \N__48340\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s3_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48333\,
            DIN => \N__48332\,
            DOUT => \N__48331\,
            PACKAGEPIN => s3_phy_wire
        );

    \s3_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48333\,
            PADOUT => \N__48332\,
            PADIN => \N__48331\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__26714\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T45_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48324\,
            DIN => \N__48323\,
            DOUT => \N__48322\,
            PACKAGEPIN => \T45_wire\
        );

    \T45_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48324\,
            PADOUT => \N__48323\,
            PADIN => \N__48322\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__36728\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_hc_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48315\,
            DIN => \N__48314\,
            DOUT => \N__48313\,
            PACKAGEPIN => delay_hc_input_wire
        );

    \delay_hc_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48315\,
            PADOUT => \N__48314\,
            PADIN => \N__48313\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_hc_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_tr_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48306\,
            DIN => \N__48305\,
            DOUT => \N__48304\,
            PACKAGEPIN => delay_tr_input_wire
        );

    \delay_tr_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48306\,
            PADOUT => \N__48305\,
            PADIN => \N__48304\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_tr_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__11505\ : InMux
    port map (
            O => \N__48287\,
            I => \N__48281\
        );

    \I__11504\ : InMux
    port map (
            O => \N__48286\,
            I => \N__48278\
        );

    \I__11503\ : InMux
    port map (
            O => \N__48285\,
            I => \N__48275\
        );

    \I__11502\ : InMux
    port map (
            O => \N__48284\,
            I => \N__48272\
        );

    \I__11501\ : LocalMux
    port map (
            O => \N__48281\,
            I => \N__48269\
        );

    \I__11500\ : LocalMux
    port map (
            O => \N__48278\,
            I => \N__48266\
        );

    \I__11499\ : LocalMux
    port map (
            O => \N__48275\,
            I => \N__48263\
        );

    \I__11498\ : LocalMux
    port map (
            O => \N__48272\,
            I => \N__48260\
        );

    \I__11497\ : Span4Mux_v
    port map (
            O => \N__48269\,
            I => \N__48257\
        );

    \I__11496\ : Span4Mux_h
    port map (
            O => \N__48266\,
            I => \N__48254\
        );

    \I__11495\ : Span4Mux_h
    port map (
            O => \N__48263\,
            I => \N__48251\
        );

    \I__11494\ : Span4Mux_h
    port map (
            O => \N__48260\,
            I => \N__48248\
        );

    \I__11493\ : Span4Mux_h
    port map (
            O => \N__48257\,
            I => \N__48245\
        );

    \I__11492\ : Span4Mux_h
    port map (
            O => \N__48254\,
            I => \N__48242\
        );

    \I__11491\ : Span4Mux_h
    port map (
            O => \N__48251\,
            I => \N__48239\
        );

    \I__11490\ : Span4Mux_v
    port map (
            O => \N__48248\,
            I => \N__48236\
        );

    \I__11489\ : Odrv4
    port map (
            O => \N__48245\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__11488\ : Odrv4
    port map (
            O => \N__48242\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__11487\ : Odrv4
    port map (
            O => \N__48239\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__11486\ : Odrv4
    port map (
            O => \N__48236\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__11485\ : InMux
    port map (
            O => \N__48227\,
            I => \N__48223\
        );

    \I__11484\ : InMux
    port map (
            O => \N__48226\,
            I => \N__48219\
        );

    \I__11483\ : LocalMux
    port map (
            O => \N__48223\,
            I => \N__48216\
        );

    \I__11482\ : InMux
    port map (
            O => \N__48222\,
            I => \N__48213\
        );

    \I__11481\ : LocalMux
    port map (
            O => \N__48219\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27\
        );

    \I__11480\ : Odrv4
    port map (
            O => \N__48216\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27\
        );

    \I__11479\ : LocalMux
    port map (
            O => \N__48213\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27\
        );

    \I__11478\ : CascadeMux
    port map (
            O => \N__48206\,
            I => \N__48190\
        );

    \I__11477\ : CascadeMux
    port map (
            O => \N__48205\,
            I => \N__48173\
        );

    \I__11476\ : CascadeMux
    port map (
            O => \N__48204\,
            I => \N__48170\
        );

    \I__11475\ : InMux
    port map (
            O => \N__48203\,
            I => \N__48160\
        );

    \I__11474\ : InMux
    port map (
            O => \N__48202\,
            I => \N__48160\
        );

    \I__11473\ : InMux
    port map (
            O => \N__48201\,
            I => \N__48160\
        );

    \I__11472\ : InMux
    port map (
            O => \N__48200\,
            I => \N__48160\
        );

    \I__11471\ : InMux
    port map (
            O => \N__48199\,
            I => \N__48155\
        );

    \I__11470\ : InMux
    port map (
            O => \N__48198\,
            I => \N__48155\
        );

    \I__11469\ : InMux
    port map (
            O => \N__48197\,
            I => \N__48133\
        );

    \I__11468\ : InMux
    port map (
            O => \N__48196\,
            I => \N__48133\
        );

    \I__11467\ : InMux
    port map (
            O => \N__48195\,
            I => \N__48133\
        );

    \I__11466\ : InMux
    port map (
            O => \N__48194\,
            I => \N__48133\
        );

    \I__11465\ : InMux
    port map (
            O => \N__48193\,
            I => \N__48133\
        );

    \I__11464\ : InMux
    port map (
            O => \N__48190\,
            I => \N__48118\
        );

    \I__11463\ : InMux
    port map (
            O => \N__48189\,
            I => \N__48118\
        );

    \I__11462\ : InMux
    port map (
            O => \N__48188\,
            I => \N__48118\
        );

    \I__11461\ : InMux
    port map (
            O => \N__48187\,
            I => \N__48118\
        );

    \I__11460\ : InMux
    port map (
            O => \N__48186\,
            I => \N__48118\
        );

    \I__11459\ : InMux
    port map (
            O => \N__48185\,
            I => \N__48105\
        );

    \I__11458\ : InMux
    port map (
            O => \N__48184\,
            I => \N__48105\
        );

    \I__11457\ : InMux
    port map (
            O => \N__48183\,
            I => \N__48105\
        );

    \I__11456\ : InMux
    port map (
            O => \N__48182\,
            I => \N__48105\
        );

    \I__11455\ : InMux
    port map (
            O => \N__48181\,
            I => \N__48105\
        );

    \I__11454\ : InMux
    port map (
            O => \N__48180\,
            I => \N__48102\
        );

    \I__11453\ : CascadeMux
    port map (
            O => \N__48179\,
            I => \N__48092\
        );

    \I__11452\ : InMux
    port map (
            O => \N__48178\,
            I => \N__48080\
        );

    \I__11451\ : InMux
    port map (
            O => \N__48177\,
            I => \N__48080\
        );

    \I__11450\ : InMux
    port map (
            O => \N__48176\,
            I => \N__48080\
        );

    \I__11449\ : InMux
    port map (
            O => \N__48173\,
            I => \N__48073\
        );

    \I__11448\ : InMux
    port map (
            O => \N__48170\,
            I => \N__48073\
        );

    \I__11447\ : InMux
    port map (
            O => \N__48169\,
            I => \N__48073\
        );

    \I__11446\ : LocalMux
    port map (
            O => \N__48160\,
            I => \N__48068\
        );

    \I__11445\ : LocalMux
    port map (
            O => \N__48155\,
            I => \N__48068\
        );

    \I__11444\ : InMux
    port map (
            O => \N__48154\,
            I => \N__48063\
        );

    \I__11443\ : InMux
    port map (
            O => \N__48153\,
            I => \N__48063\
        );

    \I__11442\ : InMux
    port map (
            O => \N__48152\,
            I => \N__48060\
        );

    \I__11441\ : InMux
    port map (
            O => \N__48151\,
            I => \N__48057\
        );

    \I__11440\ : InMux
    port map (
            O => \N__48150\,
            I => \N__48052\
        );

    \I__11439\ : InMux
    port map (
            O => \N__48149\,
            I => \N__48052\
        );

    \I__11438\ : InMux
    port map (
            O => \N__48148\,
            I => \N__48042\
        );

    \I__11437\ : InMux
    port map (
            O => \N__48147\,
            I => \N__48042\
        );

    \I__11436\ : InMux
    port map (
            O => \N__48146\,
            I => \N__48042\
        );

    \I__11435\ : InMux
    port map (
            O => \N__48145\,
            I => \N__48042\
        );

    \I__11434\ : InMux
    port map (
            O => \N__48144\,
            I => \N__48039\
        );

    \I__11433\ : LocalMux
    port map (
            O => \N__48133\,
            I => \N__48036\
        );

    \I__11432\ : InMux
    port map (
            O => \N__48132\,
            I => \N__48027\
        );

    \I__11431\ : InMux
    port map (
            O => \N__48131\,
            I => \N__48027\
        );

    \I__11430\ : InMux
    port map (
            O => \N__48130\,
            I => \N__48027\
        );

    \I__11429\ : InMux
    port map (
            O => \N__48129\,
            I => \N__48027\
        );

    \I__11428\ : LocalMux
    port map (
            O => \N__48118\,
            I => \N__48016\
        );

    \I__11427\ : InMux
    port map (
            O => \N__48117\,
            I => \N__48011\
        );

    \I__11426\ : InMux
    port map (
            O => \N__48116\,
            I => \N__48011\
        );

    \I__11425\ : LocalMux
    port map (
            O => \N__48105\,
            I => \N__47992\
        );

    \I__11424\ : LocalMux
    port map (
            O => \N__48102\,
            I => \N__47989\
        );

    \I__11423\ : InMux
    port map (
            O => \N__48101\,
            I => \N__47971\
        );

    \I__11422\ : InMux
    port map (
            O => \N__48100\,
            I => \N__47971\
        );

    \I__11421\ : InMux
    port map (
            O => \N__48099\,
            I => \N__47971\
        );

    \I__11420\ : InMux
    port map (
            O => \N__48098\,
            I => \N__47971\
        );

    \I__11419\ : InMux
    port map (
            O => \N__48097\,
            I => \N__47960\
        );

    \I__11418\ : InMux
    port map (
            O => \N__48096\,
            I => \N__47960\
        );

    \I__11417\ : InMux
    port map (
            O => \N__48095\,
            I => \N__47960\
        );

    \I__11416\ : InMux
    port map (
            O => \N__48092\,
            I => \N__47960\
        );

    \I__11415\ : InMux
    port map (
            O => \N__48091\,
            I => \N__47960\
        );

    \I__11414\ : InMux
    port map (
            O => \N__48090\,
            I => \N__47951\
        );

    \I__11413\ : InMux
    port map (
            O => \N__48089\,
            I => \N__47951\
        );

    \I__11412\ : InMux
    port map (
            O => \N__48088\,
            I => \N__47951\
        );

    \I__11411\ : InMux
    port map (
            O => \N__48087\,
            I => \N__47951\
        );

    \I__11410\ : LocalMux
    port map (
            O => \N__48080\,
            I => \N__47936\
        );

    \I__11409\ : LocalMux
    port map (
            O => \N__48073\,
            I => \N__47936\
        );

    \I__11408\ : Span4Mux_v
    port map (
            O => \N__48068\,
            I => \N__47936\
        );

    \I__11407\ : LocalMux
    port map (
            O => \N__48063\,
            I => \N__47936\
        );

    \I__11406\ : LocalMux
    port map (
            O => \N__48060\,
            I => \N__47936\
        );

    \I__11405\ : LocalMux
    port map (
            O => \N__48057\,
            I => \N__47936\
        );

    \I__11404\ : LocalMux
    port map (
            O => \N__48052\,
            I => \N__47936\
        );

    \I__11403\ : InMux
    port map (
            O => \N__48051\,
            I => \N__47933\
        );

    \I__11402\ : LocalMux
    port map (
            O => \N__48042\,
            I => \N__47928\
        );

    \I__11401\ : LocalMux
    port map (
            O => \N__48039\,
            I => \N__47928\
        );

    \I__11400\ : Span4Mux_v
    port map (
            O => \N__48036\,
            I => \N__47925\
        );

    \I__11399\ : LocalMux
    port map (
            O => \N__48027\,
            I => \N__47922\
        );

    \I__11398\ : InMux
    port map (
            O => \N__48026\,
            I => \N__47917\
        );

    \I__11397\ : InMux
    port map (
            O => \N__48025\,
            I => \N__47917\
        );

    \I__11396\ : InMux
    port map (
            O => \N__48024\,
            I => \N__47910\
        );

    \I__11395\ : InMux
    port map (
            O => \N__48023\,
            I => \N__47910\
        );

    \I__11394\ : InMux
    port map (
            O => \N__48022\,
            I => \N__47910\
        );

    \I__11393\ : InMux
    port map (
            O => \N__48021\,
            I => \N__47903\
        );

    \I__11392\ : InMux
    port map (
            O => \N__48020\,
            I => \N__47903\
        );

    \I__11391\ : InMux
    port map (
            O => \N__48019\,
            I => \N__47903\
        );

    \I__11390\ : Span4Mux_v
    port map (
            O => \N__48016\,
            I => \N__47898\
        );

    \I__11389\ : LocalMux
    port map (
            O => \N__48011\,
            I => \N__47898\
        );

    \I__11388\ : InMux
    port map (
            O => \N__48010\,
            I => \N__47895\
        );

    \I__11387\ : InMux
    port map (
            O => \N__48009\,
            I => \N__47886\
        );

    \I__11386\ : InMux
    port map (
            O => \N__48008\,
            I => \N__47886\
        );

    \I__11385\ : InMux
    port map (
            O => \N__48007\,
            I => \N__47886\
        );

    \I__11384\ : InMux
    port map (
            O => \N__48006\,
            I => \N__47886\
        );

    \I__11383\ : InMux
    port map (
            O => \N__48005\,
            I => \N__47879\
        );

    \I__11382\ : InMux
    port map (
            O => \N__48004\,
            I => \N__47879\
        );

    \I__11381\ : InMux
    port map (
            O => \N__48003\,
            I => \N__47879\
        );

    \I__11380\ : InMux
    port map (
            O => \N__48002\,
            I => \N__47870\
        );

    \I__11379\ : InMux
    port map (
            O => \N__48001\,
            I => \N__47870\
        );

    \I__11378\ : InMux
    port map (
            O => \N__48000\,
            I => \N__47870\
        );

    \I__11377\ : InMux
    port map (
            O => \N__47999\,
            I => \N__47870\
        );

    \I__11376\ : InMux
    port map (
            O => \N__47998\,
            I => \N__47861\
        );

    \I__11375\ : InMux
    port map (
            O => \N__47997\,
            I => \N__47861\
        );

    \I__11374\ : InMux
    port map (
            O => \N__47996\,
            I => \N__47861\
        );

    \I__11373\ : InMux
    port map (
            O => \N__47995\,
            I => \N__47861\
        );

    \I__11372\ : Span4Mux_h
    port map (
            O => \N__47992\,
            I => \N__47856\
        );

    \I__11371\ : Span4Mux_v
    port map (
            O => \N__47989\,
            I => \N__47856\
        );

    \I__11370\ : InMux
    port map (
            O => \N__47988\,
            I => \N__47853\
        );

    \I__11369\ : InMux
    port map (
            O => \N__47987\,
            I => \N__47848\
        );

    \I__11368\ : InMux
    port map (
            O => \N__47986\,
            I => \N__47848\
        );

    \I__11367\ : InMux
    port map (
            O => \N__47985\,
            I => \N__47839\
        );

    \I__11366\ : InMux
    port map (
            O => \N__47984\,
            I => \N__47839\
        );

    \I__11365\ : InMux
    port map (
            O => \N__47983\,
            I => \N__47839\
        );

    \I__11364\ : InMux
    port map (
            O => \N__47982\,
            I => \N__47839\
        );

    \I__11363\ : InMux
    port map (
            O => \N__47981\,
            I => \N__47834\
        );

    \I__11362\ : InMux
    port map (
            O => \N__47980\,
            I => \N__47834\
        );

    \I__11361\ : LocalMux
    port map (
            O => \N__47971\,
            I => \N__47827\
        );

    \I__11360\ : LocalMux
    port map (
            O => \N__47960\,
            I => \N__47827\
        );

    \I__11359\ : LocalMux
    port map (
            O => \N__47951\,
            I => \N__47827\
        );

    \I__11358\ : Span4Mux_v
    port map (
            O => \N__47936\,
            I => \N__47824\
        );

    \I__11357\ : LocalMux
    port map (
            O => \N__47933\,
            I => \N__47813\
        );

    \I__11356\ : Span4Mux_h
    port map (
            O => \N__47928\,
            I => \N__47813\
        );

    \I__11355\ : Span4Mux_h
    port map (
            O => \N__47925\,
            I => \N__47813\
        );

    \I__11354\ : Span4Mux_v
    port map (
            O => \N__47922\,
            I => \N__47813\
        );

    \I__11353\ : LocalMux
    port map (
            O => \N__47917\,
            I => \N__47813\
        );

    \I__11352\ : LocalMux
    port map (
            O => \N__47910\,
            I => \N__47806\
        );

    \I__11351\ : LocalMux
    port map (
            O => \N__47903\,
            I => \N__47806\
        );

    \I__11350\ : Span4Mux_h
    port map (
            O => \N__47898\,
            I => \N__47806\
        );

    \I__11349\ : LocalMux
    port map (
            O => \N__47895\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11348\ : LocalMux
    port map (
            O => \N__47886\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11347\ : LocalMux
    port map (
            O => \N__47879\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11346\ : LocalMux
    port map (
            O => \N__47870\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11345\ : LocalMux
    port map (
            O => \N__47861\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11344\ : Odrv4
    port map (
            O => \N__47856\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11343\ : LocalMux
    port map (
            O => \N__47853\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11342\ : LocalMux
    port map (
            O => \N__47848\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11341\ : LocalMux
    port map (
            O => \N__47839\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11340\ : LocalMux
    port map (
            O => \N__47834\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11339\ : Odrv4
    port map (
            O => \N__47827\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11338\ : Odrv4
    port map (
            O => \N__47824\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11337\ : Odrv4
    port map (
            O => \N__47813\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11336\ : Odrv4
    port map (
            O => \N__47806\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11335\ : CascadeMux
    port map (
            O => \N__47777\,
            I => \N__47772\
        );

    \I__11334\ : InMux
    port map (
            O => \N__47776\,
            I => \N__47769\
        );

    \I__11333\ : InMux
    port map (
            O => \N__47775\,
            I => \N__47766\
        );

    \I__11332\ : InMux
    port map (
            O => \N__47772\,
            I => \N__47763\
        );

    \I__11331\ : LocalMux
    port map (
            O => \N__47769\,
            I => \N__47759\
        );

    \I__11330\ : LocalMux
    port map (
            O => \N__47766\,
            I => \N__47756\
        );

    \I__11329\ : LocalMux
    port map (
            O => \N__47763\,
            I => \N__47753\
        );

    \I__11328\ : InMux
    port map (
            O => \N__47762\,
            I => \N__47750\
        );

    \I__11327\ : Span4Mux_h
    port map (
            O => \N__47759\,
            I => \N__47747\
        );

    \I__11326\ : Span4Mux_h
    port map (
            O => \N__47756\,
            I => \N__47744\
        );

    \I__11325\ : Span4Mux_h
    port map (
            O => \N__47753\,
            I => \N__47741\
        );

    \I__11324\ : LocalMux
    port map (
            O => \N__47750\,
            I => \N__47738\
        );

    \I__11323\ : Span4Mux_h
    port map (
            O => \N__47747\,
            I => \N__47735\
        );

    \I__11322\ : Span4Mux_h
    port map (
            O => \N__47744\,
            I => \N__47730\
        );

    \I__11321\ : Span4Mux_v
    port map (
            O => \N__47741\,
            I => \N__47730\
        );

    \I__11320\ : Odrv12
    port map (
            O => \N__47738\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__11319\ : Odrv4
    port map (
            O => \N__47735\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__11318\ : Odrv4
    port map (
            O => \N__47730\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__11317\ : InMux
    port map (
            O => \N__47723\,
            I => \N__47719\
        );

    \I__11316\ : InMux
    port map (
            O => \N__47722\,
            I => \N__47715\
        );

    \I__11315\ : LocalMux
    port map (
            O => \N__47719\,
            I => \N__47712\
        );

    \I__11314\ : InMux
    port map (
            O => \N__47718\,
            I => \N__47709\
        );

    \I__11313\ : LocalMux
    port map (
            O => \N__47715\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25\
        );

    \I__11312\ : Odrv4
    port map (
            O => \N__47712\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25\
        );

    \I__11311\ : LocalMux
    port map (
            O => \N__47709\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25\
        );

    \I__11310\ : ClkMux
    port map (
            O => \N__47702\,
            I => \N__47240\
        );

    \I__11309\ : ClkMux
    port map (
            O => \N__47701\,
            I => \N__47240\
        );

    \I__11308\ : ClkMux
    port map (
            O => \N__47700\,
            I => \N__47240\
        );

    \I__11307\ : ClkMux
    port map (
            O => \N__47699\,
            I => \N__47240\
        );

    \I__11306\ : ClkMux
    port map (
            O => \N__47698\,
            I => \N__47240\
        );

    \I__11305\ : ClkMux
    port map (
            O => \N__47697\,
            I => \N__47240\
        );

    \I__11304\ : ClkMux
    port map (
            O => \N__47696\,
            I => \N__47240\
        );

    \I__11303\ : ClkMux
    port map (
            O => \N__47695\,
            I => \N__47240\
        );

    \I__11302\ : ClkMux
    port map (
            O => \N__47694\,
            I => \N__47240\
        );

    \I__11301\ : ClkMux
    port map (
            O => \N__47693\,
            I => \N__47240\
        );

    \I__11300\ : ClkMux
    port map (
            O => \N__47692\,
            I => \N__47240\
        );

    \I__11299\ : ClkMux
    port map (
            O => \N__47691\,
            I => \N__47240\
        );

    \I__11298\ : ClkMux
    port map (
            O => \N__47690\,
            I => \N__47240\
        );

    \I__11297\ : ClkMux
    port map (
            O => \N__47689\,
            I => \N__47240\
        );

    \I__11296\ : ClkMux
    port map (
            O => \N__47688\,
            I => \N__47240\
        );

    \I__11295\ : ClkMux
    port map (
            O => \N__47687\,
            I => \N__47240\
        );

    \I__11294\ : ClkMux
    port map (
            O => \N__47686\,
            I => \N__47240\
        );

    \I__11293\ : ClkMux
    port map (
            O => \N__47685\,
            I => \N__47240\
        );

    \I__11292\ : ClkMux
    port map (
            O => \N__47684\,
            I => \N__47240\
        );

    \I__11291\ : ClkMux
    port map (
            O => \N__47683\,
            I => \N__47240\
        );

    \I__11290\ : ClkMux
    port map (
            O => \N__47682\,
            I => \N__47240\
        );

    \I__11289\ : ClkMux
    port map (
            O => \N__47681\,
            I => \N__47240\
        );

    \I__11288\ : ClkMux
    port map (
            O => \N__47680\,
            I => \N__47240\
        );

    \I__11287\ : ClkMux
    port map (
            O => \N__47679\,
            I => \N__47240\
        );

    \I__11286\ : ClkMux
    port map (
            O => \N__47678\,
            I => \N__47240\
        );

    \I__11285\ : ClkMux
    port map (
            O => \N__47677\,
            I => \N__47240\
        );

    \I__11284\ : ClkMux
    port map (
            O => \N__47676\,
            I => \N__47240\
        );

    \I__11283\ : ClkMux
    port map (
            O => \N__47675\,
            I => \N__47240\
        );

    \I__11282\ : ClkMux
    port map (
            O => \N__47674\,
            I => \N__47240\
        );

    \I__11281\ : ClkMux
    port map (
            O => \N__47673\,
            I => \N__47240\
        );

    \I__11280\ : ClkMux
    port map (
            O => \N__47672\,
            I => \N__47240\
        );

    \I__11279\ : ClkMux
    port map (
            O => \N__47671\,
            I => \N__47240\
        );

    \I__11278\ : ClkMux
    port map (
            O => \N__47670\,
            I => \N__47240\
        );

    \I__11277\ : ClkMux
    port map (
            O => \N__47669\,
            I => \N__47240\
        );

    \I__11276\ : ClkMux
    port map (
            O => \N__47668\,
            I => \N__47240\
        );

    \I__11275\ : ClkMux
    port map (
            O => \N__47667\,
            I => \N__47240\
        );

    \I__11274\ : ClkMux
    port map (
            O => \N__47666\,
            I => \N__47240\
        );

    \I__11273\ : ClkMux
    port map (
            O => \N__47665\,
            I => \N__47240\
        );

    \I__11272\ : ClkMux
    port map (
            O => \N__47664\,
            I => \N__47240\
        );

    \I__11271\ : ClkMux
    port map (
            O => \N__47663\,
            I => \N__47240\
        );

    \I__11270\ : ClkMux
    port map (
            O => \N__47662\,
            I => \N__47240\
        );

    \I__11269\ : ClkMux
    port map (
            O => \N__47661\,
            I => \N__47240\
        );

    \I__11268\ : ClkMux
    port map (
            O => \N__47660\,
            I => \N__47240\
        );

    \I__11267\ : ClkMux
    port map (
            O => \N__47659\,
            I => \N__47240\
        );

    \I__11266\ : ClkMux
    port map (
            O => \N__47658\,
            I => \N__47240\
        );

    \I__11265\ : ClkMux
    port map (
            O => \N__47657\,
            I => \N__47240\
        );

    \I__11264\ : ClkMux
    port map (
            O => \N__47656\,
            I => \N__47240\
        );

    \I__11263\ : ClkMux
    port map (
            O => \N__47655\,
            I => \N__47240\
        );

    \I__11262\ : ClkMux
    port map (
            O => \N__47654\,
            I => \N__47240\
        );

    \I__11261\ : ClkMux
    port map (
            O => \N__47653\,
            I => \N__47240\
        );

    \I__11260\ : ClkMux
    port map (
            O => \N__47652\,
            I => \N__47240\
        );

    \I__11259\ : ClkMux
    port map (
            O => \N__47651\,
            I => \N__47240\
        );

    \I__11258\ : ClkMux
    port map (
            O => \N__47650\,
            I => \N__47240\
        );

    \I__11257\ : ClkMux
    port map (
            O => \N__47649\,
            I => \N__47240\
        );

    \I__11256\ : ClkMux
    port map (
            O => \N__47648\,
            I => \N__47240\
        );

    \I__11255\ : ClkMux
    port map (
            O => \N__47647\,
            I => \N__47240\
        );

    \I__11254\ : ClkMux
    port map (
            O => \N__47646\,
            I => \N__47240\
        );

    \I__11253\ : ClkMux
    port map (
            O => \N__47645\,
            I => \N__47240\
        );

    \I__11252\ : ClkMux
    port map (
            O => \N__47644\,
            I => \N__47240\
        );

    \I__11251\ : ClkMux
    port map (
            O => \N__47643\,
            I => \N__47240\
        );

    \I__11250\ : ClkMux
    port map (
            O => \N__47642\,
            I => \N__47240\
        );

    \I__11249\ : ClkMux
    port map (
            O => \N__47641\,
            I => \N__47240\
        );

    \I__11248\ : ClkMux
    port map (
            O => \N__47640\,
            I => \N__47240\
        );

    \I__11247\ : ClkMux
    port map (
            O => \N__47639\,
            I => \N__47240\
        );

    \I__11246\ : ClkMux
    port map (
            O => \N__47638\,
            I => \N__47240\
        );

    \I__11245\ : ClkMux
    port map (
            O => \N__47637\,
            I => \N__47240\
        );

    \I__11244\ : ClkMux
    port map (
            O => \N__47636\,
            I => \N__47240\
        );

    \I__11243\ : ClkMux
    port map (
            O => \N__47635\,
            I => \N__47240\
        );

    \I__11242\ : ClkMux
    port map (
            O => \N__47634\,
            I => \N__47240\
        );

    \I__11241\ : ClkMux
    port map (
            O => \N__47633\,
            I => \N__47240\
        );

    \I__11240\ : ClkMux
    port map (
            O => \N__47632\,
            I => \N__47240\
        );

    \I__11239\ : ClkMux
    port map (
            O => \N__47631\,
            I => \N__47240\
        );

    \I__11238\ : ClkMux
    port map (
            O => \N__47630\,
            I => \N__47240\
        );

    \I__11237\ : ClkMux
    port map (
            O => \N__47629\,
            I => \N__47240\
        );

    \I__11236\ : ClkMux
    port map (
            O => \N__47628\,
            I => \N__47240\
        );

    \I__11235\ : ClkMux
    port map (
            O => \N__47627\,
            I => \N__47240\
        );

    \I__11234\ : ClkMux
    port map (
            O => \N__47626\,
            I => \N__47240\
        );

    \I__11233\ : ClkMux
    port map (
            O => \N__47625\,
            I => \N__47240\
        );

    \I__11232\ : ClkMux
    port map (
            O => \N__47624\,
            I => \N__47240\
        );

    \I__11231\ : ClkMux
    port map (
            O => \N__47623\,
            I => \N__47240\
        );

    \I__11230\ : ClkMux
    port map (
            O => \N__47622\,
            I => \N__47240\
        );

    \I__11229\ : ClkMux
    port map (
            O => \N__47621\,
            I => \N__47240\
        );

    \I__11228\ : ClkMux
    port map (
            O => \N__47620\,
            I => \N__47240\
        );

    \I__11227\ : ClkMux
    port map (
            O => \N__47619\,
            I => \N__47240\
        );

    \I__11226\ : ClkMux
    port map (
            O => \N__47618\,
            I => \N__47240\
        );

    \I__11225\ : ClkMux
    port map (
            O => \N__47617\,
            I => \N__47240\
        );

    \I__11224\ : ClkMux
    port map (
            O => \N__47616\,
            I => \N__47240\
        );

    \I__11223\ : ClkMux
    port map (
            O => \N__47615\,
            I => \N__47240\
        );

    \I__11222\ : ClkMux
    port map (
            O => \N__47614\,
            I => \N__47240\
        );

    \I__11221\ : ClkMux
    port map (
            O => \N__47613\,
            I => \N__47240\
        );

    \I__11220\ : ClkMux
    port map (
            O => \N__47612\,
            I => \N__47240\
        );

    \I__11219\ : ClkMux
    port map (
            O => \N__47611\,
            I => \N__47240\
        );

    \I__11218\ : ClkMux
    port map (
            O => \N__47610\,
            I => \N__47240\
        );

    \I__11217\ : ClkMux
    port map (
            O => \N__47609\,
            I => \N__47240\
        );

    \I__11216\ : ClkMux
    port map (
            O => \N__47608\,
            I => \N__47240\
        );

    \I__11215\ : ClkMux
    port map (
            O => \N__47607\,
            I => \N__47240\
        );

    \I__11214\ : ClkMux
    port map (
            O => \N__47606\,
            I => \N__47240\
        );

    \I__11213\ : ClkMux
    port map (
            O => \N__47605\,
            I => \N__47240\
        );

    \I__11212\ : ClkMux
    port map (
            O => \N__47604\,
            I => \N__47240\
        );

    \I__11211\ : ClkMux
    port map (
            O => \N__47603\,
            I => \N__47240\
        );

    \I__11210\ : ClkMux
    port map (
            O => \N__47602\,
            I => \N__47240\
        );

    \I__11209\ : ClkMux
    port map (
            O => \N__47601\,
            I => \N__47240\
        );

    \I__11208\ : ClkMux
    port map (
            O => \N__47600\,
            I => \N__47240\
        );

    \I__11207\ : ClkMux
    port map (
            O => \N__47599\,
            I => \N__47240\
        );

    \I__11206\ : ClkMux
    port map (
            O => \N__47598\,
            I => \N__47240\
        );

    \I__11205\ : ClkMux
    port map (
            O => \N__47597\,
            I => \N__47240\
        );

    \I__11204\ : ClkMux
    port map (
            O => \N__47596\,
            I => \N__47240\
        );

    \I__11203\ : ClkMux
    port map (
            O => \N__47595\,
            I => \N__47240\
        );

    \I__11202\ : ClkMux
    port map (
            O => \N__47594\,
            I => \N__47240\
        );

    \I__11201\ : ClkMux
    port map (
            O => \N__47593\,
            I => \N__47240\
        );

    \I__11200\ : ClkMux
    port map (
            O => \N__47592\,
            I => \N__47240\
        );

    \I__11199\ : ClkMux
    port map (
            O => \N__47591\,
            I => \N__47240\
        );

    \I__11198\ : ClkMux
    port map (
            O => \N__47590\,
            I => \N__47240\
        );

    \I__11197\ : ClkMux
    port map (
            O => \N__47589\,
            I => \N__47240\
        );

    \I__11196\ : ClkMux
    port map (
            O => \N__47588\,
            I => \N__47240\
        );

    \I__11195\ : ClkMux
    port map (
            O => \N__47587\,
            I => \N__47240\
        );

    \I__11194\ : ClkMux
    port map (
            O => \N__47586\,
            I => \N__47240\
        );

    \I__11193\ : ClkMux
    port map (
            O => \N__47585\,
            I => \N__47240\
        );

    \I__11192\ : ClkMux
    port map (
            O => \N__47584\,
            I => \N__47240\
        );

    \I__11191\ : ClkMux
    port map (
            O => \N__47583\,
            I => \N__47240\
        );

    \I__11190\ : ClkMux
    port map (
            O => \N__47582\,
            I => \N__47240\
        );

    \I__11189\ : ClkMux
    port map (
            O => \N__47581\,
            I => \N__47240\
        );

    \I__11188\ : ClkMux
    port map (
            O => \N__47580\,
            I => \N__47240\
        );

    \I__11187\ : ClkMux
    port map (
            O => \N__47579\,
            I => \N__47240\
        );

    \I__11186\ : ClkMux
    port map (
            O => \N__47578\,
            I => \N__47240\
        );

    \I__11185\ : ClkMux
    port map (
            O => \N__47577\,
            I => \N__47240\
        );

    \I__11184\ : ClkMux
    port map (
            O => \N__47576\,
            I => \N__47240\
        );

    \I__11183\ : ClkMux
    port map (
            O => \N__47575\,
            I => \N__47240\
        );

    \I__11182\ : ClkMux
    port map (
            O => \N__47574\,
            I => \N__47240\
        );

    \I__11181\ : ClkMux
    port map (
            O => \N__47573\,
            I => \N__47240\
        );

    \I__11180\ : ClkMux
    port map (
            O => \N__47572\,
            I => \N__47240\
        );

    \I__11179\ : ClkMux
    port map (
            O => \N__47571\,
            I => \N__47240\
        );

    \I__11178\ : ClkMux
    port map (
            O => \N__47570\,
            I => \N__47240\
        );

    \I__11177\ : ClkMux
    port map (
            O => \N__47569\,
            I => \N__47240\
        );

    \I__11176\ : ClkMux
    port map (
            O => \N__47568\,
            I => \N__47240\
        );

    \I__11175\ : ClkMux
    port map (
            O => \N__47567\,
            I => \N__47240\
        );

    \I__11174\ : ClkMux
    port map (
            O => \N__47566\,
            I => \N__47240\
        );

    \I__11173\ : ClkMux
    port map (
            O => \N__47565\,
            I => \N__47240\
        );

    \I__11172\ : ClkMux
    port map (
            O => \N__47564\,
            I => \N__47240\
        );

    \I__11171\ : ClkMux
    port map (
            O => \N__47563\,
            I => \N__47240\
        );

    \I__11170\ : ClkMux
    port map (
            O => \N__47562\,
            I => \N__47240\
        );

    \I__11169\ : ClkMux
    port map (
            O => \N__47561\,
            I => \N__47240\
        );

    \I__11168\ : ClkMux
    port map (
            O => \N__47560\,
            I => \N__47240\
        );

    \I__11167\ : ClkMux
    port map (
            O => \N__47559\,
            I => \N__47240\
        );

    \I__11166\ : ClkMux
    port map (
            O => \N__47558\,
            I => \N__47240\
        );

    \I__11165\ : ClkMux
    port map (
            O => \N__47557\,
            I => \N__47240\
        );

    \I__11164\ : ClkMux
    port map (
            O => \N__47556\,
            I => \N__47240\
        );

    \I__11163\ : ClkMux
    port map (
            O => \N__47555\,
            I => \N__47240\
        );

    \I__11162\ : ClkMux
    port map (
            O => \N__47554\,
            I => \N__47240\
        );

    \I__11161\ : ClkMux
    port map (
            O => \N__47553\,
            I => \N__47240\
        );

    \I__11160\ : ClkMux
    port map (
            O => \N__47552\,
            I => \N__47240\
        );

    \I__11159\ : ClkMux
    port map (
            O => \N__47551\,
            I => \N__47240\
        );

    \I__11158\ : ClkMux
    port map (
            O => \N__47550\,
            I => \N__47240\
        );

    \I__11157\ : ClkMux
    port map (
            O => \N__47549\,
            I => \N__47240\
        );

    \I__11156\ : GlobalMux
    port map (
            O => \N__47240\,
            I => clk_100mhz_0
        );

    \I__11155\ : CEMux
    port map (
            O => \N__47237\,
            I => \N__47233\
        );

    \I__11154\ : CEMux
    port map (
            O => \N__47236\,
            I => \N__47230\
        );

    \I__11153\ : LocalMux
    port map (
            O => \N__47233\,
            I => \N__47224\
        );

    \I__11152\ : LocalMux
    port map (
            O => \N__47230\,
            I => \N__47224\
        );

    \I__11151\ : CEMux
    port map (
            O => \N__47229\,
            I => \N__47221\
        );

    \I__11150\ : Span4Mux_v
    port map (
            O => \N__47224\,
            I => \N__47216\
        );

    \I__11149\ : LocalMux
    port map (
            O => \N__47221\,
            I => \N__47213\
        );

    \I__11148\ : CEMux
    port map (
            O => \N__47220\,
            I => \N__47210\
        );

    \I__11147\ : CEMux
    port map (
            O => \N__47219\,
            I => \N__47205\
        );

    \I__11146\ : Span4Mux_h
    port map (
            O => \N__47216\,
            I => \N__47195\
        );

    \I__11145\ : Span4Mux_v
    port map (
            O => \N__47213\,
            I => \N__47195\
        );

    \I__11144\ : LocalMux
    port map (
            O => \N__47210\,
            I => \N__47195\
        );

    \I__11143\ : CEMux
    port map (
            O => \N__47209\,
            I => \N__47192\
        );

    \I__11142\ : CEMux
    port map (
            O => \N__47208\,
            I => \N__47185\
        );

    \I__11141\ : LocalMux
    port map (
            O => \N__47205\,
            I => \N__47182\
        );

    \I__11140\ : CEMux
    port map (
            O => \N__47204\,
            I => \N__47179\
        );

    \I__11139\ : CEMux
    port map (
            O => \N__47203\,
            I => \N__47176\
        );

    \I__11138\ : CEMux
    port map (
            O => \N__47202\,
            I => \N__47173\
        );

    \I__11137\ : Span4Mux_v
    port map (
            O => \N__47195\,
            I => \N__47166\
        );

    \I__11136\ : LocalMux
    port map (
            O => \N__47192\,
            I => \N__47166\
        );

    \I__11135\ : InMux
    port map (
            O => \N__47191\,
            I => \N__47147\
        );

    \I__11134\ : InMux
    port map (
            O => \N__47190\,
            I => \N__47140\
        );

    \I__11133\ : InMux
    port map (
            O => \N__47189\,
            I => \N__47140\
        );

    \I__11132\ : InMux
    port map (
            O => \N__47188\,
            I => \N__47140\
        );

    \I__11131\ : LocalMux
    port map (
            O => \N__47185\,
            I => \N__47137\
        );

    \I__11130\ : Span4Mux_h
    port map (
            O => \N__47182\,
            I => \N__47134\
        );

    \I__11129\ : LocalMux
    port map (
            O => \N__47179\,
            I => \N__47131\
        );

    \I__11128\ : LocalMux
    port map (
            O => \N__47176\,
            I => \N__47126\
        );

    \I__11127\ : LocalMux
    port map (
            O => \N__47173\,
            I => \N__47126\
        );

    \I__11126\ : CEMux
    port map (
            O => \N__47172\,
            I => \N__47123\
        );

    \I__11125\ : CEMux
    port map (
            O => \N__47171\,
            I => \N__47120\
        );

    \I__11124\ : Span4Mux_v
    port map (
            O => \N__47166\,
            I => \N__47110\
        );

    \I__11123\ : InMux
    port map (
            O => \N__47165\,
            I => \N__47101\
        );

    \I__11122\ : InMux
    port map (
            O => \N__47164\,
            I => \N__47101\
        );

    \I__11121\ : InMux
    port map (
            O => \N__47163\,
            I => \N__47101\
        );

    \I__11120\ : InMux
    port map (
            O => \N__47162\,
            I => \N__47101\
        );

    \I__11119\ : InMux
    port map (
            O => \N__47161\,
            I => \N__47092\
        );

    \I__11118\ : InMux
    port map (
            O => \N__47160\,
            I => \N__47092\
        );

    \I__11117\ : InMux
    port map (
            O => \N__47159\,
            I => \N__47092\
        );

    \I__11116\ : InMux
    port map (
            O => \N__47158\,
            I => \N__47092\
        );

    \I__11115\ : InMux
    port map (
            O => \N__47157\,
            I => \N__47083\
        );

    \I__11114\ : InMux
    port map (
            O => \N__47156\,
            I => \N__47083\
        );

    \I__11113\ : InMux
    port map (
            O => \N__47155\,
            I => \N__47083\
        );

    \I__11112\ : InMux
    port map (
            O => \N__47154\,
            I => \N__47083\
        );

    \I__11111\ : InMux
    port map (
            O => \N__47153\,
            I => \N__47074\
        );

    \I__11110\ : InMux
    port map (
            O => \N__47152\,
            I => \N__47074\
        );

    \I__11109\ : InMux
    port map (
            O => \N__47151\,
            I => \N__47074\
        );

    \I__11108\ : InMux
    port map (
            O => \N__47150\,
            I => \N__47074\
        );

    \I__11107\ : LocalMux
    port map (
            O => \N__47147\,
            I => \N__47071\
        );

    \I__11106\ : LocalMux
    port map (
            O => \N__47140\,
            I => \N__47062\
        );

    \I__11105\ : Span4Mux_v
    port map (
            O => \N__47137\,
            I => \N__47062\
        );

    \I__11104\ : Span4Mux_v
    port map (
            O => \N__47134\,
            I => \N__47053\
        );

    \I__11103\ : Span4Mux_v
    port map (
            O => \N__47131\,
            I => \N__47053\
        );

    \I__11102\ : Span4Mux_h
    port map (
            O => \N__47126\,
            I => \N__47053\
        );

    \I__11101\ : LocalMux
    port map (
            O => \N__47123\,
            I => \N__47053\
        );

    \I__11100\ : LocalMux
    port map (
            O => \N__47120\,
            I => \N__47050\
        );

    \I__11099\ : InMux
    port map (
            O => \N__47119\,
            I => \N__47043\
        );

    \I__11098\ : InMux
    port map (
            O => \N__47118\,
            I => \N__47043\
        );

    \I__11097\ : InMux
    port map (
            O => \N__47117\,
            I => \N__47043\
        );

    \I__11096\ : InMux
    port map (
            O => \N__47116\,
            I => \N__47034\
        );

    \I__11095\ : InMux
    port map (
            O => \N__47115\,
            I => \N__47034\
        );

    \I__11094\ : InMux
    port map (
            O => \N__47114\,
            I => \N__47034\
        );

    \I__11093\ : InMux
    port map (
            O => \N__47113\,
            I => \N__47034\
        );

    \I__11092\ : Span4Mux_v
    port map (
            O => \N__47110\,
            I => \N__47029\
        );

    \I__11091\ : LocalMux
    port map (
            O => \N__47101\,
            I => \N__47029\
        );

    \I__11090\ : LocalMux
    port map (
            O => \N__47092\,
            I => \N__47026\
        );

    \I__11089\ : LocalMux
    port map (
            O => \N__47083\,
            I => \N__47019\
        );

    \I__11088\ : LocalMux
    port map (
            O => \N__47074\,
            I => \N__47019\
        );

    \I__11087\ : Span4Mux_h
    port map (
            O => \N__47071\,
            I => \N__47019\
        );

    \I__11086\ : InMux
    port map (
            O => \N__47070\,
            I => \N__47010\
        );

    \I__11085\ : InMux
    port map (
            O => \N__47069\,
            I => \N__47010\
        );

    \I__11084\ : InMux
    port map (
            O => \N__47068\,
            I => \N__47010\
        );

    \I__11083\ : InMux
    port map (
            O => \N__47067\,
            I => \N__47010\
        );

    \I__11082\ : Span4Mux_h
    port map (
            O => \N__47062\,
            I => \N__47005\
        );

    \I__11081\ : Span4Mux_v
    port map (
            O => \N__47053\,
            I => \N__47005\
        );

    \I__11080\ : Span4Mux_v
    port map (
            O => \N__47050\,
            I => \N__46998\
        );

    \I__11079\ : LocalMux
    port map (
            O => \N__47043\,
            I => \N__46998\
        );

    \I__11078\ : LocalMux
    port map (
            O => \N__47034\,
            I => \N__46998\
        );

    \I__11077\ : Span4Mux_v
    port map (
            O => \N__47029\,
            I => \N__46993\
        );

    \I__11076\ : Span4Mux_v
    port map (
            O => \N__47026\,
            I => \N__46993\
        );

    \I__11075\ : Span4Mux_h
    port map (
            O => \N__47019\,
            I => \N__46990\
        );

    \I__11074\ : LocalMux
    port map (
            O => \N__47010\,
            I => \N__46987\
        );

    \I__11073\ : Span4Mux_h
    port map (
            O => \N__47005\,
            I => \N__46984\
        );

    \I__11072\ : Span4Mux_h
    port map (
            O => \N__46998\,
            I => \N__46981\
        );

    \I__11071\ : Span4Mux_h
    port map (
            O => \N__46993\,
            I => \N__46978\
        );

    \I__11070\ : Span4Mux_h
    port map (
            O => \N__46990\,
            I => \N__46975\
        );

    \I__11069\ : Span4Mux_h
    port map (
            O => \N__46987\,
            I => \N__46970\
        );

    \I__11068\ : Span4Mux_s2_h
    port map (
            O => \N__46984\,
            I => \N__46970\
        );

    \I__11067\ : Odrv4
    port map (
            O => \N__46981\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__11066\ : Odrv4
    port map (
            O => \N__46978\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__11065\ : Odrv4
    port map (
            O => \N__46975\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__11064\ : Odrv4
    port map (
            O => \N__46970\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__11063\ : InMux
    port map (
            O => \N__46961\,
            I => \N__46955\
        );

    \I__11062\ : InMux
    port map (
            O => \N__46960\,
            I => \N__46950\
        );

    \I__11061\ : InMux
    port map (
            O => \N__46959\,
            I => \N__46950\
        );

    \I__11060\ : InMux
    port map (
            O => \N__46958\,
            I => \N__46947\
        );

    \I__11059\ : LocalMux
    port map (
            O => \N__46955\,
            I => \N__46944\
        );

    \I__11058\ : LocalMux
    port map (
            O => \N__46950\,
            I => \N__46941\
        );

    \I__11057\ : LocalMux
    port map (
            O => \N__46947\,
            I => \N__46933\
        );

    \I__11056\ : Glb2LocalMux
    port map (
            O => \N__46944\,
            I => \N__46466\
        );

    \I__11055\ : Glb2LocalMux
    port map (
            O => \N__46941\,
            I => \N__46466\
        );

    \I__11054\ : SRMux
    port map (
            O => \N__46940\,
            I => \N__46466\
        );

    \I__11053\ : SRMux
    port map (
            O => \N__46939\,
            I => \N__46466\
        );

    \I__11052\ : SRMux
    port map (
            O => \N__46938\,
            I => \N__46466\
        );

    \I__11051\ : SRMux
    port map (
            O => \N__46937\,
            I => \N__46466\
        );

    \I__11050\ : SRMux
    port map (
            O => \N__46936\,
            I => \N__46466\
        );

    \I__11049\ : Glb2LocalMux
    port map (
            O => \N__46933\,
            I => \N__46466\
        );

    \I__11048\ : SRMux
    port map (
            O => \N__46932\,
            I => \N__46466\
        );

    \I__11047\ : SRMux
    port map (
            O => \N__46931\,
            I => \N__46466\
        );

    \I__11046\ : SRMux
    port map (
            O => \N__46930\,
            I => \N__46466\
        );

    \I__11045\ : SRMux
    port map (
            O => \N__46929\,
            I => \N__46466\
        );

    \I__11044\ : SRMux
    port map (
            O => \N__46928\,
            I => \N__46466\
        );

    \I__11043\ : SRMux
    port map (
            O => \N__46927\,
            I => \N__46466\
        );

    \I__11042\ : SRMux
    port map (
            O => \N__46926\,
            I => \N__46466\
        );

    \I__11041\ : SRMux
    port map (
            O => \N__46925\,
            I => \N__46466\
        );

    \I__11040\ : SRMux
    port map (
            O => \N__46924\,
            I => \N__46466\
        );

    \I__11039\ : SRMux
    port map (
            O => \N__46923\,
            I => \N__46466\
        );

    \I__11038\ : SRMux
    port map (
            O => \N__46922\,
            I => \N__46466\
        );

    \I__11037\ : SRMux
    port map (
            O => \N__46921\,
            I => \N__46466\
        );

    \I__11036\ : SRMux
    port map (
            O => \N__46920\,
            I => \N__46466\
        );

    \I__11035\ : SRMux
    port map (
            O => \N__46919\,
            I => \N__46466\
        );

    \I__11034\ : SRMux
    port map (
            O => \N__46918\,
            I => \N__46466\
        );

    \I__11033\ : SRMux
    port map (
            O => \N__46917\,
            I => \N__46466\
        );

    \I__11032\ : SRMux
    port map (
            O => \N__46916\,
            I => \N__46466\
        );

    \I__11031\ : SRMux
    port map (
            O => \N__46915\,
            I => \N__46466\
        );

    \I__11030\ : SRMux
    port map (
            O => \N__46914\,
            I => \N__46466\
        );

    \I__11029\ : SRMux
    port map (
            O => \N__46913\,
            I => \N__46466\
        );

    \I__11028\ : SRMux
    port map (
            O => \N__46912\,
            I => \N__46466\
        );

    \I__11027\ : SRMux
    port map (
            O => \N__46911\,
            I => \N__46466\
        );

    \I__11026\ : SRMux
    port map (
            O => \N__46910\,
            I => \N__46466\
        );

    \I__11025\ : SRMux
    port map (
            O => \N__46909\,
            I => \N__46466\
        );

    \I__11024\ : SRMux
    port map (
            O => \N__46908\,
            I => \N__46466\
        );

    \I__11023\ : SRMux
    port map (
            O => \N__46907\,
            I => \N__46466\
        );

    \I__11022\ : SRMux
    port map (
            O => \N__46906\,
            I => \N__46466\
        );

    \I__11021\ : SRMux
    port map (
            O => \N__46905\,
            I => \N__46466\
        );

    \I__11020\ : SRMux
    port map (
            O => \N__46904\,
            I => \N__46466\
        );

    \I__11019\ : SRMux
    port map (
            O => \N__46903\,
            I => \N__46466\
        );

    \I__11018\ : SRMux
    port map (
            O => \N__46902\,
            I => \N__46466\
        );

    \I__11017\ : SRMux
    port map (
            O => \N__46901\,
            I => \N__46466\
        );

    \I__11016\ : SRMux
    port map (
            O => \N__46900\,
            I => \N__46466\
        );

    \I__11015\ : SRMux
    port map (
            O => \N__46899\,
            I => \N__46466\
        );

    \I__11014\ : SRMux
    port map (
            O => \N__46898\,
            I => \N__46466\
        );

    \I__11013\ : SRMux
    port map (
            O => \N__46897\,
            I => \N__46466\
        );

    \I__11012\ : SRMux
    port map (
            O => \N__46896\,
            I => \N__46466\
        );

    \I__11011\ : SRMux
    port map (
            O => \N__46895\,
            I => \N__46466\
        );

    \I__11010\ : SRMux
    port map (
            O => \N__46894\,
            I => \N__46466\
        );

    \I__11009\ : SRMux
    port map (
            O => \N__46893\,
            I => \N__46466\
        );

    \I__11008\ : SRMux
    port map (
            O => \N__46892\,
            I => \N__46466\
        );

    \I__11007\ : SRMux
    port map (
            O => \N__46891\,
            I => \N__46466\
        );

    \I__11006\ : SRMux
    port map (
            O => \N__46890\,
            I => \N__46466\
        );

    \I__11005\ : SRMux
    port map (
            O => \N__46889\,
            I => \N__46466\
        );

    \I__11004\ : SRMux
    port map (
            O => \N__46888\,
            I => \N__46466\
        );

    \I__11003\ : SRMux
    port map (
            O => \N__46887\,
            I => \N__46466\
        );

    \I__11002\ : SRMux
    port map (
            O => \N__46886\,
            I => \N__46466\
        );

    \I__11001\ : SRMux
    port map (
            O => \N__46885\,
            I => \N__46466\
        );

    \I__11000\ : SRMux
    port map (
            O => \N__46884\,
            I => \N__46466\
        );

    \I__10999\ : SRMux
    port map (
            O => \N__46883\,
            I => \N__46466\
        );

    \I__10998\ : SRMux
    port map (
            O => \N__46882\,
            I => \N__46466\
        );

    \I__10997\ : SRMux
    port map (
            O => \N__46881\,
            I => \N__46466\
        );

    \I__10996\ : SRMux
    port map (
            O => \N__46880\,
            I => \N__46466\
        );

    \I__10995\ : SRMux
    port map (
            O => \N__46879\,
            I => \N__46466\
        );

    \I__10994\ : SRMux
    port map (
            O => \N__46878\,
            I => \N__46466\
        );

    \I__10993\ : SRMux
    port map (
            O => \N__46877\,
            I => \N__46466\
        );

    \I__10992\ : SRMux
    port map (
            O => \N__46876\,
            I => \N__46466\
        );

    \I__10991\ : SRMux
    port map (
            O => \N__46875\,
            I => \N__46466\
        );

    \I__10990\ : SRMux
    port map (
            O => \N__46874\,
            I => \N__46466\
        );

    \I__10989\ : SRMux
    port map (
            O => \N__46873\,
            I => \N__46466\
        );

    \I__10988\ : SRMux
    port map (
            O => \N__46872\,
            I => \N__46466\
        );

    \I__10987\ : SRMux
    port map (
            O => \N__46871\,
            I => \N__46466\
        );

    \I__10986\ : SRMux
    port map (
            O => \N__46870\,
            I => \N__46466\
        );

    \I__10985\ : SRMux
    port map (
            O => \N__46869\,
            I => \N__46466\
        );

    \I__10984\ : SRMux
    port map (
            O => \N__46868\,
            I => \N__46466\
        );

    \I__10983\ : SRMux
    port map (
            O => \N__46867\,
            I => \N__46466\
        );

    \I__10982\ : SRMux
    port map (
            O => \N__46866\,
            I => \N__46466\
        );

    \I__10981\ : SRMux
    port map (
            O => \N__46865\,
            I => \N__46466\
        );

    \I__10980\ : SRMux
    port map (
            O => \N__46864\,
            I => \N__46466\
        );

    \I__10979\ : SRMux
    port map (
            O => \N__46863\,
            I => \N__46466\
        );

    \I__10978\ : SRMux
    port map (
            O => \N__46862\,
            I => \N__46466\
        );

    \I__10977\ : SRMux
    port map (
            O => \N__46861\,
            I => \N__46466\
        );

    \I__10976\ : SRMux
    port map (
            O => \N__46860\,
            I => \N__46466\
        );

    \I__10975\ : SRMux
    port map (
            O => \N__46859\,
            I => \N__46466\
        );

    \I__10974\ : SRMux
    port map (
            O => \N__46858\,
            I => \N__46466\
        );

    \I__10973\ : SRMux
    port map (
            O => \N__46857\,
            I => \N__46466\
        );

    \I__10972\ : SRMux
    port map (
            O => \N__46856\,
            I => \N__46466\
        );

    \I__10971\ : SRMux
    port map (
            O => \N__46855\,
            I => \N__46466\
        );

    \I__10970\ : SRMux
    port map (
            O => \N__46854\,
            I => \N__46466\
        );

    \I__10969\ : SRMux
    port map (
            O => \N__46853\,
            I => \N__46466\
        );

    \I__10968\ : SRMux
    port map (
            O => \N__46852\,
            I => \N__46466\
        );

    \I__10967\ : SRMux
    port map (
            O => \N__46851\,
            I => \N__46466\
        );

    \I__10966\ : SRMux
    port map (
            O => \N__46850\,
            I => \N__46466\
        );

    \I__10965\ : SRMux
    port map (
            O => \N__46849\,
            I => \N__46466\
        );

    \I__10964\ : SRMux
    port map (
            O => \N__46848\,
            I => \N__46466\
        );

    \I__10963\ : SRMux
    port map (
            O => \N__46847\,
            I => \N__46466\
        );

    \I__10962\ : SRMux
    port map (
            O => \N__46846\,
            I => \N__46466\
        );

    \I__10961\ : SRMux
    port map (
            O => \N__46845\,
            I => \N__46466\
        );

    \I__10960\ : SRMux
    port map (
            O => \N__46844\,
            I => \N__46466\
        );

    \I__10959\ : SRMux
    port map (
            O => \N__46843\,
            I => \N__46466\
        );

    \I__10958\ : SRMux
    port map (
            O => \N__46842\,
            I => \N__46466\
        );

    \I__10957\ : SRMux
    port map (
            O => \N__46841\,
            I => \N__46466\
        );

    \I__10956\ : SRMux
    port map (
            O => \N__46840\,
            I => \N__46466\
        );

    \I__10955\ : SRMux
    port map (
            O => \N__46839\,
            I => \N__46466\
        );

    \I__10954\ : SRMux
    port map (
            O => \N__46838\,
            I => \N__46466\
        );

    \I__10953\ : SRMux
    port map (
            O => \N__46837\,
            I => \N__46466\
        );

    \I__10952\ : SRMux
    port map (
            O => \N__46836\,
            I => \N__46466\
        );

    \I__10951\ : SRMux
    port map (
            O => \N__46835\,
            I => \N__46466\
        );

    \I__10950\ : SRMux
    port map (
            O => \N__46834\,
            I => \N__46466\
        );

    \I__10949\ : SRMux
    port map (
            O => \N__46833\,
            I => \N__46466\
        );

    \I__10948\ : SRMux
    port map (
            O => \N__46832\,
            I => \N__46466\
        );

    \I__10947\ : SRMux
    port map (
            O => \N__46831\,
            I => \N__46466\
        );

    \I__10946\ : SRMux
    port map (
            O => \N__46830\,
            I => \N__46466\
        );

    \I__10945\ : SRMux
    port map (
            O => \N__46829\,
            I => \N__46466\
        );

    \I__10944\ : SRMux
    port map (
            O => \N__46828\,
            I => \N__46466\
        );

    \I__10943\ : SRMux
    port map (
            O => \N__46827\,
            I => \N__46466\
        );

    \I__10942\ : SRMux
    port map (
            O => \N__46826\,
            I => \N__46466\
        );

    \I__10941\ : SRMux
    port map (
            O => \N__46825\,
            I => \N__46466\
        );

    \I__10940\ : SRMux
    port map (
            O => \N__46824\,
            I => \N__46466\
        );

    \I__10939\ : SRMux
    port map (
            O => \N__46823\,
            I => \N__46466\
        );

    \I__10938\ : SRMux
    port map (
            O => \N__46822\,
            I => \N__46466\
        );

    \I__10937\ : SRMux
    port map (
            O => \N__46821\,
            I => \N__46466\
        );

    \I__10936\ : SRMux
    port map (
            O => \N__46820\,
            I => \N__46466\
        );

    \I__10935\ : SRMux
    port map (
            O => \N__46819\,
            I => \N__46466\
        );

    \I__10934\ : SRMux
    port map (
            O => \N__46818\,
            I => \N__46466\
        );

    \I__10933\ : SRMux
    port map (
            O => \N__46817\,
            I => \N__46466\
        );

    \I__10932\ : SRMux
    port map (
            O => \N__46816\,
            I => \N__46466\
        );

    \I__10931\ : SRMux
    port map (
            O => \N__46815\,
            I => \N__46466\
        );

    \I__10930\ : SRMux
    port map (
            O => \N__46814\,
            I => \N__46466\
        );

    \I__10929\ : SRMux
    port map (
            O => \N__46813\,
            I => \N__46466\
        );

    \I__10928\ : SRMux
    port map (
            O => \N__46812\,
            I => \N__46466\
        );

    \I__10927\ : SRMux
    port map (
            O => \N__46811\,
            I => \N__46466\
        );

    \I__10926\ : SRMux
    port map (
            O => \N__46810\,
            I => \N__46466\
        );

    \I__10925\ : SRMux
    port map (
            O => \N__46809\,
            I => \N__46466\
        );

    \I__10924\ : SRMux
    port map (
            O => \N__46808\,
            I => \N__46466\
        );

    \I__10923\ : SRMux
    port map (
            O => \N__46807\,
            I => \N__46466\
        );

    \I__10922\ : SRMux
    port map (
            O => \N__46806\,
            I => \N__46466\
        );

    \I__10921\ : SRMux
    port map (
            O => \N__46805\,
            I => \N__46466\
        );

    \I__10920\ : SRMux
    port map (
            O => \N__46804\,
            I => \N__46466\
        );

    \I__10919\ : SRMux
    port map (
            O => \N__46803\,
            I => \N__46466\
        );

    \I__10918\ : SRMux
    port map (
            O => \N__46802\,
            I => \N__46466\
        );

    \I__10917\ : SRMux
    port map (
            O => \N__46801\,
            I => \N__46466\
        );

    \I__10916\ : SRMux
    port map (
            O => \N__46800\,
            I => \N__46466\
        );

    \I__10915\ : SRMux
    port map (
            O => \N__46799\,
            I => \N__46466\
        );

    \I__10914\ : SRMux
    port map (
            O => \N__46798\,
            I => \N__46466\
        );

    \I__10913\ : SRMux
    port map (
            O => \N__46797\,
            I => \N__46466\
        );

    \I__10912\ : SRMux
    port map (
            O => \N__46796\,
            I => \N__46466\
        );

    \I__10911\ : SRMux
    port map (
            O => \N__46795\,
            I => \N__46466\
        );

    \I__10910\ : SRMux
    port map (
            O => \N__46794\,
            I => \N__46466\
        );

    \I__10909\ : SRMux
    port map (
            O => \N__46793\,
            I => \N__46466\
        );

    \I__10908\ : SRMux
    port map (
            O => \N__46792\,
            I => \N__46466\
        );

    \I__10907\ : SRMux
    port map (
            O => \N__46791\,
            I => \N__46466\
        );

    \I__10906\ : SRMux
    port map (
            O => \N__46790\,
            I => \N__46466\
        );

    \I__10905\ : SRMux
    port map (
            O => \N__46789\,
            I => \N__46466\
        );

    \I__10904\ : SRMux
    port map (
            O => \N__46788\,
            I => \N__46466\
        );

    \I__10903\ : SRMux
    port map (
            O => \N__46787\,
            I => \N__46466\
        );

    \I__10902\ : SRMux
    port map (
            O => \N__46786\,
            I => \N__46466\
        );

    \I__10901\ : SRMux
    port map (
            O => \N__46785\,
            I => \N__46466\
        );

    \I__10900\ : SRMux
    port map (
            O => \N__46784\,
            I => \N__46466\
        );

    \I__10899\ : SRMux
    port map (
            O => \N__46783\,
            I => \N__46466\
        );

    \I__10898\ : GlobalMux
    port map (
            O => \N__46466\,
            I => \N__46463\
        );

    \I__10897\ : gio2CtrlBuf
    port map (
            O => \N__46463\,
            I => red_c_g
        );

    \I__10896\ : CascadeMux
    port map (
            O => \N__46460\,
            I => \N__46457\
        );

    \I__10895\ : InMux
    port map (
            O => \N__46457\,
            I => \N__46454\
        );

    \I__10894\ : LocalMux
    port map (
            O => \N__46454\,
            I => \N__46451\
        );

    \I__10893\ : Span4Mux_h
    port map (
            O => \N__46451\,
            I => \N__46448\
        );

    \I__10892\ : Odrv4
    port map (
            O => \N__46448\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt24\
        );

    \I__10891\ : InMux
    port map (
            O => \N__46445\,
            I => \N__46439\
        );

    \I__10890\ : InMux
    port map (
            O => \N__46444\,
            I => \N__46439\
        );

    \I__10889\ : LocalMux
    port map (
            O => \N__46439\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_24\
        );

    \I__10888\ : InMux
    port map (
            O => \N__46436\,
            I => \N__46429\
        );

    \I__10887\ : InMux
    port map (
            O => \N__46435\,
            I => \N__46429\
        );

    \I__10886\ : InMux
    port map (
            O => \N__46434\,
            I => \N__46426\
        );

    \I__10885\ : LocalMux
    port map (
            O => \N__46429\,
            I => \N__46423\
        );

    \I__10884\ : LocalMux
    port map (
            O => \N__46426\,
            I => \N__46418\
        );

    \I__10883\ : Span4Mux_h
    port map (
            O => \N__46423\,
            I => \N__46418\
        );

    \I__10882\ : Odrv4
    port map (
            O => \N__46418\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__10881\ : CascadeMux
    port map (
            O => \N__46415\,
            I => \N__46411\
        );

    \I__10880\ : CascadeMux
    port map (
            O => \N__46414\,
            I => \N__46408\
        );

    \I__10879\ : InMux
    port map (
            O => \N__46411\,
            I => \N__46403\
        );

    \I__10878\ : InMux
    port map (
            O => \N__46408\,
            I => \N__46403\
        );

    \I__10877\ : LocalMux
    port map (
            O => \N__46403\,
            I => \N__46399\
        );

    \I__10876\ : InMux
    port map (
            O => \N__46402\,
            I => \N__46396\
        );

    \I__10875\ : Span4Mux_h
    port map (
            O => \N__46399\,
            I => \N__46393\
        );

    \I__10874\ : LocalMux
    port map (
            O => \N__46396\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__10873\ : Odrv4
    port map (
            O => \N__46393\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__10872\ : InMux
    port map (
            O => \N__46388\,
            I => \N__46382\
        );

    \I__10871\ : InMux
    port map (
            O => \N__46387\,
            I => \N__46382\
        );

    \I__10870\ : LocalMux
    port map (
            O => \N__46382\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_25\
        );

    \I__10869\ : InMux
    port map (
            O => \N__46379\,
            I => \N__46376\
        );

    \I__10868\ : LocalMux
    port map (
            O => \N__46376\,
            I => \N__46373\
        );

    \I__10867\ : Odrv12
    port map (
            O => \N__46373\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24\
        );

    \I__10866\ : CascadeMux
    port map (
            O => \N__46370\,
            I => \N__46367\
        );

    \I__10865\ : InMux
    port map (
            O => \N__46367\,
            I => \N__46362\
        );

    \I__10864\ : InMux
    port map (
            O => \N__46366\,
            I => \N__46359\
        );

    \I__10863\ : InMux
    port map (
            O => \N__46365\,
            I => \N__46356\
        );

    \I__10862\ : LocalMux
    port map (
            O => \N__46362\,
            I => \N__46351\
        );

    \I__10861\ : LocalMux
    port map (
            O => \N__46359\,
            I => \N__46351\
        );

    \I__10860\ : LocalMux
    port map (
            O => \N__46356\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__10859\ : Odrv12
    port map (
            O => \N__46351\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__10858\ : InMux
    port map (
            O => \N__46346\,
            I => \N__46342\
        );

    \I__10857\ : InMux
    port map (
            O => \N__46345\,
            I => \N__46339\
        );

    \I__10856\ : LocalMux
    port map (
            O => \N__46342\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\
        );

    \I__10855\ : LocalMux
    port map (
            O => \N__46339\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\
        );

    \I__10854\ : CascadeMux
    port map (
            O => \N__46334\,
            I => \N__46331\
        );

    \I__10853\ : InMux
    port map (
            O => \N__46331\,
            I => \N__46326\
        );

    \I__10852\ : InMux
    port map (
            O => \N__46330\,
            I => \N__46323\
        );

    \I__10851\ : InMux
    port map (
            O => \N__46329\,
            I => \N__46320\
        );

    \I__10850\ : LocalMux
    port map (
            O => \N__46326\,
            I => \N__46317\
        );

    \I__10849\ : LocalMux
    port map (
            O => \N__46323\,
            I => \N__46314\
        );

    \I__10848\ : LocalMux
    port map (
            O => \N__46320\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__10847\ : Odrv12
    port map (
            O => \N__46317\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__10846\ : Odrv4
    port map (
            O => \N__46314\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__10845\ : InMux
    port map (
            O => \N__46307\,
            I => \N__46303\
        );

    \I__10844\ : InMux
    port map (
            O => \N__46306\,
            I => \N__46300\
        );

    \I__10843\ : LocalMux
    port map (
            O => \N__46303\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\
        );

    \I__10842\ : LocalMux
    port map (
            O => \N__46300\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\
        );

    \I__10841\ : CascadeMux
    port map (
            O => \N__46295\,
            I => \N__46292\
        );

    \I__10840\ : InMux
    port map (
            O => \N__46292\,
            I => \N__46289\
        );

    \I__10839\ : LocalMux
    port map (
            O => \N__46289\,
            I => \N__46286\
        );

    \I__10838\ : Odrv12
    port map (
            O => \N__46286\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26\
        );

    \I__10837\ : InMux
    port map (
            O => \N__46283\,
            I => \N__46280\
        );

    \I__10836\ : LocalMux
    port map (
            O => \N__46280\,
            I => \N__46277\
        );

    \I__10835\ : Span4Mux_v
    port map (
            O => \N__46277\,
            I => \N__46274\
        );

    \I__10834\ : Sp12to4
    port map (
            O => \N__46274\,
            I => \N__46271\
        );

    \I__10833\ : Span12Mux_h
    port map (
            O => \N__46271\,
            I => \N__46267\
        );

    \I__10832\ : InMux
    port map (
            O => \N__46270\,
            I => \N__46264\
        );

    \I__10831\ : Odrv12
    port map (
            O => \N__46267\,
            I => \pwm_generator_inst.un2_threshold_2_1_15\
        );

    \I__10830\ : LocalMux
    port map (
            O => \N__46264\,
            I => \pwm_generator_inst.un2_threshold_2_1_15\
        );

    \I__10829\ : CascadeMux
    port map (
            O => \N__46259\,
            I => \N__46256\
        );

    \I__10828\ : InMux
    port map (
            O => \N__46256\,
            I => \N__46250\
        );

    \I__10827\ : CascadeMux
    port map (
            O => \N__46255\,
            I => \N__46244\
        );

    \I__10826\ : CascadeMux
    port map (
            O => \N__46254\,
            I => \N__46239\
        );

    \I__10825\ : CascadeMux
    port map (
            O => \N__46253\,
            I => \N__46236\
        );

    \I__10824\ : LocalMux
    port map (
            O => \N__46250\,
            I => \N__46228\
        );

    \I__10823\ : InMux
    port map (
            O => \N__46249\,
            I => \N__46219\
        );

    \I__10822\ : InMux
    port map (
            O => \N__46248\,
            I => \N__46219\
        );

    \I__10821\ : InMux
    port map (
            O => \N__46247\,
            I => \N__46219\
        );

    \I__10820\ : InMux
    port map (
            O => \N__46244\,
            I => \N__46219\
        );

    \I__10819\ : InMux
    port map (
            O => \N__46243\,
            I => \N__46210\
        );

    \I__10818\ : InMux
    port map (
            O => \N__46242\,
            I => \N__46210\
        );

    \I__10817\ : InMux
    port map (
            O => \N__46239\,
            I => \N__46210\
        );

    \I__10816\ : InMux
    port map (
            O => \N__46236\,
            I => \N__46210\
        );

    \I__10815\ : InMux
    port map (
            O => \N__46235\,
            I => \N__46203\
        );

    \I__10814\ : InMux
    port map (
            O => \N__46234\,
            I => \N__46203\
        );

    \I__10813\ : InMux
    port map (
            O => \N__46233\,
            I => \N__46196\
        );

    \I__10812\ : InMux
    port map (
            O => \N__46232\,
            I => \N__46196\
        );

    \I__10811\ : InMux
    port map (
            O => \N__46231\,
            I => \N__46196\
        );

    \I__10810\ : Span4Mux_v
    port map (
            O => \N__46228\,
            I => \N__46191\
        );

    \I__10809\ : LocalMux
    port map (
            O => \N__46219\,
            I => \N__46191\
        );

    \I__10808\ : LocalMux
    port map (
            O => \N__46210\,
            I => \N__46188\
        );

    \I__10807\ : InMux
    port map (
            O => \N__46209\,
            I => \N__46185\
        );

    \I__10806\ : CascadeMux
    port map (
            O => \N__46208\,
            I => \N__46166\
        );

    \I__10805\ : LocalMux
    port map (
            O => \N__46203\,
            I => \N__46163\
        );

    \I__10804\ : LocalMux
    port map (
            O => \N__46196\,
            I => \N__46160\
        );

    \I__10803\ : Span4Mux_h
    port map (
            O => \N__46191\,
            I => \N__46155\
        );

    \I__10802\ : Span4Mux_v
    port map (
            O => \N__46188\,
            I => \N__46155\
        );

    \I__10801\ : LocalMux
    port map (
            O => \N__46185\,
            I => \N__46152\
        );

    \I__10800\ : InMux
    port map (
            O => \N__46184\,
            I => \N__46135\
        );

    \I__10799\ : InMux
    port map (
            O => \N__46183\,
            I => \N__46135\
        );

    \I__10798\ : InMux
    port map (
            O => \N__46182\,
            I => \N__46135\
        );

    \I__10797\ : InMux
    port map (
            O => \N__46181\,
            I => \N__46135\
        );

    \I__10796\ : InMux
    port map (
            O => \N__46180\,
            I => \N__46135\
        );

    \I__10795\ : InMux
    port map (
            O => \N__46179\,
            I => \N__46135\
        );

    \I__10794\ : InMux
    port map (
            O => \N__46178\,
            I => \N__46135\
        );

    \I__10793\ : InMux
    port map (
            O => \N__46177\,
            I => \N__46135\
        );

    \I__10792\ : InMux
    port map (
            O => \N__46176\,
            I => \N__46120\
        );

    \I__10791\ : InMux
    port map (
            O => \N__46175\,
            I => \N__46120\
        );

    \I__10790\ : InMux
    port map (
            O => \N__46174\,
            I => \N__46120\
        );

    \I__10789\ : InMux
    port map (
            O => \N__46173\,
            I => \N__46120\
        );

    \I__10788\ : InMux
    port map (
            O => \N__46172\,
            I => \N__46120\
        );

    \I__10787\ : InMux
    port map (
            O => \N__46171\,
            I => \N__46120\
        );

    \I__10786\ : InMux
    port map (
            O => \N__46170\,
            I => \N__46120\
        );

    \I__10785\ : InMux
    port map (
            O => \N__46169\,
            I => \N__46117\
        );

    \I__10784\ : InMux
    port map (
            O => \N__46166\,
            I => \N__46114\
        );

    \I__10783\ : Span4Mux_v
    port map (
            O => \N__46163\,
            I => \N__46111\
        );

    \I__10782\ : Sp12to4
    port map (
            O => \N__46160\,
            I => \N__46108\
        );

    \I__10781\ : Span4Mux_h
    port map (
            O => \N__46155\,
            I => \N__46105\
        );

    \I__10780\ : Sp12to4
    port map (
            O => \N__46152\,
            I => \N__46098\
        );

    \I__10779\ : LocalMux
    port map (
            O => \N__46135\,
            I => \N__46098\
        );

    \I__10778\ : LocalMux
    port map (
            O => \N__46120\,
            I => \N__46098\
        );

    \I__10777\ : LocalMux
    port map (
            O => \N__46117\,
            I => \N__46089\
        );

    \I__10776\ : LocalMux
    port map (
            O => \N__46114\,
            I => \N__46089\
        );

    \I__10775\ : Sp12to4
    port map (
            O => \N__46111\,
            I => \N__46089\
        );

    \I__10774\ : Span12Mux_s7_v
    port map (
            O => \N__46108\,
            I => \N__46089\
        );

    \I__10773\ : Sp12to4
    port map (
            O => \N__46105\,
            I => \N__46082\
        );

    \I__10772\ : Span12Mux_s7_v
    port map (
            O => \N__46098\,
            I => \N__46082\
        );

    \I__10771\ : Span12Mux_h
    port map (
            O => \N__46089\,
            I => \N__46082\
        );

    \I__10770\ : Odrv12
    port map (
            O => \N__46082\,
            I => \N_19_1\
        );

    \I__10769\ : InMux
    port map (
            O => \N__46079\,
            I => \N__46076\
        );

    \I__10768\ : LocalMux
    port map (
            O => \N__46076\,
            I => \N__46068\
        );

    \I__10767\ : InMux
    port map (
            O => \N__46075\,
            I => \N__46065\
        );

    \I__10766\ : CascadeMux
    port map (
            O => \N__46074\,
            I => \N__46061\
        );

    \I__10765\ : CascadeMux
    port map (
            O => \N__46073\,
            I => \N__46058\
        );

    \I__10764\ : CascadeMux
    port map (
            O => \N__46072\,
            I => \N__46054\
        );

    \I__10763\ : CascadeMux
    port map (
            O => \N__46071\,
            I => \N__46051\
        );

    \I__10762\ : Span12Mux_s7_v
    port map (
            O => \N__46068\,
            I => \N__46048\
        );

    \I__10761\ : LocalMux
    port map (
            O => \N__46065\,
            I => \N__46045\
        );

    \I__10760\ : InMux
    port map (
            O => \N__46064\,
            I => \N__46038\
        );

    \I__10759\ : InMux
    port map (
            O => \N__46061\,
            I => \N__46038\
        );

    \I__10758\ : InMux
    port map (
            O => \N__46058\,
            I => \N__46038\
        );

    \I__10757\ : InMux
    port map (
            O => \N__46057\,
            I => \N__46031\
        );

    \I__10756\ : InMux
    port map (
            O => \N__46054\,
            I => \N__46031\
        );

    \I__10755\ : InMux
    port map (
            O => \N__46051\,
            I => \N__46031\
        );

    \I__10754\ : Span12Mux_h
    port map (
            O => \N__46048\,
            I => \N__46028\
        );

    \I__10753\ : Span4Mux_v
    port map (
            O => \N__46045\,
            I => \N__46021\
        );

    \I__10752\ : LocalMux
    port map (
            O => \N__46038\,
            I => \N__46021\
        );

    \I__10751\ : LocalMux
    port map (
            O => \N__46031\,
            I => \N__46021\
        );

    \I__10750\ : Span12Mux_h
    port map (
            O => \N__46028\,
            I => \N__46018\
        );

    \I__10749\ : Span4Mux_h
    port map (
            O => \N__46021\,
            I => \N__46015\
        );

    \I__10748\ : Odrv12
    port map (
            O => \N__46018\,
            I => \pwm_generator_inst.un2_threshold_1_25\
        );

    \I__10747\ : Odrv4
    port map (
            O => \N__46015\,
            I => \pwm_generator_inst.un2_threshold_1_25\
        );

    \I__10746\ : CascadeMux
    port map (
            O => \N__46010\,
            I => \N__46007\
        );

    \I__10745\ : InMux
    port map (
            O => \N__46007\,
            I => \N__46004\
        );

    \I__10744\ : LocalMux
    port map (
            O => \N__46004\,
            I => \N__46001\
        );

    \I__10743\ : Span12Mux_s7_h
    port map (
            O => \N__46001\,
            I => \N__45998\
        );

    \I__10742\ : Span12Mux_h
    port map (
            O => \N__45998\,
            I => \N__45995\
        );

    \I__10741\ : Odrv12
    port map (
            O => \N__45995\,
            I => \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\
        );

    \I__10740\ : InMux
    port map (
            O => \N__45992\,
            I => \N__45986\
        );

    \I__10739\ : InMux
    port map (
            O => \N__45991\,
            I => \N__45986\
        );

    \I__10738\ : LocalMux
    port map (
            O => \N__45986\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_24\
        );

    \I__10737\ : CascadeMux
    port map (
            O => \N__45983\,
            I => \N__45980\
        );

    \I__10736\ : InMux
    port map (
            O => \N__45980\,
            I => \N__45974\
        );

    \I__10735\ : InMux
    port map (
            O => \N__45979\,
            I => \N__45974\
        );

    \I__10734\ : LocalMux
    port map (
            O => \N__45974\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_27\
        );

    \I__10733\ : InMux
    port map (
            O => \N__45971\,
            I => \N__45967\
        );

    \I__10732\ : InMux
    port map (
            O => \N__45970\,
            I => \N__45964\
        );

    \I__10731\ : LocalMux
    port map (
            O => \N__45967\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\
        );

    \I__10730\ : LocalMux
    port map (
            O => \N__45964\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\
        );

    \I__10729\ : CEMux
    port map (
            O => \N__45959\,
            I => \N__45935\
        );

    \I__10728\ : CEMux
    port map (
            O => \N__45958\,
            I => \N__45935\
        );

    \I__10727\ : CEMux
    port map (
            O => \N__45957\,
            I => \N__45935\
        );

    \I__10726\ : CEMux
    port map (
            O => \N__45956\,
            I => \N__45935\
        );

    \I__10725\ : CEMux
    port map (
            O => \N__45955\,
            I => \N__45935\
        );

    \I__10724\ : CEMux
    port map (
            O => \N__45954\,
            I => \N__45935\
        );

    \I__10723\ : CEMux
    port map (
            O => \N__45953\,
            I => \N__45935\
        );

    \I__10722\ : CEMux
    port map (
            O => \N__45952\,
            I => \N__45935\
        );

    \I__10721\ : GlobalMux
    port map (
            O => \N__45935\,
            I => \N__45932\
        );

    \I__10720\ : gio2CtrlBuf
    port map (
            O => \N__45932\,
            I => \phase_controller_inst2.stoper_tr.un1_start_g\
        );

    \I__10719\ : InMux
    port map (
            O => \N__45929\,
            I => \N__45923\
        );

    \I__10718\ : InMux
    port map (
            O => \N__45928\,
            I => \N__45920\
        );

    \I__10717\ : InMux
    port map (
            O => \N__45927\,
            I => \N__45917\
        );

    \I__10716\ : InMux
    port map (
            O => \N__45926\,
            I => \N__45914\
        );

    \I__10715\ : LocalMux
    port map (
            O => \N__45923\,
            I => \N__45911\
        );

    \I__10714\ : LocalMux
    port map (
            O => \N__45920\,
            I => \N__45906\
        );

    \I__10713\ : LocalMux
    port map (
            O => \N__45917\,
            I => \N__45906\
        );

    \I__10712\ : LocalMux
    port map (
            O => \N__45914\,
            I => \N__45903\
        );

    \I__10711\ : Span4Mux_h
    port map (
            O => \N__45911\,
            I => \N__45900\
        );

    \I__10710\ : Span4Mux_h
    port map (
            O => \N__45906\,
            I => \N__45895\
        );

    \I__10709\ : Span4Mux_v
    port map (
            O => \N__45903\,
            I => \N__45895\
        );

    \I__10708\ : Span4Mux_h
    port map (
            O => \N__45900\,
            I => \N__45892\
        );

    \I__10707\ : Span4Mux_h
    port map (
            O => \N__45895\,
            I => \N__45889\
        );

    \I__10706\ : Odrv4
    port map (
            O => \N__45892\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__10705\ : Odrv4
    port map (
            O => \N__45889\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__10704\ : InMux
    port map (
            O => \N__45884\,
            I => \N__45879\
        );

    \I__10703\ : InMux
    port map (
            O => \N__45883\,
            I => \N__45876\
        );

    \I__10702\ : InMux
    port map (
            O => \N__45882\,
            I => \N__45873\
        );

    \I__10701\ : LocalMux
    port map (
            O => \N__45879\,
            I => \N__45868\
        );

    \I__10700\ : LocalMux
    port map (
            O => \N__45876\,
            I => \N__45868\
        );

    \I__10699\ : LocalMux
    port map (
            O => \N__45873\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29\
        );

    \I__10698\ : Odrv4
    port map (
            O => \N__45868\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29\
        );

    \I__10697\ : InMux
    port map (
            O => \N__45863\,
            I => \N__45859\
        );

    \I__10696\ : InMux
    port map (
            O => \N__45862\,
            I => \N__45855\
        );

    \I__10695\ : LocalMux
    port map (
            O => \N__45859\,
            I => \N__45852\
        );

    \I__10694\ : InMux
    port map (
            O => \N__45858\,
            I => \N__45849\
        );

    \I__10693\ : LocalMux
    port map (
            O => \N__45855\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24\
        );

    \I__10692\ : Odrv4
    port map (
            O => \N__45852\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24\
        );

    \I__10691\ : LocalMux
    port map (
            O => \N__45849\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24\
        );

    \I__10690\ : InMux
    port map (
            O => \N__45842\,
            I => \N__45837\
        );

    \I__10689\ : InMux
    port map (
            O => \N__45841\,
            I => \N__45834\
        );

    \I__10688\ : CascadeMux
    port map (
            O => \N__45840\,
            I => \N__45831\
        );

    \I__10687\ : LocalMux
    port map (
            O => \N__45837\,
            I => \N__45827\
        );

    \I__10686\ : LocalMux
    port map (
            O => \N__45834\,
            I => \N__45824\
        );

    \I__10685\ : InMux
    port map (
            O => \N__45831\,
            I => \N__45821\
        );

    \I__10684\ : InMux
    port map (
            O => \N__45830\,
            I => \N__45818\
        );

    \I__10683\ : Span4Mux_v
    port map (
            O => \N__45827\,
            I => \N__45815\
        );

    \I__10682\ : Span4Mux_h
    port map (
            O => \N__45824\,
            I => \N__45812\
        );

    \I__10681\ : LocalMux
    port map (
            O => \N__45821\,
            I => \N__45809\
        );

    \I__10680\ : LocalMux
    port map (
            O => \N__45818\,
            I => \N__45806\
        );

    \I__10679\ : Span4Mux_h
    port map (
            O => \N__45815\,
            I => \N__45803\
        );

    \I__10678\ : Span4Mux_h
    port map (
            O => \N__45812\,
            I => \N__45800\
        );

    \I__10677\ : Span12Mux_s11_v
    port map (
            O => \N__45809\,
            I => \N__45797\
        );

    \I__10676\ : Odrv12
    port map (
            O => \N__45806\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__10675\ : Odrv4
    port map (
            O => \N__45803\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__10674\ : Odrv4
    port map (
            O => \N__45800\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__10673\ : Odrv12
    port map (
            O => \N__45797\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__10672\ : InMux
    port map (
            O => \N__45788\,
            I => \N__45783\
        );

    \I__10671\ : InMux
    port map (
            O => \N__45787\,
            I => \N__45780\
        );

    \I__10670\ : InMux
    port map (
            O => \N__45786\,
            I => \N__45777\
        );

    \I__10669\ : LocalMux
    port map (
            O => \N__45783\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26\
        );

    \I__10668\ : LocalMux
    port map (
            O => \N__45780\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26\
        );

    \I__10667\ : LocalMux
    port map (
            O => \N__45777\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26\
        );

    \I__10666\ : InMux
    port map (
            O => \N__45770\,
            I => \N__45766\
        );

    \I__10665\ : InMux
    port map (
            O => \N__45769\,
            I => \N__45763\
        );

    \I__10664\ : LocalMux
    port map (
            O => \N__45766\,
            I => \N__45758\
        );

    \I__10663\ : LocalMux
    port map (
            O => \N__45763\,
            I => \N__45758\
        );

    \I__10662\ : Span4Mux_v
    port map (
            O => \N__45758\,
            I => \N__45753\
        );

    \I__10661\ : InMux
    port map (
            O => \N__45757\,
            I => \N__45750\
        );

    \I__10660\ : InMux
    port map (
            O => \N__45756\,
            I => \N__45747\
        );

    \I__10659\ : Sp12to4
    port map (
            O => \N__45753\,
            I => \N__45742\
        );

    \I__10658\ : LocalMux
    port map (
            O => \N__45750\,
            I => \N__45742\
        );

    \I__10657\ : LocalMux
    port map (
            O => \N__45747\,
            I => \N__45739\
        );

    \I__10656\ : Span12Mux_s10_h
    port map (
            O => \N__45742\,
            I => \N__45736\
        );

    \I__10655\ : Odrv12
    port map (
            O => \N__45739\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__10654\ : Odrv12
    port map (
            O => \N__45736\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__10653\ : CascadeMux
    port map (
            O => \N__45731\,
            I => \N__45728\
        );

    \I__10652\ : InMux
    port map (
            O => \N__45728\,
            I => \N__45725\
        );

    \I__10651\ : LocalMux
    port map (
            O => \N__45725\,
            I => \N__45722\
        );

    \I__10650\ : Span4Mux_h
    port map (
            O => \N__45722\,
            I => \N__45719\
        );

    \I__10649\ : Span4Mux_h
    port map (
            O => \N__45719\,
            I => \N__45716\
        );

    \I__10648\ : Odrv4
    port map (
            O => \N__45716\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28\
        );

    \I__10647\ : InMux
    port map (
            O => \N__45713\,
            I => \N__45709\
        );

    \I__10646\ : InMux
    port map (
            O => \N__45712\,
            I => \N__45706\
        );

    \I__10645\ : LocalMux
    port map (
            O => \N__45709\,
            I => \N__45699\
        );

    \I__10644\ : LocalMux
    port map (
            O => \N__45706\,
            I => \N__45699\
        );

    \I__10643\ : InMux
    port map (
            O => \N__45705\,
            I => \N__45696\
        );

    \I__10642\ : InMux
    port map (
            O => \N__45704\,
            I => \N__45693\
        );

    \I__10641\ : Span4Mux_v
    port map (
            O => \N__45699\,
            I => \N__45688\
        );

    \I__10640\ : LocalMux
    port map (
            O => \N__45696\,
            I => \N__45688\
        );

    \I__10639\ : LocalMux
    port map (
            O => \N__45693\,
            I => \N__45685\
        );

    \I__10638\ : Span4Mux_h
    port map (
            O => \N__45688\,
            I => \N__45682\
        );

    \I__10637\ : Span4Mux_h
    port map (
            O => \N__45685\,
            I => \N__45679\
        );

    \I__10636\ : Span4Mux_v
    port map (
            O => \N__45682\,
            I => \N__45676\
        );

    \I__10635\ : Span4Mux_v
    port map (
            O => \N__45679\,
            I => \N__45673\
        );

    \I__10634\ : Odrv4
    port map (
            O => \N__45676\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__10633\ : Odrv4
    port map (
            O => \N__45673\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__10632\ : InMux
    port map (
            O => \N__45668\,
            I => \N__45664\
        );

    \I__10631\ : InMux
    port map (
            O => \N__45667\,
            I => \N__45660\
        );

    \I__10630\ : LocalMux
    port map (
            O => \N__45664\,
            I => \N__45657\
        );

    \I__10629\ : InMux
    port map (
            O => \N__45663\,
            I => \N__45654\
        );

    \I__10628\ : LocalMux
    port map (
            O => \N__45660\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28\
        );

    \I__10627\ : Odrv4
    port map (
            O => \N__45657\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28\
        );

    \I__10626\ : LocalMux
    port map (
            O => \N__45654\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28\
        );

    \I__10625\ : InMux
    port map (
            O => \N__45647\,
            I => \N__45644\
        );

    \I__10624\ : LocalMux
    port map (
            O => \N__45644\,
            I => \N__45641\
        );

    \I__10623\ : Odrv12
    port map (
            O => \N__45641\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28\
        );

    \I__10622\ : InMux
    port map (
            O => \N__45638\,
            I => \N__45632\
        );

    \I__10621\ : InMux
    port map (
            O => \N__45637\,
            I => \N__45632\
        );

    \I__10620\ : LocalMux
    port map (
            O => \N__45632\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_29\
        );

    \I__10619\ : InMux
    port map (
            O => \N__45629\,
            I => \N__45623\
        );

    \I__10618\ : InMux
    port map (
            O => \N__45628\,
            I => \N__45623\
        );

    \I__10617\ : LocalMux
    port map (
            O => \N__45623\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_28\
        );

    \I__10616\ : CascadeMux
    port map (
            O => \N__45620\,
            I => \N__45616\
        );

    \I__10615\ : InMux
    port map (
            O => \N__45619\,
            I => \N__45610\
        );

    \I__10614\ : InMux
    port map (
            O => \N__45616\,
            I => \N__45610\
        );

    \I__10613\ : InMux
    port map (
            O => \N__45615\,
            I => \N__45607\
        );

    \I__10612\ : LocalMux
    port map (
            O => \N__45610\,
            I => \N__45604\
        );

    \I__10611\ : LocalMux
    port map (
            O => \N__45607\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__10610\ : Odrv4
    port map (
            O => \N__45604\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__10609\ : CascadeMux
    port map (
            O => \N__45599\,
            I => \N__45595\
        );

    \I__10608\ : InMux
    port map (
            O => \N__45598\,
            I => \N__45589\
        );

    \I__10607\ : InMux
    port map (
            O => \N__45595\,
            I => \N__45589\
        );

    \I__10606\ : InMux
    port map (
            O => \N__45594\,
            I => \N__45586\
        );

    \I__10605\ : LocalMux
    port map (
            O => \N__45589\,
            I => \N__45583\
        );

    \I__10604\ : LocalMux
    port map (
            O => \N__45586\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__10603\ : Odrv4
    port map (
            O => \N__45583\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__10602\ : CascadeMux
    port map (
            O => \N__45578\,
            I => \N__45575\
        );

    \I__10601\ : InMux
    port map (
            O => \N__45575\,
            I => \N__45572\
        );

    \I__10600\ : LocalMux
    port map (
            O => \N__45572\,
            I => \N__45569\
        );

    \I__10599\ : Odrv12
    port map (
            O => \N__45569\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt28\
        );

    \I__10598\ : InMux
    port map (
            O => \N__45566\,
            I => \N__45563\
        );

    \I__10597\ : LocalMux
    port map (
            O => \N__45563\,
            I => \N__45560\
        );

    \I__10596\ : Odrv12
    port map (
            O => \N__45560\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt26\
        );

    \I__10595\ : InMux
    port map (
            O => \N__45557\,
            I => \N__45552\
        );

    \I__10594\ : InMux
    port map (
            O => \N__45556\,
            I => \N__45549\
        );

    \I__10593\ : InMux
    port map (
            O => \N__45555\,
            I => \N__45546\
        );

    \I__10592\ : LocalMux
    port map (
            O => \N__45552\,
            I => \N__45543\
        );

    \I__10591\ : LocalMux
    port map (
            O => \N__45549\,
            I => \N__45540\
        );

    \I__10590\ : LocalMux
    port map (
            O => \N__45546\,
            I => \N__45536\
        );

    \I__10589\ : Span4Mux_h
    port map (
            O => \N__45543\,
            I => \N__45531\
        );

    \I__10588\ : Span4Mux_v
    port map (
            O => \N__45540\,
            I => \N__45531\
        );

    \I__10587\ : CascadeMux
    port map (
            O => \N__45539\,
            I => \N__45528\
        );

    \I__10586\ : Sp12to4
    port map (
            O => \N__45536\,
            I => \N__45525\
        );

    \I__10585\ : Span4Mux_v
    port map (
            O => \N__45531\,
            I => \N__45522\
        );

    \I__10584\ : InMux
    port map (
            O => \N__45528\,
            I => \N__45519\
        );

    \I__10583\ : Span12Mux_v
    port map (
            O => \N__45525\,
            I => \N__45516\
        );

    \I__10582\ : Span4Mux_h
    port map (
            O => \N__45522\,
            I => \N__45513\
        );

    \I__10581\ : LocalMux
    port map (
            O => \N__45519\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__10580\ : Odrv12
    port map (
            O => \N__45516\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__10579\ : Odrv4
    port map (
            O => \N__45513\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__10578\ : CascadeMux
    port map (
            O => \N__45506\,
            I => \N__45503\
        );

    \I__10577\ : InMux
    port map (
            O => \N__45503\,
            I => \N__45500\
        );

    \I__10576\ : LocalMux
    port map (
            O => \N__45500\,
            I => \N__45494\
        );

    \I__10575\ : InMux
    port map (
            O => \N__45499\,
            I => \N__45489\
        );

    \I__10574\ : InMux
    port map (
            O => \N__45498\,
            I => \N__45489\
        );

    \I__10573\ : InMux
    port map (
            O => \N__45497\,
            I => \N__45485\
        );

    \I__10572\ : Span4Mux_h
    port map (
            O => \N__45494\,
            I => \N__45482\
        );

    \I__10571\ : LocalMux
    port map (
            O => \N__45489\,
            I => \N__45479\
        );

    \I__10570\ : InMux
    port map (
            O => \N__45488\,
            I => \N__45476\
        );

    \I__10569\ : LocalMux
    port map (
            O => \N__45485\,
            I => \N__45473\
        );

    \I__10568\ : Span4Mux_h
    port map (
            O => \N__45482\,
            I => \N__45470\
        );

    \I__10567\ : Span4Mux_h
    port map (
            O => \N__45479\,
            I => \N__45467\
        );

    \I__10566\ : LocalMux
    port map (
            O => \N__45476\,
            I => \N__45462\
        );

    \I__10565\ : Span4Mux_h
    port map (
            O => \N__45473\,
            I => \N__45462\
        );

    \I__10564\ : Span4Mux_v
    port map (
            O => \N__45470\,
            I => \N__45457\
        );

    \I__10563\ : Span4Mux_v
    port map (
            O => \N__45467\,
            I => \N__45457\
        );

    \I__10562\ : Span4Mux_v
    port map (
            O => \N__45462\,
            I => \N__45454\
        );

    \I__10561\ : Odrv4
    port map (
            O => \N__45457\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__10560\ : Odrv4
    port map (
            O => \N__45454\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__10559\ : CascadeMux
    port map (
            O => \N__45449\,
            I => \N__45445\
        );

    \I__10558\ : InMux
    port map (
            O => \N__45448\,
            I => \N__45440\
        );

    \I__10557\ : InMux
    port map (
            O => \N__45445\,
            I => \N__45440\
        );

    \I__10556\ : LocalMux
    port map (
            O => \N__45440\,
            I => \N__45437\
        );

    \I__10555\ : Span4Mux_h
    port map (
            O => \N__45437\,
            I => \N__45433\
        );

    \I__10554\ : InMux
    port map (
            O => \N__45436\,
            I => \N__45430\
        );

    \I__10553\ : Span4Mux_h
    port map (
            O => \N__45433\,
            I => \N__45427\
        );

    \I__10552\ : LocalMux
    port map (
            O => \N__45430\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__10551\ : Odrv4
    port map (
            O => \N__45427\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__10550\ : CascadeMux
    port map (
            O => \N__45422\,
            I => \N__45419\
        );

    \I__10549\ : InMux
    port map (
            O => \N__45419\,
            I => \N__45415\
        );

    \I__10548\ : InMux
    port map (
            O => \N__45418\,
            I => \N__45412\
        );

    \I__10547\ : LocalMux
    port map (
            O => \N__45415\,
            I => \N__45407\
        );

    \I__10546\ : LocalMux
    port map (
            O => \N__45412\,
            I => \N__45407\
        );

    \I__10545\ : Span4Mux_h
    port map (
            O => \N__45407\,
            I => \N__45403\
        );

    \I__10544\ : InMux
    port map (
            O => \N__45406\,
            I => \N__45400\
        );

    \I__10543\ : Span4Mux_h
    port map (
            O => \N__45403\,
            I => \N__45397\
        );

    \I__10542\ : LocalMux
    port map (
            O => \N__45400\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__10541\ : Odrv4
    port map (
            O => \N__45397\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__10540\ : InMux
    port map (
            O => \N__45392\,
            I => \N__45389\
        );

    \I__10539\ : LocalMux
    port map (
            O => \N__45389\,
            I => \N__45386\
        );

    \I__10538\ : Span4Mux_h
    port map (
            O => \N__45386\,
            I => \N__45383\
        );

    \I__10537\ : Odrv4
    port map (
            O => \N__45383\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24\
        );

    \I__10536\ : InMux
    port map (
            O => \N__45380\,
            I => \N__45377\
        );

    \I__10535\ : LocalMux
    port map (
            O => \N__45377\,
            I => \N__45374\
        );

    \I__10534\ : Odrv12
    port map (
            O => \N__45374\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26\
        );

    \I__10533\ : InMux
    port map (
            O => \N__45371\,
            I => \N__45365\
        );

    \I__10532\ : InMux
    port map (
            O => \N__45370\,
            I => \N__45365\
        );

    \I__10531\ : LocalMux
    port map (
            O => \N__45365\,
            I => \N__45362\
        );

    \I__10530\ : Span4Mux_h
    port map (
            O => \N__45362\,
            I => \N__45358\
        );

    \I__10529\ : InMux
    port map (
            O => \N__45361\,
            I => \N__45355\
        );

    \I__10528\ : Span4Mux_h
    port map (
            O => \N__45358\,
            I => \N__45352\
        );

    \I__10527\ : LocalMux
    port map (
            O => \N__45355\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__10526\ : Odrv4
    port map (
            O => \N__45352\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__10525\ : CascadeMux
    port map (
            O => \N__45347\,
            I => \N__45343\
        );

    \I__10524\ : InMux
    port map (
            O => \N__45346\,
            I => \N__45338\
        );

    \I__10523\ : InMux
    port map (
            O => \N__45343\,
            I => \N__45338\
        );

    \I__10522\ : LocalMux
    port map (
            O => \N__45338\,
            I => \N__45334\
        );

    \I__10521\ : InMux
    port map (
            O => \N__45337\,
            I => \N__45331\
        );

    \I__10520\ : Span12Mux_s10_v
    port map (
            O => \N__45334\,
            I => \N__45328\
        );

    \I__10519\ : LocalMux
    port map (
            O => \N__45331\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__10518\ : Odrv12
    port map (
            O => \N__45328\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__10517\ : CascadeMux
    port map (
            O => \N__45323\,
            I => \N__45320\
        );

    \I__10516\ : InMux
    port map (
            O => \N__45320\,
            I => \N__45317\
        );

    \I__10515\ : LocalMux
    port map (
            O => \N__45317\,
            I => \N__45314\
        );

    \I__10514\ : Odrv12
    port map (
            O => \N__45314\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt26\
        );

    \I__10513\ : InMux
    port map (
            O => \N__45311\,
            I => \N__45305\
        );

    \I__10512\ : InMux
    port map (
            O => \N__45310\,
            I => \N__45305\
        );

    \I__10511\ : LocalMux
    port map (
            O => \N__45305\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_26\
        );

    \I__10510\ : InMux
    port map (
            O => \N__45302\,
            I => \N__45299\
        );

    \I__10509\ : LocalMux
    port map (
            O => \N__45299\,
            I => \N__45296\
        );

    \I__10508\ : Span4Mux_h
    port map (
            O => \N__45296\,
            I => \N__45293\
        );

    \I__10507\ : Span4Mux_h
    port map (
            O => \N__45293\,
            I => \N__45290\
        );

    \I__10506\ : Odrv4
    port map (
            O => \N__45290\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt28\
        );

    \I__10505\ : InMux
    port map (
            O => \N__45287\,
            I => \N__45281\
        );

    \I__10504\ : InMux
    port map (
            O => \N__45286\,
            I => \N__45281\
        );

    \I__10503\ : LocalMux
    port map (
            O => \N__45281\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_28\
        );

    \I__10502\ : InMux
    port map (
            O => \N__45278\,
            I => \N__45273\
        );

    \I__10501\ : InMux
    port map (
            O => \N__45277\,
            I => \N__45270\
        );

    \I__10500\ : InMux
    port map (
            O => \N__45276\,
            I => \N__45267\
        );

    \I__10499\ : LocalMux
    port map (
            O => \N__45273\,
            I => \N__45262\
        );

    \I__10498\ : LocalMux
    port map (
            O => \N__45270\,
            I => \N__45262\
        );

    \I__10497\ : LocalMux
    port map (
            O => \N__45267\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__10496\ : Odrv12
    port map (
            O => \N__45262\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__10495\ : CascadeMux
    port map (
            O => \N__45257\,
            I => \N__45253\
        );

    \I__10494\ : CascadeMux
    port map (
            O => \N__45256\,
            I => \N__45250\
        );

    \I__10493\ : InMux
    port map (
            O => \N__45253\,
            I => \N__45247\
        );

    \I__10492\ : InMux
    port map (
            O => \N__45250\,
            I => \N__45244\
        );

    \I__10491\ : LocalMux
    port map (
            O => \N__45247\,
            I => \N__45238\
        );

    \I__10490\ : LocalMux
    port map (
            O => \N__45244\,
            I => \N__45238\
        );

    \I__10489\ : InMux
    port map (
            O => \N__45243\,
            I => \N__45235\
        );

    \I__10488\ : Span4Mux_h
    port map (
            O => \N__45238\,
            I => \N__45232\
        );

    \I__10487\ : LocalMux
    port map (
            O => \N__45235\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__10486\ : Odrv4
    port map (
            O => \N__45232\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__10485\ : InMux
    port map (
            O => \N__45227\,
            I => \N__45221\
        );

    \I__10484\ : InMux
    port map (
            O => \N__45226\,
            I => \N__45221\
        );

    \I__10483\ : LocalMux
    port map (
            O => \N__45221\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\
        );

    \I__10482\ : InMux
    port map (
            O => \N__45218\,
            I => \N__45212\
        );

    \I__10481\ : InMux
    port map (
            O => \N__45217\,
            I => \N__45212\
        );

    \I__10480\ : LocalMux
    port map (
            O => \N__45212\,
            I => \N__45208\
        );

    \I__10479\ : InMux
    port map (
            O => \N__45211\,
            I => \N__45205\
        );

    \I__10478\ : Span4Mux_v
    port map (
            O => \N__45208\,
            I => \N__45202\
        );

    \I__10477\ : LocalMux
    port map (
            O => \N__45205\,
            I => \N__45199\
        );

    \I__10476\ : Odrv4
    port map (
            O => \N__45202\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__10475\ : Odrv12
    port map (
            O => \N__45199\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__10474\ : InMux
    port map (
            O => \N__45194\,
            I => \N__45191\
        );

    \I__10473\ : LocalMux
    port map (
            O => \N__45191\,
            I => \N__45187\
        );

    \I__10472\ : CascadeMux
    port map (
            O => \N__45190\,
            I => \N__45183\
        );

    \I__10471\ : Span4Mux_h
    port map (
            O => \N__45187\,
            I => \N__45179\
        );

    \I__10470\ : InMux
    port map (
            O => \N__45186\,
            I => \N__45172\
        );

    \I__10469\ : InMux
    port map (
            O => \N__45183\,
            I => \N__45172\
        );

    \I__10468\ : InMux
    port map (
            O => \N__45182\,
            I => \N__45172\
        );

    \I__10467\ : Odrv4
    port map (
            O => \N__45179\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__10466\ : LocalMux
    port map (
            O => \N__45172\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__10465\ : CascadeMux
    port map (
            O => \N__45167\,
            I => \N__45163\
        );

    \I__10464\ : InMux
    port map (
            O => \N__45166\,
            I => \N__45158\
        );

    \I__10463\ : InMux
    port map (
            O => \N__45163\,
            I => \N__45158\
        );

    \I__10462\ : LocalMux
    port map (
            O => \N__45158\,
            I => \N__45154\
        );

    \I__10461\ : InMux
    port map (
            O => \N__45157\,
            I => \N__45151\
        );

    \I__10460\ : Span4Mux_v
    port map (
            O => \N__45154\,
            I => \N__45147\
        );

    \I__10459\ : LocalMux
    port map (
            O => \N__45151\,
            I => \N__45144\
        );

    \I__10458\ : InMux
    port map (
            O => \N__45150\,
            I => \N__45141\
        );

    \I__10457\ : Span4Mux_h
    port map (
            O => \N__45147\,
            I => \N__45136\
        );

    \I__10456\ : Span4Mux_h
    port map (
            O => \N__45144\,
            I => \N__45136\
        );

    \I__10455\ : LocalMux
    port map (
            O => \N__45141\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__10454\ : Odrv4
    port map (
            O => \N__45136\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__10453\ : CascadeMux
    port map (
            O => \N__45131\,
            I => \N__45128\
        );

    \I__10452\ : InMux
    port map (
            O => \N__45128\,
            I => \N__45125\
        );

    \I__10451\ : LocalMux
    port map (
            O => \N__45125\,
            I => \N__45122\
        );

    \I__10450\ : Span4Mux_h
    port map (
            O => \N__45122\,
            I => \N__45119\
        );

    \I__10449\ : Span4Mux_h
    port map (
            O => \N__45119\,
            I => \N__45116\
        );

    \I__10448\ : Odrv4
    port map (
            O => \N__45116\,
            I => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\
        );

    \I__10447\ : CascadeMux
    port map (
            O => \N__45113\,
            I => \N__45110\
        );

    \I__10446\ : InMux
    port map (
            O => \N__45110\,
            I => \N__45107\
        );

    \I__10445\ : LocalMux
    port map (
            O => \N__45107\,
            I => \N__45104\
        );

    \I__10444\ : Odrv12
    port map (
            O => \N__45104\,
            I => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\
        );

    \I__10443\ : InMux
    port map (
            O => \N__45101\,
            I => \N__45095\
        );

    \I__10442\ : InMux
    port map (
            O => \N__45100\,
            I => \N__45095\
        );

    \I__10441\ : LocalMux
    port map (
            O => \N__45095\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__10440\ : CascadeMux
    port map (
            O => \N__45092\,
            I => \N__45089\
        );

    \I__10439\ : InMux
    port map (
            O => \N__45089\,
            I => \N__45083\
        );

    \I__10438\ : InMux
    port map (
            O => \N__45088\,
            I => \N__45083\
        );

    \I__10437\ : LocalMux
    port map (
            O => \N__45083\,
            I => \N__45080\
        );

    \I__10436\ : Span4Mux_v
    port map (
            O => \N__45080\,
            I => \N__45076\
        );

    \I__10435\ : InMux
    port map (
            O => \N__45079\,
            I => \N__45073\
        );

    \I__10434\ : Sp12to4
    port map (
            O => \N__45076\,
            I => \N__45066\
        );

    \I__10433\ : LocalMux
    port map (
            O => \N__45073\,
            I => \N__45066\
        );

    \I__10432\ : InMux
    port map (
            O => \N__45072\,
            I => \N__45061\
        );

    \I__10431\ : InMux
    port map (
            O => \N__45071\,
            I => \N__45061\
        );

    \I__10430\ : Odrv12
    port map (
            O => \N__45066\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__10429\ : LocalMux
    port map (
            O => \N__45061\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__10428\ : CascadeMux
    port map (
            O => \N__45056\,
            I => \N__45047\
        );

    \I__10427\ : CascadeMux
    port map (
            O => \N__45055\,
            I => \N__45040\
        );

    \I__10426\ : CascadeMux
    port map (
            O => \N__45054\,
            I => \N__45024\
        );

    \I__10425\ : CascadeMux
    port map (
            O => \N__45053\,
            I => \N__45020\
        );

    \I__10424\ : CascadeMux
    port map (
            O => \N__45052\,
            I => \N__45016\
        );

    \I__10423\ : CascadeMux
    port map (
            O => \N__45051\,
            I => \N__45000\
        );

    \I__10422\ : InMux
    port map (
            O => \N__45050\,
            I => \N__44989\
        );

    \I__10421\ : InMux
    port map (
            O => \N__45047\,
            I => \N__44989\
        );

    \I__10420\ : CascadeMux
    port map (
            O => \N__45046\,
            I => \N__44986\
        );

    \I__10419\ : CascadeMux
    port map (
            O => \N__45045\,
            I => \N__44983\
        );

    \I__10418\ : CascadeMux
    port map (
            O => \N__45044\,
            I => \N__44980\
        );

    \I__10417\ : CascadeMux
    port map (
            O => \N__45043\,
            I => \N__44976\
        );

    \I__10416\ : InMux
    port map (
            O => \N__45040\,
            I => \N__44966\
        );

    \I__10415\ : CascadeMux
    port map (
            O => \N__45039\,
            I => \N__44962\
        );

    \I__10414\ : CascadeMux
    port map (
            O => \N__45038\,
            I => \N__44958\
        );

    \I__10413\ : CascadeMux
    port map (
            O => \N__45037\,
            I => \N__44955\
        );

    \I__10412\ : InMux
    port map (
            O => \N__45036\,
            I => \N__44949\
        );

    \I__10411\ : InMux
    port map (
            O => \N__45035\,
            I => \N__44949\
        );

    \I__10410\ : InMux
    port map (
            O => \N__45034\,
            I => \N__44939\
        );

    \I__10409\ : InMux
    port map (
            O => \N__45033\,
            I => \N__44939\
        );

    \I__10408\ : InMux
    port map (
            O => \N__45032\,
            I => \N__44939\
        );

    \I__10407\ : InMux
    port map (
            O => \N__45031\,
            I => \N__44939\
        );

    \I__10406\ : CascadeMux
    port map (
            O => \N__45030\,
            I => \N__44928\
        );

    \I__10405\ : CascadeMux
    port map (
            O => \N__45029\,
            I => \N__44920\
        );

    \I__10404\ : InMux
    port map (
            O => \N__45028\,
            I => \N__44902\
        );

    \I__10403\ : InMux
    port map (
            O => \N__45027\,
            I => \N__44902\
        );

    \I__10402\ : InMux
    port map (
            O => \N__45024\,
            I => \N__44902\
        );

    \I__10401\ : InMux
    port map (
            O => \N__45023\,
            I => \N__44902\
        );

    \I__10400\ : InMux
    port map (
            O => \N__45020\,
            I => \N__44902\
        );

    \I__10399\ : InMux
    port map (
            O => \N__45019\,
            I => \N__44902\
        );

    \I__10398\ : InMux
    port map (
            O => \N__45016\,
            I => \N__44902\
        );

    \I__10397\ : InMux
    port map (
            O => \N__45015\,
            I => \N__44902\
        );

    \I__10396\ : CascadeMux
    port map (
            O => \N__45014\,
            I => \N__44899\
        );

    \I__10395\ : CascadeMux
    port map (
            O => \N__45013\,
            I => \N__44895\
        );

    \I__10394\ : CascadeMux
    port map (
            O => \N__45012\,
            I => \N__44891\
        );

    \I__10393\ : CascadeMux
    port map (
            O => \N__45011\,
            I => \N__44887\
        );

    \I__10392\ : CascadeMux
    port map (
            O => \N__45010\,
            I => \N__44883\
        );

    \I__10391\ : CascadeMux
    port map (
            O => \N__45009\,
            I => \N__44879\
        );

    \I__10390\ : CascadeMux
    port map (
            O => \N__45008\,
            I => \N__44875\
        );

    \I__10389\ : CascadeMux
    port map (
            O => \N__45007\,
            I => \N__44871\
        );

    \I__10388\ : CascadeMux
    port map (
            O => \N__45006\,
            I => \N__44867\
        );

    \I__10387\ : CascadeMux
    port map (
            O => \N__45005\,
            I => \N__44863\
        );

    \I__10386\ : CascadeMux
    port map (
            O => \N__45004\,
            I => \N__44859\
        );

    \I__10385\ : InMux
    port map (
            O => \N__45003\,
            I => \N__44853\
        );

    \I__10384\ : InMux
    port map (
            O => \N__45000\,
            I => \N__44853\
        );

    \I__10383\ : CascadeMux
    port map (
            O => \N__44999\,
            I => \N__44847\
        );

    \I__10382\ : CascadeMux
    port map (
            O => \N__44998\,
            I => \N__44844\
        );

    \I__10381\ : CascadeMux
    port map (
            O => \N__44997\,
            I => \N__44841\
        );

    \I__10380\ : CascadeMux
    port map (
            O => \N__44996\,
            I => \N__44838\
        );

    \I__10379\ : CascadeMux
    port map (
            O => \N__44995\,
            I => \N__44835\
        );

    \I__10378\ : CascadeMux
    port map (
            O => \N__44994\,
            I => \N__44830\
        );

    \I__10377\ : LocalMux
    port map (
            O => \N__44989\,
            I => \N__44824\
        );

    \I__10376\ : InMux
    port map (
            O => \N__44986\,
            I => \N__44821\
        );

    \I__10375\ : InMux
    port map (
            O => \N__44983\,
            I => \N__44818\
        );

    \I__10374\ : InMux
    port map (
            O => \N__44980\,
            I => \N__44811\
        );

    \I__10373\ : InMux
    port map (
            O => \N__44979\,
            I => \N__44811\
        );

    \I__10372\ : InMux
    port map (
            O => \N__44976\,
            I => \N__44811\
        );

    \I__10371\ : CascadeMux
    port map (
            O => \N__44975\,
            I => \N__44807\
        );

    \I__10370\ : CascadeMux
    port map (
            O => \N__44974\,
            I => \N__44803\
        );

    \I__10369\ : CascadeMux
    port map (
            O => \N__44973\,
            I => \N__44799\
        );

    \I__10368\ : CascadeMux
    port map (
            O => \N__44972\,
            I => \N__44795\
        );

    \I__10367\ : CascadeMux
    port map (
            O => \N__44971\,
            I => \N__44791\
        );

    \I__10366\ : CascadeMux
    port map (
            O => \N__44970\,
            I => \N__44787\
        );

    \I__10365\ : CascadeMux
    port map (
            O => \N__44969\,
            I => \N__44783\
        );

    \I__10364\ : LocalMux
    port map (
            O => \N__44966\,
            I => \N__44772\
        );

    \I__10363\ : InMux
    port map (
            O => \N__44965\,
            I => \N__44769\
        );

    \I__10362\ : InMux
    port map (
            O => \N__44962\,
            I => \N__44764\
        );

    \I__10361\ : InMux
    port map (
            O => \N__44961\,
            I => \N__44764\
        );

    \I__10360\ : InMux
    port map (
            O => \N__44958\,
            I => \N__44761\
        );

    \I__10359\ : InMux
    port map (
            O => \N__44955\,
            I => \N__44756\
        );

    \I__10358\ : InMux
    port map (
            O => \N__44954\,
            I => \N__44756\
        );

    \I__10357\ : LocalMux
    port map (
            O => \N__44949\,
            I => \N__44753\
        );

    \I__10356\ : InMux
    port map (
            O => \N__44948\,
            I => \N__44750\
        );

    \I__10355\ : LocalMux
    port map (
            O => \N__44939\,
            I => \N__44747\
        );

    \I__10354\ : InMux
    port map (
            O => \N__44938\,
            I => \N__44732\
        );

    \I__10353\ : InMux
    port map (
            O => \N__44937\,
            I => \N__44732\
        );

    \I__10352\ : InMux
    port map (
            O => \N__44936\,
            I => \N__44732\
        );

    \I__10351\ : InMux
    port map (
            O => \N__44935\,
            I => \N__44732\
        );

    \I__10350\ : InMux
    port map (
            O => \N__44934\,
            I => \N__44732\
        );

    \I__10349\ : InMux
    port map (
            O => \N__44933\,
            I => \N__44732\
        );

    \I__10348\ : InMux
    port map (
            O => \N__44932\,
            I => \N__44732\
        );

    \I__10347\ : InMux
    port map (
            O => \N__44931\,
            I => \N__44717\
        );

    \I__10346\ : InMux
    port map (
            O => \N__44928\,
            I => \N__44717\
        );

    \I__10345\ : InMux
    port map (
            O => \N__44927\,
            I => \N__44717\
        );

    \I__10344\ : InMux
    port map (
            O => \N__44926\,
            I => \N__44717\
        );

    \I__10343\ : InMux
    port map (
            O => \N__44925\,
            I => \N__44717\
        );

    \I__10342\ : InMux
    port map (
            O => \N__44924\,
            I => \N__44717\
        );

    \I__10341\ : InMux
    port map (
            O => \N__44923\,
            I => \N__44717\
        );

    \I__10340\ : InMux
    port map (
            O => \N__44920\,
            I => \N__44712\
        );

    \I__10339\ : InMux
    port map (
            O => \N__44919\,
            I => \N__44712\
        );

    \I__10338\ : LocalMux
    port map (
            O => \N__44902\,
            I => \N__44709\
        );

    \I__10337\ : InMux
    port map (
            O => \N__44899\,
            I => \N__44692\
        );

    \I__10336\ : InMux
    port map (
            O => \N__44898\,
            I => \N__44692\
        );

    \I__10335\ : InMux
    port map (
            O => \N__44895\,
            I => \N__44692\
        );

    \I__10334\ : InMux
    port map (
            O => \N__44894\,
            I => \N__44692\
        );

    \I__10333\ : InMux
    port map (
            O => \N__44891\,
            I => \N__44692\
        );

    \I__10332\ : InMux
    port map (
            O => \N__44890\,
            I => \N__44692\
        );

    \I__10331\ : InMux
    port map (
            O => \N__44887\,
            I => \N__44692\
        );

    \I__10330\ : InMux
    port map (
            O => \N__44886\,
            I => \N__44692\
        );

    \I__10329\ : InMux
    port map (
            O => \N__44883\,
            I => \N__44675\
        );

    \I__10328\ : InMux
    port map (
            O => \N__44882\,
            I => \N__44675\
        );

    \I__10327\ : InMux
    port map (
            O => \N__44879\,
            I => \N__44675\
        );

    \I__10326\ : InMux
    port map (
            O => \N__44878\,
            I => \N__44675\
        );

    \I__10325\ : InMux
    port map (
            O => \N__44875\,
            I => \N__44675\
        );

    \I__10324\ : InMux
    port map (
            O => \N__44874\,
            I => \N__44675\
        );

    \I__10323\ : InMux
    port map (
            O => \N__44871\,
            I => \N__44675\
        );

    \I__10322\ : InMux
    port map (
            O => \N__44870\,
            I => \N__44675\
        );

    \I__10321\ : InMux
    port map (
            O => \N__44867\,
            I => \N__44662\
        );

    \I__10320\ : InMux
    port map (
            O => \N__44866\,
            I => \N__44662\
        );

    \I__10319\ : InMux
    port map (
            O => \N__44863\,
            I => \N__44662\
        );

    \I__10318\ : InMux
    port map (
            O => \N__44862\,
            I => \N__44662\
        );

    \I__10317\ : InMux
    port map (
            O => \N__44859\,
            I => \N__44662\
        );

    \I__10316\ : InMux
    port map (
            O => \N__44858\,
            I => \N__44662\
        );

    \I__10315\ : LocalMux
    port map (
            O => \N__44853\,
            I => \N__44659\
        );

    \I__10314\ : InMux
    port map (
            O => \N__44852\,
            I => \N__44652\
        );

    \I__10313\ : InMux
    port map (
            O => \N__44851\,
            I => \N__44652\
        );

    \I__10312\ : InMux
    port map (
            O => \N__44850\,
            I => \N__44652\
        );

    \I__10311\ : InMux
    port map (
            O => \N__44847\,
            I => \N__44645\
        );

    \I__10310\ : InMux
    port map (
            O => \N__44844\,
            I => \N__44645\
        );

    \I__10309\ : InMux
    port map (
            O => \N__44841\,
            I => \N__44645\
        );

    \I__10308\ : InMux
    port map (
            O => \N__44838\,
            I => \N__44628\
        );

    \I__10307\ : InMux
    port map (
            O => \N__44835\,
            I => \N__44628\
        );

    \I__10306\ : InMux
    port map (
            O => \N__44834\,
            I => \N__44628\
        );

    \I__10305\ : InMux
    port map (
            O => \N__44833\,
            I => \N__44628\
        );

    \I__10304\ : InMux
    port map (
            O => \N__44830\,
            I => \N__44628\
        );

    \I__10303\ : InMux
    port map (
            O => \N__44829\,
            I => \N__44628\
        );

    \I__10302\ : InMux
    port map (
            O => \N__44828\,
            I => \N__44628\
        );

    \I__10301\ : InMux
    port map (
            O => \N__44827\,
            I => \N__44628\
        );

    \I__10300\ : Span4Mux_v
    port map (
            O => \N__44824\,
            I => \N__44619\
        );

    \I__10299\ : LocalMux
    port map (
            O => \N__44821\,
            I => \N__44612\
        );

    \I__10298\ : LocalMux
    port map (
            O => \N__44818\,
            I => \N__44612\
        );

    \I__10297\ : LocalMux
    port map (
            O => \N__44811\,
            I => \N__44612\
        );

    \I__10296\ : InMux
    port map (
            O => \N__44810\,
            I => \N__44597\
        );

    \I__10295\ : InMux
    port map (
            O => \N__44807\,
            I => \N__44597\
        );

    \I__10294\ : InMux
    port map (
            O => \N__44806\,
            I => \N__44597\
        );

    \I__10293\ : InMux
    port map (
            O => \N__44803\,
            I => \N__44597\
        );

    \I__10292\ : InMux
    port map (
            O => \N__44802\,
            I => \N__44597\
        );

    \I__10291\ : InMux
    port map (
            O => \N__44799\,
            I => \N__44597\
        );

    \I__10290\ : InMux
    port map (
            O => \N__44798\,
            I => \N__44597\
        );

    \I__10289\ : InMux
    port map (
            O => \N__44795\,
            I => \N__44580\
        );

    \I__10288\ : InMux
    port map (
            O => \N__44794\,
            I => \N__44580\
        );

    \I__10287\ : InMux
    port map (
            O => \N__44791\,
            I => \N__44580\
        );

    \I__10286\ : InMux
    port map (
            O => \N__44790\,
            I => \N__44580\
        );

    \I__10285\ : InMux
    port map (
            O => \N__44787\,
            I => \N__44580\
        );

    \I__10284\ : InMux
    port map (
            O => \N__44786\,
            I => \N__44580\
        );

    \I__10283\ : InMux
    port map (
            O => \N__44783\,
            I => \N__44580\
        );

    \I__10282\ : InMux
    port map (
            O => \N__44782\,
            I => \N__44580\
        );

    \I__10281\ : CascadeMux
    port map (
            O => \N__44781\,
            I => \N__44577\
        );

    \I__10280\ : CascadeMux
    port map (
            O => \N__44780\,
            I => \N__44573\
        );

    \I__10279\ : CascadeMux
    port map (
            O => \N__44779\,
            I => \N__44569\
        );

    \I__10278\ : CascadeMux
    port map (
            O => \N__44778\,
            I => \N__44565\
        );

    \I__10277\ : CascadeMux
    port map (
            O => \N__44777\,
            I => \N__44561\
        );

    \I__10276\ : CascadeMux
    port map (
            O => \N__44776\,
            I => \N__44557\
        );

    \I__10275\ : CascadeMux
    port map (
            O => \N__44775\,
            I => \N__44553\
        );

    \I__10274\ : Span4Mux_h
    port map (
            O => \N__44772\,
            I => \N__44545\
        );

    \I__10273\ : LocalMux
    port map (
            O => \N__44769\,
            I => \N__44545\
        );

    \I__10272\ : LocalMux
    port map (
            O => \N__44764\,
            I => \N__44545\
        );

    \I__10271\ : LocalMux
    port map (
            O => \N__44761\,
            I => \N__44542\
        );

    \I__10270\ : LocalMux
    port map (
            O => \N__44756\,
            I => \N__44539\
        );

    \I__10269\ : Span4Mux_h
    port map (
            O => \N__44753\,
            I => \N__44518\
        );

    \I__10268\ : LocalMux
    port map (
            O => \N__44750\,
            I => \N__44518\
        );

    \I__10267\ : Span4Mux_h
    port map (
            O => \N__44747\,
            I => \N__44518\
        );

    \I__10266\ : LocalMux
    port map (
            O => \N__44732\,
            I => \N__44518\
        );

    \I__10265\ : LocalMux
    port map (
            O => \N__44717\,
            I => \N__44518\
        );

    \I__10264\ : LocalMux
    port map (
            O => \N__44712\,
            I => \N__44518\
        );

    \I__10263\ : Span4Mux_v
    port map (
            O => \N__44709\,
            I => \N__44518\
        );

    \I__10262\ : LocalMux
    port map (
            O => \N__44692\,
            I => \N__44518\
        );

    \I__10261\ : LocalMux
    port map (
            O => \N__44675\,
            I => \N__44518\
        );

    \I__10260\ : LocalMux
    port map (
            O => \N__44662\,
            I => \N__44518\
        );

    \I__10259\ : Span4Mux_h
    port map (
            O => \N__44659\,
            I => \N__44515\
        );

    \I__10258\ : LocalMux
    port map (
            O => \N__44652\,
            I => \N__44508\
        );

    \I__10257\ : LocalMux
    port map (
            O => \N__44645\,
            I => \N__44508\
        );

    \I__10256\ : LocalMux
    port map (
            O => \N__44628\,
            I => \N__44508\
        );

    \I__10255\ : InMux
    port map (
            O => \N__44627\,
            I => \N__44505\
        );

    \I__10254\ : InMux
    port map (
            O => \N__44626\,
            I => \N__44494\
        );

    \I__10253\ : InMux
    port map (
            O => \N__44625\,
            I => \N__44494\
        );

    \I__10252\ : InMux
    port map (
            O => \N__44624\,
            I => \N__44494\
        );

    \I__10251\ : InMux
    port map (
            O => \N__44623\,
            I => \N__44494\
        );

    \I__10250\ : InMux
    port map (
            O => \N__44622\,
            I => \N__44494\
        );

    \I__10249\ : Span4Mux_h
    port map (
            O => \N__44619\,
            I => \N__44485\
        );

    \I__10248\ : Span4Mux_v
    port map (
            O => \N__44612\,
            I => \N__44485\
        );

    \I__10247\ : LocalMux
    port map (
            O => \N__44597\,
            I => \N__44485\
        );

    \I__10246\ : LocalMux
    port map (
            O => \N__44580\,
            I => \N__44485\
        );

    \I__10245\ : InMux
    port map (
            O => \N__44577\,
            I => \N__44468\
        );

    \I__10244\ : InMux
    port map (
            O => \N__44576\,
            I => \N__44468\
        );

    \I__10243\ : InMux
    port map (
            O => \N__44573\,
            I => \N__44468\
        );

    \I__10242\ : InMux
    port map (
            O => \N__44572\,
            I => \N__44468\
        );

    \I__10241\ : InMux
    port map (
            O => \N__44569\,
            I => \N__44468\
        );

    \I__10240\ : InMux
    port map (
            O => \N__44568\,
            I => \N__44468\
        );

    \I__10239\ : InMux
    port map (
            O => \N__44565\,
            I => \N__44468\
        );

    \I__10238\ : InMux
    port map (
            O => \N__44564\,
            I => \N__44468\
        );

    \I__10237\ : InMux
    port map (
            O => \N__44561\,
            I => \N__44455\
        );

    \I__10236\ : InMux
    port map (
            O => \N__44560\,
            I => \N__44455\
        );

    \I__10235\ : InMux
    port map (
            O => \N__44557\,
            I => \N__44455\
        );

    \I__10234\ : InMux
    port map (
            O => \N__44556\,
            I => \N__44455\
        );

    \I__10233\ : InMux
    port map (
            O => \N__44553\,
            I => \N__44455\
        );

    \I__10232\ : InMux
    port map (
            O => \N__44552\,
            I => \N__44455\
        );

    \I__10231\ : Span4Mux_v
    port map (
            O => \N__44545\,
            I => \N__44446\
        );

    \I__10230\ : Span4Mux_v
    port map (
            O => \N__44542\,
            I => \N__44446\
        );

    \I__10229\ : Span4Mux_h
    port map (
            O => \N__44539\,
            I => \N__44446\
        );

    \I__10228\ : Span4Mux_v
    port map (
            O => \N__44518\,
            I => \N__44446\
        );

    \I__10227\ : Odrv4
    port map (
            O => \N__44515\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10226\ : Odrv4
    port map (
            O => \N__44508\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10225\ : LocalMux
    port map (
            O => \N__44505\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10224\ : LocalMux
    port map (
            O => \N__44494\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10223\ : Odrv4
    port map (
            O => \N__44485\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10222\ : LocalMux
    port map (
            O => \N__44468\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10221\ : LocalMux
    port map (
            O => \N__44455\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10220\ : Odrv4
    port map (
            O => \N__44446\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10219\ : CascadeMux
    port map (
            O => \N__44429\,
            I => \N__44411\
        );

    \I__10218\ : CascadeMux
    port map (
            O => \N__44428\,
            I => \N__44408\
        );

    \I__10217\ : InMux
    port map (
            O => \N__44427\,
            I => \N__44385\
        );

    \I__10216\ : InMux
    port map (
            O => \N__44426\,
            I => \N__44382\
        );

    \I__10215\ : InMux
    port map (
            O => \N__44425\,
            I => \N__44369\
        );

    \I__10214\ : InMux
    port map (
            O => \N__44424\,
            I => \N__44369\
        );

    \I__10213\ : InMux
    port map (
            O => \N__44423\,
            I => \N__44369\
        );

    \I__10212\ : InMux
    port map (
            O => \N__44422\,
            I => \N__44369\
        );

    \I__10211\ : InMux
    port map (
            O => \N__44421\,
            I => \N__44369\
        );

    \I__10210\ : InMux
    port map (
            O => \N__44420\,
            I => \N__44369\
        );

    \I__10209\ : CascadeMux
    port map (
            O => \N__44419\,
            I => \N__44366\
        );

    \I__10208\ : InMux
    port map (
            O => \N__44418\,
            I => \N__44356\
        );

    \I__10207\ : InMux
    port map (
            O => \N__44417\,
            I => \N__44352\
        );

    \I__10206\ : CascadeMux
    port map (
            O => \N__44416\,
            I => \N__44349\
        );

    \I__10205\ : InMux
    port map (
            O => \N__44415\,
            I => \N__44344\
        );

    \I__10204\ : InMux
    port map (
            O => \N__44414\,
            I => \N__44344\
        );

    \I__10203\ : InMux
    port map (
            O => \N__44411\,
            I => \N__44339\
        );

    \I__10202\ : InMux
    port map (
            O => \N__44408\,
            I => \N__44339\
        );

    \I__10201\ : InMux
    port map (
            O => \N__44407\,
            I => \N__44336\
        );

    \I__10200\ : InMux
    port map (
            O => \N__44406\,
            I => \N__44323\
        );

    \I__10199\ : InMux
    port map (
            O => \N__44405\,
            I => \N__44323\
        );

    \I__10198\ : InMux
    port map (
            O => \N__44404\,
            I => \N__44323\
        );

    \I__10197\ : InMux
    port map (
            O => \N__44403\,
            I => \N__44323\
        );

    \I__10196\ : InMux
    port map (
            O => \N__44402\,
            I => \N__44323\
        );

    \I__10195\ : InMux
    port map (
            O => \N__44401\,
            I => \N__44323\
        );

    \I__10194\ : InMux
    port map (
            O => \N__44400\,
            I => \N__44316\
        );

    \I__10193\ : InMux
    port map (
            O => \N__44399\,
            I => \N__44316\
        );

    \I__10192\ : InMux
    port map (
            O => \N__44398\,
            I => \N__44316\
        );

    \I__10191\ : InMux
    port map (
            O => \N__44397\,
            I => \N__44311\
        );

    \I__10190\ : InMux
    port map (
            O => \N__44396\,
            I => \N__44311\
        );

    \I__10189\ : InMux
    port map (
            O => \N__44395\,
            I => \N__44302\
        );

    \I__10188\ : InMux
    port map (
            O => \N__44394\,
            I => \N__44302\
        );

    \I__10187\ : InMux
    port map (
            O => \N__44393\,
            I => \N__44302\
        );

    \I__10186\ : InMux
    port map (
            O => \N__44392\,
            I => \N__44302\
        );

    \I__10185\ : InMux
    port map (
            O => \N__44391\,
            I => \N__44299\
        );

    \I__10184\ : InMux
    port map (
            O => \N__44390\,
            I => \N__44288\
        );

    \I__10183\ : InMux
    port map (
            O => \N__44389\,
            I => \N__44283\
        );

    \I__10182\ : InMux
    port map (
            O => \N__44388\,
            I => \N__44283\
        );

    \I__10181\ : LocalMux
    port map (
            O => \N__44385\,
            I => \N__44272\
        );

    \I__10180\ : LocalMux
    port map (
            O => \N__44382\,
            I => \N__44272\
        );

    \I__10179\ : LocalMux
    port map (
            O => \N__44369\,
            I => \N__44269\
        );

    \I__10178\ : InMux
    port map (
            O => \N__44366\,
            I => \N__44252\
        );

    \I__10177\ : InMux
    port map (
            O => \N__44365\,
            I => \N__44252\
        );

    \I__10176\ : InMux
    port map (
            O => \N__44364\,
            I => \N__44252\
        );

    \I__10175\ : InMux
    port map (
            O => \N__44363\,
            I => \N__44252\
        );

    \I__10174\ : InMux
    port map (
            O => \N__44362\,
            I => \N__44252\
        );

    \I__10173\ : InMux
    port map (
            O => \N__44361\,
            I => \N__44252\
        );

    \I__10172\ : InMux
    port map (
            O => \N__44360\,
            I => \N__44252\
        );

    \I__10171\ : InMux
    port map (
            O => \N__44359\,
            I => \N__44252\
        );

    \I__10170\ : LocalMux
    port map (
            O => \N__44356\,
            I => \N__44249\
        );

    \I__10169\ : InMux
    port map (
            O => \N__44355\,
            I => \N__44246\
        );

    \I__10168\ : LocalMux
    port map (
            O => \N__44352\,
            I => \N__44243\
        );

    \I__10167\ : InMux
    port map (
            O => \N__44349\,
            I => \N__44240\
        );

    \I__10166\ : LocalMux
    port map (
            O => \N__44344\,
            I => \N__44236\
        );

    \I__10165\ : LocalMux
    port map (
            O => \N__44339\,
            I => \N__44227\
        );

    \I__10164\ : LocalMux
    port map (
            O => \N__44336\,
            I => \N__44227\
        );

    \I__10163\ : LocalMux
    port map (
            O => \N__44323\,
            I => \N__44227\
        );

    \I__10162\ : LocalMux
    port map (
            O => \N__44316\,
            I => \N__44227\
        );

    \I__10161\ : LocalMux
    port map (
            O => \N__44311\,
            I => \N__44222\
        );

    \I__10160\ : LocalMux
    port map (
            O => \N__44302\,
            I => \N__44222\
        );

    \I__10159\ : LocalMux
    port map (
            O => \N__44299\,
            I => \N__44219\
        );

    \I__10158\ : InMux
    port map (
            O => \N__44298\,
            I => \N__44216\
        );

    \I__10157\ : InMux
    port map (
            O => \N__44297\,
            I => \N__44201\
        );

    \I__10156\ : InMux
    port map (
            O => \N__44296\,
            I => \N__44201\
        );

    \I__10155\ : InMux
    port map (
            O => \N__44295\,
            I => \N__44201\
        );

    \I__10154\ : InMux
    port map (
            O => \N__44294\,
            I => \N__44201\
        );

    \I__10153\ : InMux
    port map (
            O => \N__44293\,
            I => \N__44201\
        );

    \I__10152\ : InMux
    port map (
            O => \N__44292\,
            I => \N__44201\
        );

    \I__10151\ : InMux
    port map (
            O => \N__44291\,
            I => \N__44201\
        );

    \I__10150\ : LocalMux
    port map (
            O => \N__44288\,
            I => \N__44184\
        );

    \I__10149\ : LocalMux
    port map (
            O => \N__44283\,
            I => \N__44184\
        );

    \I__10148\ : InMux
    port map (
            O => \N__44282\,
            I => \N__44171\
        );

    \I__10147\ : InMux
    port map (
            O => \N__44281\,
            I => \N__44171\
        );

    \I__10146\ : InMux
    port map (
            O => \N__44280\,
            I => \N__44171\
        );

    \I__10145\ : InMux
    port map (
            O => \N__44279\,
            I => \N__44171\
        );

    \I__10144\ : InMux
    port map (
            O => \N__44278\,
            I => \N__44171\
        );

    \I__10143\ : InMux
    port map (
            O => \N__44277\,
            I => \N__44171\
        );

    \I__10142\ : Span4Mux_v
    port map (
            O => \N__44272\,
            I => \N__44162\
        );

    \I__10141\ : Span4Mux_v
    port map (
            O => \N__44269\,
            I => \N__44162\
        );

    \I__10140\ : LocalMux
    port map (
            O => \N__44252\,
            I => \N__44162\
        );

    \I__10139\ : Span4Mux_h
    port map (
            O => \N__44249\,
            I => \N__44162\
        );

    \I__10138\ : LocalMux
    port map (
            O => \N__44246\,
            I => \N__44155\
        );

    \I__10137\ : Span4Mux_h
    port map (
            O => \N__44243\,
            I => \N__44155\
        );

    \I__10136\ : LocalMux
    port map (
            O => \N__44240\,
            I => \N__44155\
        );

    \I__10135\ : InMux
    port map (
            O => \N__44239\,
            I => \N__44152\
        );

    \I__10134\ : Span4Mux_v
    port map (
            O => \N__44236\,
            I => \N__44145\
        );

    \I__10133\ : Span4Mux_v
    port map (
            O => \N__44227\,
            I => \N__44145\
        );

    \I__10132\ : Span4Mux_v
    port map (
            O => \N__44222\,
            I => \N__44145\
        );

    \I__10131\ : Span4Mux_v
    port map (
            O => \N__44219\,
            I => \N__44138\
        );

    \I__10130\ : LocalMux
    port map (
            O => \N__44216\,
            I => \N__44138\
        );

    \I__10129\ : LocalMux
    port map (
            O => \N__44201\,
            I => \N__44138\
        );

    \I__10128\ : InMux
    port map (
            O => \N__44200\,
            I => \N__44123\
        );

    \I__10127\ : InMux
    port map (
            O => \N__44199\,
            I => \N__44123\
        );

    \I__10126\ : InMux
    port map (
            O => \N__44198\,
            I => \N__44123\
        );

    \I__10125\ : InMux
    port map (
            O => \N__44197\,
            I => \N__44123\
        );

    \I__10124\ : InMux
    port map (
            O => \N__44196\,
            I => \N__44123\
        );

    \I__10123\ : InMux
    port map (
            O => \N__44195\,
            I => \N__44123\
        );

    \I__10122\ : InMux
    port map (
            O => \N__44194\,
            I => \N__44123\
        );

    \I__10121\ : InMux
    port map (
            O => \N__44193\,
            I => \N__44118\
        );

    \I__10120\ : InMux
    port map (
            O => \N__44192\,
            I => \N__44118\
        );

    \I__10119\ : InMux
    port map (
            O => \N__44191\,
            I => \N__44115\
        );

    \I__10118\ : InMux
    port map (
            O => \N__44190\,
            I => \N__44110\
        );

    \I__10117\ : InMux
    port map (
            O => \N__44189\,
            I => \N__44110\
        );

    \I__10116\ : Span4Mux_v
    port map (
            O => \N__44184\,
            I => \N__44105\
        );

    \I__10115\ : LocalMux
    port map (
            O => \N__44171\,
            I => \N__44105\
        );

    \I__10114\ : Span4Mux_h
    port map (
            O => \N__44162\,
            I => \N__44102\
        );

    \I__10113\ : Span4Mux_v
    port map (
            O => \N__44155\,
            I => \N__44095\
        );

    \I__10112\ : LocalMux
    port map (
            O => \N__44152\,
            I => \N__44095\
        );

    \I__10111\ : Span4Mux_h
    port map (
            O => \N__44145\,
            I => \N__44095\
        );

    \I__10110\ : Odrv4
    port map (
            O => \N__44138\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10109\ : LocalMux
    port map (
            O => \N__44123\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10108\ : LocalMux
    port map (
            O => \N__44118\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10107\ : LocalMux
    port map (
            O => \N__44115\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10106\ : LocalMux
    port map (
            O => \N__44110\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10105\ : Odrv4
    port map (
            O => \N__44105\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10104\ : Odrv4
    port map (
            O => \N__44102\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10103\ : Odrv4
    port map (
            O => \N__44095\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10102\ : CascadeMux
    port map (
            O => \N__44078\,
            I => \N__44075\
        );

    \I__10101\ : InMux
    port map (
            O => \N__44075\,
            I => \N__44072\
        );

    \I__10100\ : LocalMux
    port map (
            O => \N__44072\,
            I => \N__44069\
        );

    \I__10099\ : Span4Mux_h
    port map (
            O => \N__44069\,
            I => \N__44066\
        );

    \I__10098\ : Odrv4
    port map (
            O => \N__44066\,
            I => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\
        );

    \I__10097\ : InMux
    port map (
            O => \N__44063\,
            I => \N__44058\
        );

    \I__10096\ : InMux
    port map (
            O => \N__44062\,
            I => \N__44055\
        );

    \I__10095\ : InMux
    port map (
            O => \N__44061\,
            I => \N__44052\
        );

    \I__10094\ : LocalMux
    port map (
            O => \N__44058\,
            I => \N__44047\
        );

    \I__10093\ : LocalMux
    port map (
            O => \N__44055\,
            I => \N__44047\
        );

    \I__10092\ : LocalMux
    port map (
            O => \N__44052\,
            I => \N__44043\
        );

    \I__10091\ : Span4Mux_h
    port map (
            O => \N__44047\,
            I => \N__44040\
        );

    \I__10090\ : InMux
    port map (
            O => \N__44046\,
            I => \N__44037\
        );

    \I__10089\ : Span4Mux_v
    port map (
            O => \N__44043\,
            I => \N__44034\
        );

    \I__10088\ : Span4Mux_v
    port map (
            O => \N__44040\,
            I => \N__44029\
        );

    \I__10087\ : LocalMux
    port map (
            O => \N__44037\,
            I => \N__44029\
        );

    \I__10086\ : Odrv4
    port map (
            O => \N__44034\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__10085\ : Odrv4
    port map (
            O => \N__44029\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__10084\ : InMux
    port map (
            O => \N__44024\,
            I => \N__44021\
        );

    \I__10083\ : LocalMux
    port map (
            O => \N__44021\,
            I => \N__44018\
        );

    \I__10082\ : Span4Mux_h
    port map (
            O => \N__44018\,
            I => \N__44015\
        );

    \I__10081\ : Odrv4
    port map (
            O => \N__44015\,
            I => \current_shift_inst.un4_control_input_1_axb_14\
        );

    \I__10080\ : InMux
    port map (
            O => \N__44012\,
            I => \N__44009\
        );

    \I__10079\ : LocalMux
    port map (
            O => \N__44009\,
            I => \N__44004\
        );

    \I__10078\ : InMux
    port map (
            O => \N__44008\,
            I => \N__44001\
        );

    \I__10077\ : InMux
    port map (
            O => \N__44007\,
            I => \N__43998\
        );

    \I__10076\ : Span4Mux_h
    port map (
            O => \N__44004\,
            I => \N__43990\
        );

    \I__10075\ : LocalMux
    port map (
            O => \N__44001\,
            I => \N__43990\
        );

    \I__10074\ : LocalMux
    port map (
            O => \N__43998\,
            I => \N__43990\
        );

    \I__10073\ : InMux
    port map (
            O => \N__43997\,
            I => \N__43987\
        );

    \I__10072\ : Span4Mux_h
    port map (
            O => \N__43990\,
            I => \N__43982\
        );

    \I__10071\ : LocalMux
    port map (
            O => \N__43987\,
            I => \N__43982\
        );

    \I__10070\ : Span4Mux_v
    port map (
            O => \N__43982\,
            I => \N__43979\
        );

    \I__10069\ : Odrv4
    port map (
            O => \N__43979\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__10068\ : InMux
    port map (
            O => \N__43976\,
            I => \N__43973\
        );

    \I__10067\ : LocalMux
    port map (
            O => \N__43973\,
            I => \N__43970\
        );

    \I__10066\ : Odrv4
    port map (
            O => \N__43970\,
            I => \current_shift_inst.un4_control_input_1_axb_29\
        );

    \I__10065\ : CascadeMux
    port map (
            O => \N__43967\,
            I => \N__43963\
        );

    \I__10064\ : CascadeMux
    port map (
            O => \N__43966\,
            I => \N__43960\
        );

    \I__10063\ : InMux
    port map (
            O => \N__43963\,
            I => \N__43956\
        );

    \I__10062\ : InMux
    port map (
            O => \N__43960\,
            I => \N__43953\
        );

    \I__10061\ : InMux
    port map (
            O => \N__43959\,
            I => \N__43950\
        );

    \I__10060\ : LocalMux
    port map (
            O => \N__43956\,
            I => \N__43946\
        );

    \I__10059\ : LocalMux
    port map (
            O => \N__43953\,
            I => \N__43943\
        );

    \I__10058\ : LocalMux
    port map (
            O => \N__43950\,
            I => \N__43940\
        );

    \I__10057\ : InMux
    port map (
            O => \N__43949\,
            I => \N__43937\
        );

    \I__10056\ : Span4Mux_h
    port map (
            O => \N__43946\,
            I => \N__43934\
        );

    \I__10055\ : Span4Mux_v
    port map (
            O => \N__43943\,
            I => \N__43931\
        );

    \I__10054\ : Span4Mux_h
    port map (
            O => \N__43940\,
            I => \N__43928\
        );

    \I__10053\ : LocalMux
    port map (
            O => \N__43937\,
            I => \N__43925\
        );

    \I__10052\ : Odrv4
    port map (
            O => \N__43934\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__10051\ : Odrv4
    port map (
            O => \N__43931\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__10050\ : Odrv4
    port map (
            O => \N__43928\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__10049\ : Odrv12
    port map (
            O => \N__43925\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__10048\ : InMux
    port map (
            O => \N__43916\,
            I => \N__43913\
        );

    \I__10047\ : LocalMux
    port map (
            O => \N__43913\,
            I => \N__43910\
        );

    \I__10046\ : Odrv12
    port map (
            O => \N__43910\,
            I => \current_shift_inst.un4_control_input_1_axb_17\
        );

    \I__10045\ : CascadeMux
    port map (
            O => \N__43907\,
            I => \N__43904\
        );

    \I__10044\ : InMux
    port map (
            O => \N__43904\,
            I => \N__43901\
        );

    \I__10043\ : LocalMux
    port map (
            O => \N__43901\,
            I => \N__43896\
        );

    \I__10042\ : InMux
    port map (
            O => \N__43900\,
            I => \N__43891\
        );

    \I__10041\ : InMux
    port map (
            O => \N__43899\,
            I => \N__43891\
        );

    \I__10040\ : Span4Mux_h
    port map (
            O => \N__43896\,
            I => \N__43885\
        );

    \I__10039\ : LocalMux
    port map (
            O => \N__43891\,
            I => \N__43885\
        );

    \I__10038\ : InMux
    port map (
            O => \N__43890\,
            I => \N__43882\
        );

    \I__10037\ : Span4Mux_h
    port map (
            O => \N__43885\,
            I => \N__43879\
        );

    \I__10036\ : LocalMux
    port map (
            O => \N__43882\,
            I => \N__43876\
        );

    \I__10035\ : Odrv4
    port map (
            O => \N__43879\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__10034\ : Odrv4
    port map (
            O => \N__43876\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__10033\ : InMux
    port map (
            O => \N__43871\,
            I => \N__43868\
        );

    \I__10032\ : LocalMux
    port map (
            O => \N__43868\,
            I => \N__43865\
        );

    \I__10031\ : Odrv12
    port map (
            O => \N__43865\,
            I => \current_shift_inst.un4_control_input_1_axb_19\
        );

    \I__10030\ : InMux
    port map (
            O => \N__43862\,
            I => \N__43859\
        );

    \I__10029\ : LocalMux
    port map (
            O => \N__43859\,
            I => \N__43856\
        );

    \I__10028\ : Span4Mux_v
    port map (
            O => \N__43856\,
            I => \N__43852\
        );

    \I__10027\ : CascadeMux
    port map (
            O => \N__43855\,
            I => \N__43848\
        );

    \I__10026\ : Span4Mux_h
    port map (
            O => \N__43852\,
            I => \N__43840\
        );

    \I__10025\ : InMux
    port map (
            O => \N__43851\,
            I => \N__43837\
        );

    \I__10024\ : InMux
    port map (
            O => \N__43848\,
            I => \N__43830\
        );

    \I__10023\ : InMux
    port map (
            O => \N__43847\,
            I => \N__43830\
        );

    \I__10022\ : InMux
    port map (
            O => \N__43846\,
            I => \N__43830\
        );

    \I__10021\ : InMux
    port map (
            O => \N__43845\,
            I => \N__43827\
        );

    \I__10020\ : InMux
    port map (
            O => \N__43844\,
            I => \N__43822\
        );

    \I__10019\ : InMux
    port map (
            O => \N__43843\,
            I => \N__43822\
        );

    \I__10018\ : Span4Mux_h
    port map (
            O => \N__43840\,
            I => \N__43818\
        );

    \I__10017\ : LocalMux
    port map (
            O => \N__43837\,
            I => \N__43811\
        );

    \I__10016\ : LocalMux
    port map (
            O => \N__43830\,
            I => \N__43811\
        );

    \I__10015\ : LocalMux
    port map (
            O => \N__43827\,
            I => \N__43811\
        );

    \I__10014\ : LocalMux
    port map (
            O => \N__43822\,
            I => \N__43808\
        );

    \I__10013\ : InMux
    port map (
            O => \N__43821\,
            I => \N__43805\
        );

    \I__10012\ : Span4Mux_h
    port map (
            O => \N__43818\,
            I => \N__43799\
        );

    \I__10011\ : Span4Mux_v
    port map (
            O => \N__43811\,
            I => \N__43799\
        );

    \I__10010\ : Span4Mux_h
    port map (
            O => \N__43808\,
            I => \N__43796\
        );

    \I__10009\ : LocalMux
    port map (
            O => \N__43805\,
            I => \N__43793\
        );

    \I__10008\ : InMux
    port map (
            O => \N__43804\,
            I => \N__43790\
        );

    \I__10007\ : Odrv4
    port map (
            O => \N__43799\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__10006\ : Odrv4
    port map (
            O => \N__43796\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__10005\ : Odrv4
    port map (
            O => \N__43793\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__10004\ : LocalMux
    port map (
            O => \N__43790\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__10003\ : CascadeMux
    port map (
            O => \N__43781\,
            I => \N__43778\
        );

    \I__10002\ : InMux
    port map (
            O => \N__43778\,
            I => \N__43775\
        );

    \I__10001\ : LocalMux
    port map (
            O => \N__43775\,
            I => \N__43772\
        );

    \I__10000\ : Span4Mux_h
    port map (
            O => \N__43772\,
            I => \N__43769\
        );

    \I__9999\ : Odrv4
    port map (
            O => \N__43769\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt24\
        );

    \I__9998\ : InMux
    port map (
            O => \N__43766\,
            I => \N__43763\
        );

    \I__9997\ : LocalMux
    port map (
            O => \N__43763\,
            I => \N__43760\
        );

    \I__9996\ : Span12Mux_v
    port map (
            O => \N__43760\,
            I => \N__43757\
        );

    \I__9995\ : Odrv12
    port map (
            O => \N__43757\,
            I => \current_shift_inst.un4_control_input_1_axb_28\
        );

    \I__9994\ : CascadeMux
    port map (
            O => \N__43754\,
            I => \N__43751\
        );

    \I__9993\ : InMux
    port map (
            O => \N__43751\,
            I => \N__43747\
        );

    \I__9992\ : CascadeMux
    port map (
            O => \N__43750\,
            I => \N__43744\
        );

    \I__9991\ : LocalMux
    port map (
            O => \N__43747\,
            I => \N__43740\
        );

    \I__9990\ : InMux
    port map (
            O => \N__43744\,
            I => \N__43735\
        );

    \I__9989\ : InMux
    port map (
            O => \N__43743\,
            I => \N__43735\
        );

    \I__9988\ : Odrv4
    port map (
            O => \N__43740\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__9987\ : LocalMux
    port map (
            O => \N__43735\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__9986\ : InMux
    port map (
            O => \N__43730\,
            I => \current_shift_inst.un4_control_input_1_cry_27\
        );

    \I__9985\ : CascadeMux
    port map (
            O => \N__43727\,
            I => \N__43723\
        );

    \I__9984\ : InMux
    port map (
            O => \N__43726\,
            I => \N__43720\
        );

    \I__9983\ : InMux
    port map (
            O => \N__43723\,
            I => \N__43717\
        );

    \I__9982\ : LocalMux
    port map (
            O => \N__43720\,
            I => \N__43711\
        );

    \I__9981\ : LocalMux
    port map (
            O => \N__43717\,
            I => \N__43711\
        );

    \I__9980\ : InMux
    port map (
            O => \N__43716\,
            I => \N__43708\
        );

    \I__9979\ : Odrv12
    port map (
            O => \N__43711\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__9978\ : LocalMux
    port map (
            O => \N__43708\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__9977\ : InMux
    port map (
            O => \N__43703\,
            I => \current_shift_inst.un4_control_input_1_cry_28\
        );

    \I__9976\ : InMux
    port map (
            O => \N__43700\,
            I => \current_shift_inst.un4_control_input1_31\
        );

    \I__9975\ : CascadeMux
    port map (
            O => \N__43697\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO_cascade_\
        );

    \I__9974\ : InMux
    port map (
            O => \N__43694\,
            I => \N__43691\
        );

    \I__9973\ : LocalMux
    port map (
            O => \N__43691\,
            I => \N__43688\
        );

    \I__9972\ : Odrv4
    port map (
            O => \N__43688\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\
        );

    \I__9971\ : InMux
    port map (
            O => \N__43685\,
            I => \N__43681\
        );

    \I__9970\ : InMux
    port map (
            O => \N__43684\,
            I => \N__43676\
        );

    \I__9969\ : LocalMux
    port map (
            O => \N__43681\,
            I => \N__43673\
        );

    \I__9968\ : InMux
    port map (
            O => \N__43680\,
            I => \N__43668\
        );

    \I__9967\ : InMux
    port map (
            O => \N__43679\,
            I => \N__43668\
        );

    \I__9966\ : LocalMux
    port map (
            O => \N__43676\,
            I => \N__43665\
        );

    \I__9965\ : Span4Mux_h
    port map (
            O => \N__43673\,
            I => \N__43660\
        );

    \I__9964\ : LocalMux
    port map (
            O => \N__43668\,
            I => \N__43660\
        );

    \I__9963\ : Span4Mux_h
    port map (
            O => \N__43665\,
            I => \N__43657\
        );

    \I__9962\ : Span4Mux_v
    port map (
            O => \N__43660\,
            I => \N__43654\
        );

    \I__9961\ : Odrv4
    port map (
            O => \N__43657\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__9960\ : Odrv4
    port map (
            O => \N__43654\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__9959\ : InMux
    port map (
            O => \N__43649\,
            I => \N__43646\
        );

    \I__9958\ : LocalMux
    port map (
            O => \N__43646\,
            I => \N__43641\
        );

    \I__9957\ : InMux
    port map (
            O => \N__43645\,
            I => \N__43638\
        );

    \I__9956\ : InMux
    port map (
            O => \N__43644\,
            I => \N__43635\
        );

    \I__9955\ : Odrv4
    port map (
            O => \N__43641\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__9954\ : LocalMux
    port map (
            O => \N__43638\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__9953\ : LocalMux
    port map (
            O => \N__43635\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__9952\ : CascadeMux
    port map (
            O => \N__43628\,
            I => \N__43625\
        );

    \I__9951\ : InMux
    port map (
            O => \N__43625\,
            I => \N__43622\
        );

    \I__9950\ : LocalMux
    port map (
            O => \N__43622\,
            I => \N__43619\
        );

    \I__9949\ : Span4Mux_h
    port map (
            O => \N__43619\,
            I => \N__43616\
        );

    \I__9948\ : Span4Mux_v
    port map (
            O => \N__43616\,
            I => \N__43613\
        );

    \I__9947\ : Odrv4
    port map (
            O => \N__43613\,
            I => \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0\
        );

    \I__9946\ : CascadeMux
    port map (
            O => \N__43610\,
            I => \N__43607\
        );

    \I__9945\ : InMux
    port map (
            O => \N__43607\,
            I => \N__43604\
        );

    \I__9944\ : LocalMux
    port map (
            O => \N__43604\,
            I => \N__43601\
        );

    \I__9943\ : Span12Mux_v
    port map (
            O => \N__43601\,
            I => \N__43598\
        );

    \I__9942\ : Odrv12
    port map (
            O => \N__43598\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2\
        );

    \I__9941\ : InMux
    port map (
            O => \N__43595\,
            I => \N__43590\
        );

    \I__9940\ : InMux
    port map (
            O => \N__43594\,
            I => \N__43587\
        );

    \I__9939\ : InMux
    port map (
            O => \N__43593\,
            I => \N__43584\
        );

    \I__9938\ : LocalMux
    port map (
            O => \N__43590\,
            I => \N__43581\
        );

    \I__9937\ : LocalMux
    port map (
            O => \N__43587\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__9936\ : LocalMux
    port map (
            O => \N__43584\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__9935\ : Odrv4
    port map (
            O => \N__43581\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__9934\ : CEMux
    port map (
            O => \N__43574\,
            I => \N__43550\
        );

    \I__9933\ : CEMux
    port map (
            O => \N__43573\,
            I => \N__43550\
        );

    \I__9932\ : CEMux
    port map (
            O => \N__43572\,
            I => \N__43550\
        );

    \I__9931\ : CEMux
    port map (
            O => \N__43571\,
            I => \N__43550\
        );

    \I__9930\ : CEMux
    port map (
            O => \N__43570\,
            I => \N__43550\
        );

    \I__9929\ : CEMux
    port map (
            O => \N__43569\,
            I => \N__43550\
        );

    \I__9928\ : CEMux
    port map (
            O => \N__43568\,
            I => \N__43550\
        );

    \I__9927\ : CEMux
    port map (
            O => \N__43567\,
            I => \N__43550\
        );

    \I__9926\ : GlobalMux
    port map (
            O => \N__43550\,
            I => \N__43547\
        );

    \I__9925\ : gio2CtrlBuf
    port map (
            O => \N__43547\,
            I => \current_shift_inst.timer_s1.N_162_i_g\
        );

    \I__9924\ : InMux
    port map (
            O => \N__43544\,
            I => \N__43541\
        );

    \I__9923\ : LocalMux
    port map (
            O => \N__43541\,
            I => \N__43538\
        );

    \I__9922\ : Span4Mux_h
    port map (
            O => \N__43538\,
            I => \N__43535\
        );

    \I__9921\ : Odrv4
    port map (
            O => \N__43535\,
            I => \current_shift_inst.un4_control_input_1_axb_1\
        );

    \I__9920\ : InMux
    port map (
            O => \N__43532\,
            I => \N__43529\
        );

    \I__9919\ : LocalMux
    port map (
            O => \N__43529\,
            I => \N__43526\
        );

    \I__9918\ : Span4Mux_h
    port map (
            O => \N__43526\,
            I => \N__43523\
        );

    \I__9917\ : Odrv4
    port map (
            O => \N__43523\,
            I => \current_shift_inst.un4_control_input_1_axb_20\
        );

    \I__9916\ : CascadeMux
    port map (
            O => \N__43520\,
            I => \N__43517\
        );

    \I__9915\ : InMux
    port map (
            O => \N__43517\,
            I => \N__43513\
        );

    \I__9914\ : InMux
    port map (
            O => \N__43516\,
            I => \N__43510\
        );

    \I__9913\ : LocalMux
    port map (
            O => \N__43513\,
            I => \N__43507\
        );

    \I__9912\ : LocalMux
    port map (
            O => \N__43510\,
            I => \N__43501\
        );

    \I__9911\ : Span4Mux_h
    port map (
            O => \N__43507\,
            I => \N__43501\
        );

    \I__9910\ : InMux
    port map (
            O => \N__43506\,
            I => \N__43498\
        );

    \I__9909\ : Odrv4
    port map (
            O => \N__43501\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__9908\ : LocalMux
    port map (
            O => \N__43498\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__9907\ : InMux
    port map (
            O => \N__43493\,
            I => \current_shift_inst.un4_control_input_1_cry_19\
        );

    \I__9906\ : InMux
    port map (
            O => \N__43490\,
            I => \N__43487\
        );

    \I__9905\ : LocalMux
    port map (
            O => \N__43487\,
            I => \N__43484\
        );

    \I__9904\ : Span4Mux_v
    port map (
            O => \N__43484\,
            I => \N__43481\
        );

    \I__9903\ : Odrv4
    port map (
            O => \N__43481\,
            I => \current_shift_inst.un4_control_input_1_axb_21\
        );

    \I__9902\ : InMux
    port map (
            O => \N__43478\,
            I => \N__43475\
        );

    \I__9901\ : LocalMux
    port map (
            O => \N__43475\,
            I => \N__43470\
        );

    \I__9900\ : InMux
    port map (
            O => \N__43474\,
            I => \N__43467\
        );

    \I__9899\ : InMux
    port map (
            O => \N__43473\,
            I => \N__43464\
        );

    \I__9898\ : Odrv4
    port map (
            O => \N__43470\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__9897\ : LocalMux
    port map (
            O => \N__43467\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__9896\ : LocalMux
    port map (
            O => \N__43464\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__9895\ : InMux
    port map (
            O => \N__43457\,
            I => \current_shift_inst.un4_control_input_1_cry_20\
        );

    \I__9894\ : InMux
    port map (
            O => \N__43454\,
            I => \N__43451\
        );

    \I__9893\ : LocalMux
    port map (
            O => \N__43451\,
            I => \N__43448\
        );

    \I__9892\ : Span4Mux_h
    port map (
            O => \N__43448\,
            I => \N__43445\
        );

    \I__9891\ : Odrv4
    port map (
            O => \N__43445\,
            I => \current_shift_inst.un4_control_input_1_axb_22\
        );

    \I__9890\ : CascadeMux
    port map (
            O => \N__43442\,
            I => \N__43438\
        );

    \I__9889\ : InMux
    port map (
            O => \N__43441\,
            I => \N__43435\
        );

    \I__9888\ : InMux
    port map (
            O => \N__43438\,
            I => \N__43432\
        );

    \I__9887\ : LocalMux
    port map (
            O => \N__43435\,
            I => \N__43429\
        );

    \I__9886\ : LocalMux
    port map (
            O => \N__43432\,
            I => \N__43424\
        );

    \I__9885\ : Span4Mux_v
    port map (
            O => \N__43429\,
            I => \N__43424\
        );

    \I__9884\ : Sp12to4
    port map (
            O => \N__43424\,
            I => \N__43420\
        );

    \I__9883\ : InMux
    port map (
            O => \N__43423\,
            I => \N__43417\
        );

    \I__9882\ : Odrv12
    port map (
            O => \N__43420\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__9881\ : LocalMux
    port map (
            O => \N__43417\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__9880\ : InMux
    port map (
            O => \N__43412\,
            I => \current_shift_inst.un4_control_input_1_cry_21\
        );

    \I__9879\ : InMux
    port map (
            O => \N__43409\,
            I => \N__43406\
        );

    \I__9878\ : LocalMux
    port map (
            O => \N__43406\,
            I => \N__43403\
        );

    \I__9877\ : Span4Mux_h
    port map (
            O => \N__43403\,
            I => \N__43400\
        );

    \I__9876\ : Odrv4
    port map (
            O => \N__43400\,
            I => \current_shift_inst.un4_control_input_1_axb_23\
        );

    \I__9875\ : CascadeMux
    port map (
            O => \N__43397\,
            I => \N__43393\
        );

    \I__9874\ : InMux
    port map (
            O => \N__43396\,
            I => \N__43389\
        );

    \I__9873\ : InMux
    port map (
            O => \N__43393\,
            I => \N__43386\
        );

    \I__9872\ : InMux
    port map (
            O => \N__43392\,
            I => \N__43383\
        );

    \I__9871\ : LocalMux
    port map (
            O => \N__43389\,
            I => \N__43378\
        );

    \I__9870\ : LocalMux
    port map (
            O => \N__43386\,
            I => \N__43378\
        );

    \I__9869\ : LocalMux
    port map (
            O => \N__43383\,
            I => \N__43375\
        );

    \I__9868\ : Odrv12
    port map (
            O => \N__43378\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__9867\ : Odrv4
    port map (
            O => \N__43375\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__9866\ : InMux
    port map (
            O => \N__43370\,
            I => \current_shift_inst.un4_control_input_1_cry_22\
        );

    \I__9865\ : InMux
    port map (
            O => \N__43367\,
            I => \N__43364\
        );

    \I__9864\ : LocalMux
    port map (
            O => \N__43364\,
            I => \N__43361\
        );

    \I__9863\ : Span12Mux_v
    port map (
            O => \N__43361\,
            I => \N__43358\
        );

    \I__9862\ : Odrv12
    port map (
            O => \N__43358\,
            I => \current_shift_inst.un4_control_input_1_axb_24\
        );

    \I__9861\ : InMux
    port map (
            O => \N__43355\,
            I => \N__43352\
        );

    \I__9860\ : LocalMux
    port map (
            O => \N__43352\,
            I => \N__43349\
        );

    \I__9859\ : Span4Mux_h
    port map (
            O => \N__43349\,
            I => \N__43345\
        );

    \I__9858\ : InMux
    port map (
            O => \N__43348\,
            I => \N__43342\
        );

    \I__9857\ : Span4Mux_h
    port map (
            O => \N__43345\,
            I => \N__43338\
        );

    \I__9856\ : LocalMux
    port map (
            O => \N__43342\,
            I => \N__43335\
        );

    \I__9855\ : InMux
    port map (
            O => \N__43341\,
            I => \N__43332\
        );

    \I__9854\ : Odrv4
    port map (
            O => \N__43338\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__9853\ : Odrv4
    port map (
            O => \N__43335\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__9852\ : LocalMux
    port map (
            O => \N__43332\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__9851\ : InMux
    port map (
            O => \N__43325\,
            I => \current_shift_inst.un4_control_input_1_cry_23\
        );

    \I__9850\ : InMux
    port map (
            O => \N__43322\,
            I => \N__43319\
        );

    \I__9849\ : LocalMux
    port map (
            O => \N__43319\,
            I => \N__43316\
        );

    \I__9848\ : Span4Mux_h
    port map (
            O => \N__43316\,
            I => \N__43313\
        );

    \I__9847\ : Odrv4
    port map (
            O => \N__43313\,
            I => \current_shift_inst.un4_control_input_1_axb_25\
        );

    \I__9846\ : CascadeMux
    port map (
            O => \N__43310\,
            I => \N__43306\
        );

    \I__9845\ : CascadeMux
    port map (
            O => \N__43309\,
            I => \N__43303\
        );

    \I__9844\ : InMux
    port map (
            O => \N__43306\,
            I => \N__43300\
        );

    \I__9843\ : InMux
    port map (
            O => \N__43303\,
            I => \N__43297\
        );

    \I__9842\ : LocalMux
    port map (
            O => \N__43300\,
            I => \N__43294\
        );

    \I__9841\ : LocalMux
    port map (
            O => \N__43297\,
            I => \N__43291\
        );

    \I__9840\ : Sp12to4
    port map (
            O => \N__43294\,
            I => \N__43285\
        );

    \I__9839\ : Span12Mux_h
    port map (
            O => \N__43291\,
            I => \N__43285\
        );

    \I__9838\ : InMux
    port map (
            O => \N__43290\,
            I => \N__43282\
        );

    \I__9837\ : Odrv12
    port map (
            O => \N__43285\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__9836\ : LocalMux
    port map (
            O => \N__43282\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__9835\ : InMux
    port map (
            O => \N__43277\,
            I => \bfn_18_17_0_\
        );

    \I__9834\ : InMux
    port map (
            O => \N__43274\,
            I => \N__43271\
        );

    \I__9833\ : LocalMux
    port map (
            O => \N__43271\,
            I => \N__43268\
        );

    \I__9832\ : Span4Mux_h
    port map (
            O => \N__43268\,
            I => \N__43265\
        );

    \I__9831\ : Odrv4
    port map (
            O => \N__43265\,
            I => \current_shift_inst.un4_control_input_1_axb_26\
        );

    \I__9830\ : InMux
    port map (
            O => \N__43262\,
            I => \N__43258\
        );

    \I__9829\ : InMux
    port map (
            O => \N__43261\,
            I => \N__43255\
        );

    \I__9828\ : LocalMux
    port map (
            O => \N__43258\,
            I => \N__43252\
        );

    \I__9827\ : LocalMux
    port map (
            O => \N__43255\,
            I => \N__43249\
        );

    \I__9826\ : Span4Mux_h
    port map (
            O => \N__43252\,
            I => \N__43245\
        );

    \I__9825\ : Span4Mux_v
    port map (
            O => \N__43249\,
            I => \N__43242\
        );

    \I__9824\ : InMux
    port map (
            O => \N__43248\,
            I => \N__43239\
        );

    \I__9823\ : Odrv4
    port map (
            O => \N__43245\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__9822\ : Odrv4
    port map (
            O => \N__43242\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__9821\ : LocalMux
    port map (
            O => \N__43239\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__9820\ : InMux
    port map (
            O => \N__43232\,
            I => \current_shift_inst.un4_control_input_1_cry_25\
        );

    \I__9819\ : InMux
    port map (
            O => \N__43229\,
            I => \N__43226\
        );

    \I__9818\ : LocalMux
    port map (
            O => \N__43226\,
            I => \N__43223\
        );

    \I__9817\ : Span4Mux_h
    port map (
            O => \N__43223\,
            I => \N__43220\
        );

    \I__9816\ : Odrv4
    port map (
            O => \N__43220\,
            I => \current_shift_inst.un4_control_input_1_axb_27\
        );

    \I__9815\ : InMux
    port map (
            O => \N__43217\,
            I => \N__43211\
        );

    \I__9814\ : InMux
    port map (
            O => \N__43216\,
            I => \N__43211\
        );

    \I__9813\ : LocalMux
    port map (
            O => \N__43211\,
            I => \N__43207\
        );

    \I__9812\ : InMux
    port map (
            O => \N__43210\,
            I => \N__43204\
        );

    \I__9811\ : Odrv4
    port map (
            O => \N__43207\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__9810\ : LocalMux
    port map (
            O => \N__43204\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__9809\ : InMux
    port map (
            O => \N__43199\,
            I => \current_shift_inst.un4_control_input_1_cry_26\
        );

    \I__9808\ : InMux
    port map (
            O => \N__43196\,
            I => \N__43193\
        );

    \I__9807\ : LocalMux
    port map (
            O => \N__43193\,
            I => \N__43190\
        );

    \I__9806\ : Span4Mux_h
    port map (
            O => \N__43190\,
            I => \N__43187\
        );

    \I__9805\ : Odrv4
    port map (
            O => \N__43187\,
            I => \current_shift_inst.un4_control_input_1_axb_12\
        );

    \I__9804\ : InMux
    port map (
            O => \N__43184\,
            I => \N__43178\
        );

    \I__9803\ : InMux
    port map (
            O => \N__43183\,
            I => \N__43178\
        );

    \I__9802\ : LocalMux
    port map (
            O => \N__43178\,
            I => \N__43174\
        );

    \I__9801\ : InMux
    port map (
            O => \N__43177\,
            I => \N__43171\
        );

    \I__9800\ : Odrv12
    port map (
            O => \N__43174\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__9799\ : LocalMux
    port map (
            O => \N__43171\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__9798\ : InMux
    port map (
            O => \N__43166\,
            I => \current_shift_inst.un4_control_input_1_cry_11\
        );

    \I__9797\ : InMux
    port map (
            O => \N__43163\,
            I => \N__43160\
        );

    \I__9796\ : LocalMux
    port map (
            O => \N__43160\,
            I => \N__43157\
        );

    \I__9795\ : Span12Mux_v
    port map (
            O => \N__43157\,
            I => \N__43154\
        );

    \I__9794\ : Odrv12
    port map (
            O => \N__43154\,
            I => \current_shift_inst.un4_control_input_1_axb_13\
        );

    \I__9793\ : InMux
    port map (
            O => \N__43151\,
            I => \N__43148\
        );

    \I__9792\ : LocalMux
    port map (
            O => \N__43148\,
            I => \N__43144\
        );

    \I__9791\ : InMux
    port map (
            O => \N__43147\,
            I => \N__43141\
        );

    \I__9790\ : Span4Mux_h
    port map (
            O => \N__43144\,
            I => \N__43137\
        );

    \I__9789\ : LocalMux
    port map (
            O => \N__43141\,
            I => \N__43134\
        );

    \I__9788\ : InMux
    port map (
            O => \N__43140\,
            I => \N__43131\
        );

    \I__9787\ : Odrv4
    port map (
            O => \N__43137\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__9786\ : Odrv12
    port map (
            O => \N__43134\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__9785\ : LocalMux
    port map (
            O => \N__43131\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__9784\ : InMux
    port map (
            O => \N__43124\,
            I => \current_shift_inst.un4_control_input_1_cry_12\
        );

    \I__9783\ : CascadeMux
    port map (
            O => \N__43121\,
            I => \N__43118\
        );

    \I__9782\ : InMux
    port map (
            O => \N__43118\,
            I => \N__43114\
        );

    \I__9781\ : CascadeMux
    port map (
            O => \N__43117\,
            I => \N__43111\
        );

    \I__9780\ : LocalMux
    port map (
            O => \N__43114\,
            I => \N__43108\
        );

    \I__9779\ : InMux
    port map (
            O => \N__43111\,
            I => \N__43105\
        );

    \I__9778\ : Span4Mux_v
    port map (
            O => \N__43108\,
            I => \N__43102\
        );

    \I__9777\ : LocalMux
    port map (
            O => \N__43105\,
            I => \N__43098\
        );

    \I__9776\ : Span4Mux_h
    port map (
            O => \N__43102\,
            I => \N__43095\
        );

    \I__9775\ : InMux
    port map (
            O => \N__43101\,
            I => \N__43092\
        );

    \I__9774\ : Odrv4
    port map (
            O => \N__43098\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__9773\ : Odrv4
    port map (
            O => \N__43095\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__9772\ : LocalMux
    port map (
            O => \N__43092\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__9771\ : InMux
    port map (
            O => \N__43085\,
            I => \current_shift_inst.un4_control_input_1_cry_13\
        );

    \I__9770\ : InMux
    port map (
            O => \N__43082\,
            I => \N__43079\
        );

    \I__9769\ : LocalMux
    port map (
            O => \N__43079\,
            I => \N__43076\
        );

    \I__9768\ : Span4Mux_h
    port map (
            O => \N__43076\,
            I => \N__43073\
        );

    \I__9767\ : Odrv4
    port map (
            O => \N__43073\,
            I => \current_shift_inst.un4_control_input_1_axb_15\
        );

    \I__9766\ : InMux
    port map (
            O => \N__43070\,
            I => \N__43066\
        );

    \I__9765\ : InMux
    port map (
            O => \N__43069\,
            I => \N__43063\
        );

    \I__9764\ : LocalMux
    port map (
            O => \N__43066\,
            I => \N__43059\
        );

    \I__9763\ : LocalMux
    port map (
            O => \N__43063\,
            I => \N__43056\
        );

    \I__9762\ : InMux
    port map (
            O => \N__43062\,
            I => \N__43053\
        );

    \I__9761\ : Odrv12
    port map (
            O => \N__43059\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__9760\ : Odrv4
    port map (
            O => \N__43056\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__9759\ : LocalMux
    port map (
            O => \N__43053\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__9758\ : InMux
    port map (
            O => \N__43046\,
            I => \current_shift_inst.un4_control_input_1_cry_14\
        );

    \I__9757\ : InMux
    port map (
            O => \N__43043\,
            I => \N__43040\
        );

    \I__9756\ : LocalMux
    port map (
            O => \N__43040\,
            I => \N__43037\
        );

    \I__9755\ : Span4Mux_h
    port map (
            O => \N__43037\,
            I => \N__43034\
        );

    \I__9754\ : Odrv4
    port map (
            O => \N__43034\,
            I => \current_shift_inst.un4_control_input_1_axb_16\
        );

    \I__9753\ : InMux
    port map (
            O => \N__43031\,
            I => \N__43028\
        );

    \I__9752\ : LocalMux
    port map (
            O => \N__43028\,
            I => \N__43024\
        );

    \I__9751\ : InMux
    port map (
            O => \N__43027\,
            I => \N__43021\
        );

    \I__9750\ : Span4Mux_h
    port map (
            O => \N__43024\,
            I => \N__43018\
        );

    \I__9749\ : LocalMux
    port map (
            O => \N__43021\,
            I => \N__43014\
        );

    \I__9748\ : Span4Mux_h
    port map (
            O => \N__43018\,
            I => \N__43011\
        );

    \I__9747\ : InMux
    port map (
            O => \N__43017\,
            I => \N__43008\
        );

    \I__9746\ : Odrv4
    port map (
            O => \N__43014\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__9745\ : Odrv4
    port map (
            O => \N__43011\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__9744\ : LocalMux
    port map (
            O => \N__43008\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__9743\ : InMux
    port map (
            O => \N__43001\,
            I => \current_shift_inst.un4_control_input_1_cry_15\
        );

    \I__9742\ : InMux
    port map (
            O => \N__42998\,
            I => \N__42995\
        );

    \I__9741\ : LocalMux
    port map (
            O => \N__42995\,
            I => \N__42990\
        );

    \I__9740\ : CascadeMux
    port map (
            O => \N__42994\,
            I => \N__42987\
        );

    \I__9739\ : InMux
    port map (
            O => \N__42993\,
            I => \N__42984\
        );

    \I__9738\ : Span4Mux_h
    port map (
            O => \N__42990\,
            I => \N__42981\
        );

    \I__9737\ : InMux
    port map (
            O => \N__42987\,
            I => \N__42978\
        );

    \I__9736\ : LocalMux
    port map (
            O => \N__42984\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__9735\ : Odrv4
    port map (
            O => \N__42981\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__9734\ : LocalMux
    port map (
            O => \N__42978\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__9733\ : InMux
    port map (
            O => \N__42971\,
            I => \bfn_18_16_0_\
        );

    \I__9732\ : InMux
    port map (
            O => \N__42968\,
            I => \N__42965\
        );

    \I__9731\ : LocalMux
    port map (
            O => \N__42965\,
            I => \N__42962\
        );

    \I__9730\ : Span4Mux_h
    port map (
            O => \N__42962\,
            I => \N__42959\
        );

    \I__9729\ : Odrv4
    port map (
            O => \N__42959\,
            I => \current_shift_inst.un4_control_input_1_axb_18\
        );

    \I__9728\ : InMux
    port map (
            O => \N__42956\,
            I => \N__42952\
        );

    \I__9727\ : InMux
    port map (
            O => \N__42955\,
            I => \N__42949\
        );

    \I__9726\ : LocalMux
    port map (
            O => \N__42952\,
            I => \N__42943\
        );

    \I__9725\ : LocalMux
    port map (
            O => \N__42949\,
            I => \N__42943\
        );

    \I__9724\ : InMux
    port map (
            O => \N__42948\,
            I => \N__42940\
        );

    \I__9723\ : Odrv12
    port map (
            O => \N__42943\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__9722\ : LocalMux
    port map (
            O => \N__42940\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__9721\ : InMux
    port map (
            O => \N__42935\,
            I => \current_shift_inst.un4_control_input_1_cry_17\
        );

    \I__9720\ : CascadeMux
    port map (
            O => \N__42932\,
            I => \N__42928\
        );

    \I__9719\ : InMux
    port map (
            O => \N__42931\,
            I => \N__42924\
        );

    \I__9718\ : InMux
    port map (
            O => \N__42928\,
            I => \N__42921\
        );

    \I__9717\ : InMux
    port map (
            O => \N__42927\,
            I => \N__42918\
        );

    \I__9716\ : LocalMux
    port map (
            O => \N__42924\,
            I => \N__42915\
        );

    \I__9715\ : LocalMux
    port map (
            O => \N__42921\,
            I => \N__42910\
        );

    \I__9714\ : LocalMux
    port map (
            O => \N__42918\,
            I => \N__42910\
        );

    \I__9713\ : Odrv12
    port map (
            O => \N__42915\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__9712\ : Odrv4
    port map (
            O => \N__42910\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__9711\ : InMux
    port map (
            O => \N__42905\,
            I => \current_shift_inst.un4_control_input_1_cry_18\
        );

    \I__9710\ : InMux
    port map (
            O => \N__42902\,
            I => \N__42899\
        );

    \I__9709\ : LocalMux
    port map (
            O => \N__42899\,
            I => \N__42896\
        );

    \I__9708\ : Span4Mux_h
    port map (
            O => \N__42896\,
            I => \N__42893\
        );

    \I__9707\ : Odrv4
    port map (
            O => \N__42893\,
            I => \current_shift_inst.un4_control_input_1_axb_4\
        );

    \I__9706\ : CascadeMux
    port map (
            O => \N__42890\,
            I => \N__42886\
        );

    \I__9705\ : CascadeMux
    port map (
            O => \N__42889\,
            I => \N__42883\
        );

    \I__9704\ : InMux
    port map (
            O => \N__42886\,
            I => \N__42880\
        );

    \I__9703\ : InMux
    port map (
            O => \N__42883\,
            I => \N__42877\
        );

    \I__9702\ : LocalMux
    port map (
            O => \N__42880\,
            I => \N__42871\
        );

    \I__9701\ : LocalMux
    port map (
            O => \N__42877\,
            I => \N__42871\
        );

    \I__9700\ : InMux
    port map (
            O => \N__42876\,
            I => \N__42868\
        );

    \I__9699\ : Odrv12
    port map (
            O => \N__42871\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__9698\ : LocalMux
    port map (
            O => \N__42868\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__9697\ : InMux
    port map (
            O => \N__42863\,
            I => \current_shift_inst.un4_control_input_1_cry_3\
        );

    \I__9696\ : InMux
    port map (
            O => \N__42860\,
            I => \N__42857\
        );

    \I__9695\ : LocalMux
    port map (
            O => \N__42857\,
            I => \N__42854\
        );

    \I__9694\ : Span4Mux_h
    port map (
            O => \N__42854\,
            I => \N__42851\
        );

    \I__9693\ : Span4Mux_v
    port map (
            O => \N__42851\,
            I => \N__42848\
        );

    \I__9692\ : Odrv4
    port map (
            O => \N__42848\,
            I => \current_shift_inst.un4_control_input_1_axb_5\
        );

    \I__9691\ : InMux
    port map (
            O => \N__42845\,
            I => \N__42839\
        );

    \I__9690\ : InMux
    port map (
            O => \N__42844\,
            I => \N__42839\
        );

    \I__9689\ : LocalMux
    port map (
            O => \N__42839\,
            I => \N__42835\
        );

    \I__9688\ : InMux
    port map (
            O => \N__42838\,
            I => \N__42832\
        );

    \I__9687\ : Odrv4
    port map (
            O => \N__42835\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__9686\ : LocalMux
    port map (
            O => \N__42832\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__9685\ : InMux
    port map (
            O => \N__42827\,
            I => \current_shift_inst.un4_control_input_1_cry_4\
        );

    \I__9684\ : InMux
    port map (
            O => \N__42824\,
            I => \N__42821\
        );

    \I__9683\ : LocalMux
    port map (
            O => \N__42821\,
            I => \current_shift_inst.un4_control_input_1_axb_6\
        );

    \I__9682\ : InMux
    port map (
            O => \N__42818\,
            I => \current_shift_inst.un4_control_input_1_cry_5\
        );

    \I__9681\ : InMux
    port map (
            O => \N__42815\,
            I => \N__42812\
        );

    \I__9680\ : LocalMux
    port map (
            O => \N__42812\,
            I => \N__42809\
        );

    \I__9679\ : Span12Mux_v
    port map (
            O => \N__42809\,
            I => \N__42806\
        );

    \I__9678\ : Odrv12
    port map (
            O => \N__42806\,
            I => \current_shift_inst.un4_control_input_1_axb_7\
        );

    \I__9677\ : InMux
    port map (
            O => \N__42803\,
            I => \N__42800\
        );

    \I__9676\ : LocalMux
    port map (
            O => \N__42800\,
            I => \N__42796\
        );

    \I__9675\ : InMux
    port map (
            O => \N__42799\,
            I => \N__42793\
        );

    \I__9674\ : Span4Mux_h
    port map (
            O => \N__42796\,
            I => \N__42789\
        );

    \I__9673\ : LocalMux
    port map (
            O => \N__42793\,
            I => \N__42786\
        );

    \I__9672\ : InMux
    port map (
            O => \N__42792\,
            I => \N__42783\
        );

    \I__9671\ : Odrv4
    port map (
            O => \N__42789\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__9670\ : Odrv12
    port map (
            O => \N__42786\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__9669\ : LocalMux
    port map (
            O => \N__42783\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__9668\ : InMux
    port map (
            O => \N__42776\,
            I => \current_shift_inst.un4_control_input_1_cry_6\
        );

    \I__9667\ : InMux
    port map (
            O => \N__42773\,
            I => \N__42770\
        );

    \I__9666\ : LocalMux
    port map (
            O => \N__42770\,
            I => \N__42767\
        );

    \I__9665\ : Span4Mux_v
    port map (
            O => \N__42767\,
            I => \N__42764\
        );

    \I__9664\ : Odrv4
    port map (
            O => \N__42764\,
            I => \current_shift_inst.un4_control_input_1_axb_8\
        );

    \I__9663\ : InMux
    port map (
            O => \N__42761\,
            I => \N__42757\
        );

    \I__9662\ : CascadeMux
    port map (
            O => \N__42760\,
            I => \N__42754\
        );

    \I__9661\ : LocalMux
    port map (
            O => \N__42757\,
            I => \N__42751\
        );

    \I__9660\ : InMux
    port map (
            O => \N__42754\,
            I => \N__42748\
        );

    \I__9659\ : Span4Mux_v
    port map (
            O => \N__42751\,
            I => \N__42742\
        );

    \I__9658\ : LocalMux
    port map (
            O => \N__42748\,
            I => \N__42742\
        );

    \I__9657\ : InMux
    port map (
            O => \N__42747\,
            I => \N__42739\
        );

    \I__9656\ : Odrv4
    port map (
            O => \N__42742\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__9655\ : LocalMux
    port map (
            O => \N__42739\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__9654\ : InMux
    port map (
            O => \N__42734\,
            I => \current_shift_inst.un4_control_input_1_cry_7\
        );

    \I__9653\ : InMux
    port map (
            O => \N__42731\,
            I => \N__42728\
        );

    \I__9652\ : LocalMux
    port map (
            O => \N__42728\,
            I => \N__42725\
        );

    \I__9651\ : Span4Mux_h
    port map (
            O => \N__42725\,
            I => \N__42722\
        );

    \I__9650\ : Odrv4
    port map (
            O => \N__42722\,
            I => \current_shift_inst.un4_control_input_1_axb_9\
        );

    \I__9649\ : CascadeMux
    port map (
            O => \N__42719\,
            I => \N__42716\
        );

    \I__9648\ : InMux
    port map (
            O => \N__42716\,
            I => \N__42712\
        );

    \I__9647\ : InMux
    port map (
            O => \N__42715\,
            I => \N__42709\
        );

    \I__9646\ : LocalMux
    port map (
            O => \N__42712\,
            I => \N__42706\
        );

    \I__9645\ : LocalMux
    port map (
            O => \N__42709\,
            I => \N__42703\
        );

    \I__9644\ : Span4Mux_h
    port map (
            O => \N__42706\,
            I => \N__42697\
        );

    \I__9643\ : Span4Mux_h
    port map (
            O => \N__42703\,
            I => \N__42697\
        );

    \I__9642\ : InMux
    port map (
            O => \N__42702\,
            I => \N__42694\
        );

    \I__9641\ : Odrv4
    port map (
            O => \N__42697\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__9640\ : LocalMux
    port map (
            O => \N__42694\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__9639\ : InMux
    port map (
            O => \N__42689\,
            I => \bfn_18_15_0_\
        );

    \I__9638\ : InMux
    port map (
            O => \N__42686\,
            I => \N__42683\
        );

    \I__9637\ : LocalMux
    port map (
            O => \N__42683\,
            I => \N__42680\
        );

    \I__9636\ : Span4Mux_h
    port map (
            O => \N__42680\,
            I => \N__42677\
        );

    \I__9635\ : Span4Mux_h
    port map (
            O => \N__42677\,
            I => \N__42674\
        );

    \I__9634\ : Odrv4
    port map (
            O => \N__42674\,
            I => \current_shift_inst.un4_control_input_1_axb_10\
        );

    \I__9633\ : CascadeMux
    port map (
            O => \N__42671\,
            I => \N__42667\
        );

    \I__9632\ : InMux
    port map (
            O => \N__42670\,
            I => \N__42664\
        );

    \I__9631\ : InMux
    port map (
            O => \N__42667\,
            I => \N__42661\
        );

    \I__9630\ : LocalMux
    port map (
            O => \N__42664\,
            I => \N__42655\
        );

    \I__9629\ : LocalMux
    port map (
            O => \N__42661\,
            I => \N__42655\
        );

    \I__9628\ : InMux
    port map (
            O => \N__42660\,
            I => \N__42652\
        );

    \I__9627\ : Odrv12
    port map (
            O => \N__42655\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__9626\ : LocalMux
    port map (
            O => \N__42652\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__9625\ : InMux
    port map (
            O => \N__42647\,
            I => \current_shift_inst.un4_control_input_1_cry_9\
        );

    \I__9624\ : InMux
    port map (
            O => \N__42644\,
            I => \N__42641\
        );

    \I__9623\ : LocalMux
    port map (
            O => \N__42641\,
            I => \N__42638\
        );

    \I__9622\ : Span4Mux_v
    port map (
            O => \N__42638\,
            I => \N__42635\
        );

    \I__9621\ : Odrv4
    port map (
            O => \N__42635\,
            I => \current_shift_inst.un4_control_input_1_axb_11\
        );

    \I__9620\ : InMux
    port map (
            O => \N__42632\,
            I => \N__42628\
        );

    \I__9619\ : InMux
    port map (
            O => \N__42631\,
            I => \N__42625\
        );

    \I__9618\ : LocalMux
    port map (
            O => \N__42628\,
            I => \N__42622\
        );

    \I__9617\ : LocalMux
    port map (
            O => \N__42625\,
            I => \N__42618\
        );

    \I__9616\ : Span4Mux_h
    port map (
            O => \N__42622\,
            I => \N__42615\
        );

    \I__9615\ : InMux
    port map (
            O => \N__42621\,
            I => \N__42612\
        );

    \I__9614\ : Odrv12
    port map (
            O => \N__42618\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__9613\ : Odrv4
    port map (
            O => \N__42615\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__9612\ : LocalMux
    port map (
            O => \N__42612\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__9611\ : InMux
    port map (
            O => \N__42605\,
            I => \current_shift_inst.un4_control_input_1_cry_10\
        );

    \I__9610\ : CascadeMux
    port map (
            O => \N__42602\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18_cascade_\
        );

    \I__9609\ : InMux
    port map (
            O => \N__42599\,
            I => \N__42593\
        );

    \I__9608\ : InMux
    port map (
            O => \N__42598\,
            I => \N__42588\
        );

    \I__9607\ : InMux
    port map (
            O => \N__42597\,
            I => \N__42588\
        );

    \I__9606\ : InMux
    port map (
            O => \N__42596\,
            I => \N__42585\
        );

    \I__9605\ : LocalMux
    port map (
            O => \N__42593\,
            I => \N__42582\
        );

    \I__9604\ : LocalMux
    port map (
            O => \N__42588\,
            I => \N__42579\
        );

    \I__9603\ : LocalMux
    port map (
            O => \N__42585\,
            I => \N__42576\
        );

    \I__9602\ : Span4Mux_v
    port map (
            O => \N__42582\,
            I => \N__42573\
        );

    \I__9601\ : Span4Mux_h
    port map (
            O => \N__42579\,
            I => \N__42570\
        );

    \I__9600\ : Span12Mux_s10_h
    port map (
            O => \N__42576\,
            I => \N__42567\
        );

    \I__9599\ : Odrv4
    port map (
            O => \N__42573\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__9598\ : Odrv4
    port map (
            O => \N__42570\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__9597\ : Odrv12
    port map (
            O => \N__42567\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__9596\ : InMux
    port map (
            O => \N__42560\,
            I => \N__42554\
        );

    \I__9595\ : InMux
    port map (
            O => \N__42559\,
            I => \N__42554\
        );

    \I__9594\ : LocalMux
    port map (
            O => \N__42554\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\
        );

    \I__9593\ : InMux
    port map (
            O => \N__42551\,
            I => \N__42548\
        );

    \I__9592\ : LocalMux
    port map (
            O => \N__42548\,
            I => \N__42542\
        );

    \I__9591\ : InMux
    port map (
            O => \N__42547\,
            I => \N__42537\
        );

    \I__9590\ : InMux
    port map (
            O => \N__42546\,
            I => \N__42537\
        );

    \I__9589\ : InMux
    port map (
            O => \N__42545\,
            I => \N__42534\
        );

    \I__9588\ : Span4Mux_v
    port map (
            O => \N__42542\,
            I => \N__42529\
        );

    \I__9587\ : LocalMux
    port map (
            O => \N__42537\,
            I => \N__42529\
        );

    \I__9586\ : LocalMux
    port map (
            O => \N__42534\,
            I => \N__42526\
        );

    \I__9585\ : Span4Mux_h
    port map (
            O => \N__42529\,
            I => \N__42523\
        );

    \I__9584\ : Odrv12
    port map (
            O => \N__42526\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\
        );

    \I__9583\ : Odrv4
    port map (
            O => \N__42523\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\
        );

    \I__9582\ : InMux
    port map (
            O => \N__42518\,
            I => \N__42514\
        );

    \I__9581\ : InMux
    port map (
            O => \N__42517\,
            I => \N__42511\
        );

    \I__9580\ : LocalMux
    port map (
            O => \N__42514\,
            I => \N__42507\
        );

    \I__9579\ : LocalMux
    port map (
            O => \N__42511\,
            I => \N__42504\
        );

    \I__9578\ : InMux
    port map (
            O => \N__42510\,
            I => \N__42501\
        );

    \I__9577\ : Span4Mux_h
    port map (
            O => \N__42507\,
            I => \N__42498\
        );

    \I__9576\ : Span4Mux_v
    port map (
            O => \N__42504\,
            I => \N__42495\
        );

    \I__9575\ : LocalMux
    port map (
            O => \N__42501\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15\
        );

    \I__9574\ : Odrv4
    port map (
            O => \N__42498\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15\
        );

    \I__9573\ : Odrv4
    port map (
            O => \N__42495\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15\
        );

    \I__9572\ : InMux
    port map (
            O => \N__42488\,
            I => \N__42485\
        );

    \I__9571\ : LocalMux
    port map (
            O => \N__42485\,
            I => \N__42482\
        );

    \I__9570\ : Odrv4
    port map (
            O => \N__42482\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\
        );

    \I__9569\ : InMux
    port map (
            O => \N__42479\,
            I => \N__42476\
        );

    \I__9568\ : LocalMux
    port map (
            O => \N__42476\,
            I => \N__42473\
        );

    \I__9567\ : Span4Mux_v
    port map (
            O => \N__42473\,
            I => \N__42470\
        );

    \I__9566\ : Odrv4
    port map (
            O => \N__42470\,
            I => \current_shift_inst.un38_control_input_axb_31_s0\
        );

    \I__9565\ : InMux
    port map (
            O => \N__42467\,
            I => \N__42463\
        );

    \I__9564\ : InMux
    port map (
            O => \N__42466\,
            I => \N__42459\
        );

    \I__9563\ : LocalMux
    port map (
            O => \N__42463\,
            I => \N__42456\
        );

    \I__9562\ : InMux
    port map (
            O => \N__42462\,
            I => \N__42453\
        );

    \I__9561\ : LocalMux
    port map (
            O => \N__42459\,
            I => \N__42450\
        );

    \I__9560\ : Span4Mux_v
    port map (
            O => \N__42456\,
            I => \N__42445\
        );

    \I__9559\ : LocalMux
    port map (
            O => \N__42453\,
            I => \N__42445\
        );

    \I__9558\ : Span4Mux_h
    port map (
            O => \N__42450\,
            I => \N__42441\
        );

    \I__9557\ : Span4Mux_h
    port map (
            O => \N__42445\,
            I => \N__42438\
        );

    \I__9556\ : InMux
    port map (
            O => \N__42444\,
            I => \N__42435\
        );

    \I__9555\ : Odrv4
    port map (
            O => \N__42441\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__9554\ : Odrv4
    port map (
            O => \N__42438\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__9553\ : LocalMux
    port map (
            O => \N__42435\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__9552\ : InMux
    port map (
            O => \N__42428\,
            I => \N__42425\
        );

    \I__9551\ : LocalMux
    port map (
            O => \N__42425\,
            I => \N__42422\
        );

    \I__9550\ : Span4Mux_h
    port map (
            O => \N__42422\,
            I => \N__42419\
        );

    \I__9549\ : Odrv4
    port map (
            O => \N__42419\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\
        );

    \I__9548\ : InMux
    port map (
            O => \N__42416\,
            I => \N__42411\
        );

    \I__9547\ : InMux
    port map (
            O => \N__42415\,
            I => \N__42408\
        );

    \I__9546\ : InMux
    port map (
            O => \N__42414\,
            I => \N__42405\
        );

    \I__9545\ : LocalMux
    port map (
            O => \N__42411\,
            I => \N__42400\
        );

    \I__9544\ : LocalMux
    port map (
            O => \N__42408\,
            I => \N__42400\
        );

    \I__9543\ : LocalMux
    port map (
            O => \N__42405\,
            I => \N__42397\
        );

    \I__9542\ : Span4Mux_v
    port map (
            O => \N__42400\,
            I => \N__42394\
        );

    \I__9541\ : Span12Mux_s10_h
    port map (
            O => \N__42397\,
            I => \N__42391\
        );

    \I__9540\ : Span4Mux_v
    port map (
            O => \N__42394\,
            I => \N__42388\
        );

    \I__9539\ : Odrv12
    port map (
            O => \N__42391\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__9538\ : Odrv4
    port map (
            O => \N__42388\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__9537\ : InMux
    port map (
            O => \N__42383\,
            I => \N__42377\
        );

    \I__9536\ : InMux
    port map (
            O => \N__42382\,
            I => \N__42374\
        );

    \I__9535\ : InMux
    port map (
            O => \N__42381\,
            I => \N__42371\
        );

    \I__9534\ : InMux
    port map (
            O => \N__42380\,
            I => \N__42355\
        );

    \I__9533\ : LocalMux
    port map (
            O => \N__42377\,
            I => \N__42352\
        );

    \I__9532\ : LocalMux
    port map (
            O => \N__42374\,
            I => \N__42349\
        );

    \I__9531\ : LocalMux
    port map (
            O => \N__42371\,
            I => \N__42346\
        );

    \I__9530\ : InMux
    port map (
            O => \N__42370\,
            I => \N__42331\
        );

    \I__9529\ : InMux
    port map (
            O => \N__42369\,
            I => \N__42331\
        );

    \I__9528\ : InMux
    port map (
            O => \N__42368\,
            I => \N__42331\
        );

    \I__9527\ : InMux
    port map (
            O => \N__42367\,
            I => \N__42331\
        );

    \I__9526\ : InMux
    port map (
            O => \N__42366\,
            I => \N__42331\
        );

    \I__9525\ : InMux
    port map (
            O => \N__42365\,
            I => \N__42331\
        );

    \I__9524\ : InMux
    port map (
            O => \N__42364\,
            I => \N__42331\
        );

    \I__9523\ : InMux
    port map (
            O => \N__42363\,
            I => \N__42318\
        );

    \I__9522\ : InMux
    port map (
            O => \N__42362\,
            I => \N__42318\
        );

    \I__9521\ : InMux
    port map (
            O => \N__42361\,
            I => \N__42318\
        );

    \I__9520\ : InMux
    port map (
            O => \N__42360\,
            I => \N__42318\
        );

    \I__9519\ : InMux
    port map (
            O => \N__42359\,
            I => \N__42318\
        );

    \I__9518\ : InMux
    port map (
            O => \N__42358\,
            I => \N__42318\
        );

    \I__9517\ : LocalMux
    port map (
            O => \N__42355\,
            I => \N__42305\
        );

    \I__9516\ : Span4Mux_h
    port map (
            O => \N__42352\,
            I => \N__42305\
        );

    \I__9515\ : Span4Mux_v
    port map (
            O => \N__42349\,
            I => \N__42296\
        );

    \I__9514\ : Span4Mux_h
    port map (
            O => \N__42346\,
            I => \N__42296\
        );

    \I__9513\ : LocalMux
    port map (
            O => \N__42331\,
            I => \N__42296\
        );

    \I__9512\ : LocalMux
    port map (
            O => \N__42318\,
            I => \N__42296\
        );

    \I__9511\ : InMux
    port map (
            O => \N__42317\,
            I => \N__42287\
        );

    \I__9510\ : InMux
    port map (
            O => \N__42316\,
            I => \N__42287\
        );

    \I__9509\ : InMux
    port map (
            O => \N__42315\,
            I => \N__42287\
        );

    \I__9508\ : InMux
    port map (
            O => \N__42314\,
            I => \N__42287\
        );

    \I__9507\ : InMux
    port map (
            O => \N__42313\,
            I => \N__42278\
        );

    \I__9506\ : InMux
    port map (
            O => \N__42312\,
            I => \N__42278\
        );

    \I__9505\ : InMux
    port map (
            O => \N__42311\,
            I => \N__42278\
        );

    \I__9504\ : InMux
    port map (
            O => \N__42310\,
            I => \N__42278\
        );

    \I__9503\ : Span4Mux_h
    port map (
            O => \N__42305\,
            I => \N__42275\
        );

    \I__9502\ : Odrv4
    port map (
            O => \N__42296\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__9501\ : LocalMux
    port map (
            O => \N__42287\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__9500\ : LocalMux
    port map (
            O => \N__42278\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__9499\ : Odrv4
    port map (
            O => \N__42275\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__9498\ : CascadeMux
    port map (
            O => \N__42266\,
            I => \N__42262\
        );

    \I__9497\ : InMux
    port map (
            O => \N__42265\,
            I => \N__42258\
        );

    \I__9496\ : InMux
    port map (
            O => \N__42262\,
            I => \N__42255\
        );

    \I__9495\ : InMux
    port map (
            O => \N__42261\,
            I => \N__42252\
        );

    \I__9494\ : LocalMux
    port map (
            O => \N__42258\,
            I => \N__42247\
        );

    \I__9493\ : LocalMux
    port map (
            O => \N__42255\,
            I => \N__42247\
        );

    \I__9492\ : LocalMux
    port map (
            O => \N__42252\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__9491\ : Odrv12
    port map (
            O => \N__42247\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__9490\ : InMux
    port map (
            O => \N__42242\,
            I => \N__42239\
        );

    \I__9489\ : LocalMux
    port map (
            O => \N__42239\,
            I => \N__42236\
        );

    \I__9488\ : Span4Mux_h
    port map (
            O => \N__42236\,
            I => \N__42233\
        );

    \I__9487\ : Span4Mux_v
    port map (
            O => \N__42233\,
            I => \N__42230\
        );

    \I__9486\ : Odrv4
    port map (
            O => \N__42230\,
            I => \current_shift_inst.un4_control_input_1_axb_2\
        );

    \I__9485\ : InMux
    port map (
            O => \N__42227\,
            I => \N__42221\
        );

    \I__9484\ : InMux
    port map (
            O => \N__42226\,
            I => \N__42221\
        );

    \I__9483\ : LocalMux
    port map (
            O => \N__42221\,
            I => \N__42218\
        );

    \I__9482\ : Span4Mux_h
    port map (
            O => \N__42218\,
            I => \N__42214\
        );

    \I__9481\ : InMux
    port map (
            O => \N__42217\,
            I => \N__42211\
        );

    \I__9480\ : Odrv4
    port map (
            O => \N__42214\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__9479\ : LocalMux
    port map (
            O => \N__42211\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__9478\ : InMux
    port map (
            O => \N__42206\,
            I => \current_shift_inst.un4_control_input_1_cry_1\
        );

    \I__9477\ : InMux
    port map (
            O => \N__42203\,
            I => \N__42200\
        );

    \I__9476\ : LocalMux
    port map (
            O => \N__42200\,
            I => \N__42197\
        );

    \I__9475\ : Span4Mux_h
    port map (
            O => \N__42197\,
            I => \N__42194\
        );

    \I__9474\ : Odrv4
    port map (
            O => \N__42194\,
            I => \current_shift_inst.un4_control_input_1_axb_3\
        );

    \I__9473\ : InMux
    port map (
            O => \N__42191\,
            I => \N__42187\
        );

    \I__9472\ : InMux
    port map (
            O => \N__42190\,
            I => \N__42184\
        );

    \I__9471\ : LocalMux
    port map (
            O => \N__42187\,
            I => \N__42181\
        );

    \I__9470\ : LocalMux
    port map (
            O => \N__42184\,
            I => \N__42178\
        );

    \I__9469\ : Span4Mux_v
    port map (
            O => \N__42181\,
            I => \N__42172\
        );

    \I__9468\ : Span4Mux_h
    port map (
            O => \N__42178\,
            I => \N__42172\
        );

    \I__9467\ : InMux
    port map (
            O => \N__42177\,
            I => \N__42169\
        );

    \I__9466\ : Odrv4
    port map (
            O => \N__42172\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__9465\ : LocalMux
    port map (
            O => \N__42169\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__9464\ : InMux
    port map (
            O => \N__42164\,
            I => \current_shift_inst.un4_control_input_1_cry_2\
        );

    \I__9463\ : CascadeMux
    port map (
            O => \N__42161\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0_cascade_\
        );

    \I__9462\ : CascadeMux
    port map (
            O => \N__42158\,
            I => \N__42155\
        );

    \I__9461\ : InMux
    port map (
            O => \N__42155\,
            I => \N__42152\
        );

    \I__9460\ : LocalMux
    port map (
            O => \N__42152\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4Z0Z_28\
        );

    \I__9459\ : CascadeMux
    port map (
            O => \N__42149\,
            I => \N__42146\
        );

    \I__9458\ : InMux
    port map (
            O => \N__42146\,
            I => \N__42142\
        );

    \I__9457\ : InMux
    port map (
            O => \N__42145\,
            I => \N__42139\
        );

    \I__9456\ : LocalMux
    port map (
            O => \N__42142\,
            I => \N__42136\
        );

    \I__9455\ : LocalMux
    port map (
            O => \N__42139\,
            I => \N__42133\
        );

    \I__9454\ : Span4Mux_h
    port map (
            O => \N__42136\,
            I => \N__42130\
        );

    \I__9453\ : Span12Mux_v
    port map (
            O => \N__42133\,
            I => \N__42127\
        );

    \I__9452\ : Odrv4
    port map (
            O => \N__42130\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__9451\ : Odrv12
    port map (
            O => \N__42127\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__9450\ : InMux
    port map (
            O => \N__42122\,
            I => \N__42118\
        );

    \I__9449\ : InMux
    port map (
            O => \N__42121\,
            I => \N__42115\
        );

    \I__9448\ : LocalMux
    port map (
            O => \N__42118\,
            I => \phase_controller_inst1.stoper_tr.runningZ0\
        );

    \I__9447\ : LocalMux
    port map (
            O => \N__42115\,
            I => \phase_controller_inst1.stoper_tr.runningZ0\
        );

    \I__9446\ : InMux
    port map (
            O => \N__42110\,
            I => \N__42106\
        );

    \I__9445\ : InMux
    port map (
            O => \N__42109\,
            I => \N__42103\
        );

    \I__9444\ : LocalMux
    port map (
            O => \N__42106\,
            I => \N__42100\
        );

    \I__9443\ : LocalMux
    port map (
            O => \N__42103\,
            I => \N__42097\
        );

    \I__9442\ : Span4Mux_h
    port map (
            O => \N__42100\,
            I => \N__42094\
        );

    \I__9441\ : Span4Mux_v
    port map (
            O => \N__42097\,
            I => \N__42091\
        );

    \I__9440\ : Odrv4
    port map (
            O => \N__42094\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt30\
        );

    \I__9439\ : Odrv4
    port map (
            O => \N__42091\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt30\
        );

    \I__9438\ : CascadeMux
    port map (
            O => \N__42086\,
            I => \N__42083\
        );

    \I__9437\ : InMux
    port map (
            O => \N__42083\,
            I => \N__42080\
        );

    \I__9436\ : LocalMux
    port map (
            O => \N__42080\,
            I => \N__42077\
        );

    \I__9435\ : Odrv4
    port map (
            O => \N__42077\,
            I => \phase_controller_inst1.stoper_tr.un4_running_df30\
        );

    \I__9434\ : InMux
    port map (
            O => \N__42074\,
            I => \N__42071\
        );

    \I__9433\ : LocalMux
    port map (
            O => \N__42071\,
            I => \N__42068\
        );

    \I__9432\ : Span4Mux_h
    port map (
            O => \N__42068\,
            I => \N__42065\
        );

    \I__9431\ : Odrv4
    port map (
            O => \N__42065\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO\
        );

    \I__9430\ : InMux
    port map (
            O => \N__42062\,
            I => \N__42059\
        );

    \I__9429\ : LocalMux
    port map (
            O => \N__42059\,
            I => \N__42055\
        );

    \I__9428\ : InMux
    port map (
            O => \N__42058\,
            I => \N__42052\
        );

    \I__9427\ : Odrv12
    port map (
            O => \N__42055\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\
        );

    \I__9426\ : LocalMux
    port map (
            O => \N__42052\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\
        );

    \I__9425\ : CascadeMux
    port map (
            O => \N__42047\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\
        );

    \I__9424\ : InMux
    port map (
            O => \N__42044\,
            I => \N__42041\
        );

    \I__9423\ : LocalMux
    port map (
            O => \N__42041\,
            I => \N__42037\
        );

    \I__9422\ : InMux
    port map (
            O => \N__42040\,
            I => \N__42034\
        );

    \I__9421\ : Span4Mux_v
    port map (
            O => \N__42037\,
            I => \N__42031\
        );

    \I__9420\ : LocalMux
    port map (
            O => \N__42034\,
            I => \N__42028\
        );

    \I__9419\ : Span4Mux_v
    port map (
            O => \N__42031\,
            I => \N__42025\
        );

    \I__9418\ : Span4Mux_v
    port map (
            O => \N__42028\,
            I => \N__42022\
        );

    \I__9417\ : Span4Mux_h
    port map (
            O => \N__42025\,
            I => \N__42017\
        );

    \I__9416\ : Span4Mux_h
    port map (
            O => \N__42022\,
            I => \N__42014\
        );

    \I__9415\ : InMux
    port map (
            O => \N__42021\,
            I => \N__42009\
        );

    \I__9414\ : InMux
    port map (
            O => \N__42020\,
            I => \N__42009\
        );

    \I__9413\ : Odrv4
    port map (
            O => \N__42017\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__9412\ : Odrv4
    port map (
            O => \N__42014\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__9411\ : LocalMux
    port map (
            O => \N__42009\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__9410\ : InMux
    port map (
            O => \N__42002\,
            I => \N__41999\
        );

    \I__9409\ : LocalMux
    port map (
            O => \N__41999\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\
        );

    \I__9408\ : InMux
    port map (
            O => \N__41996\,
            I => \N__41993\
        );

    \I__9407\ : LocalMux
    port map (
            O => \N__41993\,
            I => \N__41990\
        );

    \I__9406\ : Span4Mux_h
    port map (
            O => \N__41990\,
            I => \N__41987\
        );

    \I__9405\ : Odrv4
    port map (
            O => \N__41987\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt18\
        );

    \I__9404\ : InMux
    port map (
            O => \N__41984\,
            I => \N__41979\
        );

    \I__9403\ : InMux
    port map (
            O => \N__41983\,
            I => \N__41974\
        );

    \I__9402\ : InMux
    port map (
            O => \N__41982\,
            I => \N__41974\
        );

    \I__9401\ : LocalMux
    port map (
            O => \N__41979\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__9400\ : LocalMux
    port map (
            O => \N__41974\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__9399\ : CascadeMux
    port map (
            O => \N__41969\,
            I => \N__41965\
        );

    \I__9398\ : InMux
    port map (
            O => \N__41968\,
            I => \N__41961\
        );

    \I__9397\ : InMux
    port map (
            O => \N__41965\,
            I => \N__41956\
        );

    \I__9396\ : InMux
    port map (
            O => \N__41964\,
            I => \N__41956\
        );

    \I__9395\ : LocalMux
    port map (
            O => \N__41961\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__9394\ : LocalMux
    port map (
            O => \N__41956\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__9393\ : CascadeMux
    port map (
            O => \N__41951\,
            I => \N__41948\
        );

    \I__9392\ : InMux
    port map (
            O => \N__41948\,
            I => \N__41945\
        );

    \I__9391\ : LocalMux
    port map (
            O => \N__41945\,
            I => \N__41942\
        );

    \I__9390\ : Span4Mux_h
    port map (
            O => \N__41942\,
            I => \N__41939\
        );

    \I__9389\ : Odrv4
    port map (
            O => \N__41939\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\
        );

    \I__9388\ : InMux
    port map (
            O => \N__41936\,
            I => \N__41932\
        );

    \I__9387\ : CascadeMux
    port map (
            O => \N__41935\,
            I => \N__41929\
        );

    \I__9386\ : LocalMux
    port map (
            O => \N__41932\,
            I => \N__41926\
        );

    \I__9385\ : InMux
    port map (
            O => \N__41929\,
            I => \N__41922\
        );

    \I__9384\ : Span4Mux_v
    port map (
            O => \N__41926\,
            I => \N__41919\
        );

    \I__9383\ : InMux
    port map (
            O => \N__41925\,
            I => \N__41916\
        );

    \I__9382\ : LocalMux
    port map (
            O => \N__41922\,
            I => \N__41911\
        );

    \I__9381\ : Span4Mux_h
    port map (
            O => \N__41919\,
            I => \N__41911\
        );

    \I__9380\ : LocalMux
    port map (
            O => \N__41916\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19\
        );

    \I__9379\ : Odrv4
    port map (
            O => \N__41911\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19\
        );

    \I__9378\ : InMux
    port map (
            O => \N__41906\,
            I => \N__41901\
        );

    \I__9377\ : InMux
    port map (
            O => \N__41905\,
            I => \N__41897\
        );

    \I__9376\ : InMux
    port map (
            O => \N__41904\,
            I => \N__41894\
        );

    \I__9375\ : LocalMux
    port map (
            O => \N__41901\,
            I => \N__41891\
        );

    \I__9374\ : InMux
    port map (
            O => \N__41900\,
            I => \N__41888\
        );

    \I__9373\ : LocalMux
    port map (
            O => \N__41897\,
            I => \N__41885\
        );

    \I__9372\ : LocalMux
    port map (
            O => \N__41894\,
            I => \N__41880\
        );

    \I__9371\ : Span4Mux_h
    port map (
            O => \N__41891\,
            I => \N__41880\
        );

    \I__9370\ : LocalMux
    port map (
            O => \N__41888\,
            I => \N__41877\
        );

    \I__9369\ : Span4Mux_h
    port map (
            O => \N__41885\,
            I => \N__41872\
        );

    \I__9368\ : Span4Mux_v
    port map (
            O => \N__41880\,
            I => \N__41872\
        );

    \I__9367\ : Odrv4
    port map (
            O => \N__41877\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__9366\ : Odrv4
    port map (
            O => \N__41872\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__9365\ : CascadeMux
    port map (
            O => \N__41867\,
            I => \N__41864\
        );

    \I__9364\ : InMux
    port map (
            O => \N__41864\,
            I => \N__41858\
        );

    \I__9363\ : InMux
    port map (
            O => \N__41863\,
            I => \N__41858\
        );

    \I__9362\ : LocalMux
    port map (
            O => \N__41858\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\
        );

    \I__9361\ : InMux
    port map (
            O => \N__41855\,
            I => \N__41852\
        );

    \I__9360\ : LocalMux
    port map (
            O => \N__41852\,
            I => \N__41849\
        );

    \I__9359\ : Span4Mux_h
    port map (
            O => \N__41849\,
            I => \N__41846\
        );

    \I__9358\ : Span4Mux_v
    port map (
            O => \N__41846\,
            I => \N__41842\
        );

    \I__9357\ : InMux
    port map (
            O => \N__41845\,
            I => \N__41839\
        );

    \I__9356\ : Odrv4
    port map (
            O => \N__41842\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18\
        );

    \I__9355\ : LocalMux
    port map (
            O => \N__41839\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18\
        );

    \I__9354\ : InMux
    port map (
            O => \N__41834\,
            I => \N__41830\
        );

    \I__9353\ : InMux
    port map (
            O => \N__41833\,
            I => \N__41826\
        );

    \I__9352\ : LocalMux
    port map (
            O => \N__41830\,
            I => \N__41823\
        );

    \I__9351\ : InMux
    port map (
            O => \N__41829\,
            I => \N__41820\
        );

    \I__9350\ : LocalMux
    port map (
            O => \N__41826\,
            I => \elapsed_time_ns_1_RNILK91B_0_9\
        );

    \I__9349\ : Odrv4
    port map (
            O => \N__41823\,
            I => \elapsed_time_ns_1_RNILK91B_0_9\
        );

    \I__9348\ : LocalMux
    port map (
            O => \N__41820\,
            I => \elapsed_time_ns_1_RNILK91B_0_9\
        );

    \I__9347\ : InMux
    port map (
            O => \N__41813\,
            I => \N__41810\
        );

    \I__9346\ : LocalMux
    port map (
            O => \N__41810\,
            I => \N__41805\
        );

    \I__9345\ : InMux
    port map (
            O => \N__41809\,
            I => \N__41802\
        );

    \I__9344\ : InMux
    port map (
            O => \N__41808\,
            I => \N__41799\
        );

    \I__9343\ : Span4Mux_v
    port map (
            O => \N__41805\,
            I => \N__41792\
        );

    \I__9342\ : LocalMux
    port map (
            O => \N__41802\,
            I => \N__41792\
        );

    \I__9341\ : LocalMux
    port map (
            O => \N__41799\,
            I => \N__41792\
        );

    \I__9340\ : Span4Mux_h
    port map (
            O => \N__41792\,
            I => \N__41788\
        );

    \I__9339\ : InMux
    port map (
            O => \N__41791\,
            I => \N__41785\
        );

    \I__9338\ : Odrv4
    port map (
            O => \N__41788\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\
        );

    \I__9337\ : LocalMux
    port map (
            O => \N__41785\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\
        );

    \I__9336\ : CascadeMux
    port map (
            O => \N__41780\,
            I => \N__41777\
        );

    \I__9335\ : InMux
    port map (
            O => \N__41777\,
            I => \N__41774\
        );

    \I__9334\ : LocalMux
    port map (
            O => \N__41774\,
            I => \N__41771\
        );

    \I__9333\ : Span4Mux_v
    port map (
            O => \N__41771\,
            I => \N__41768\
        );

    \I__9332\ : Odrv4
    port map (
            O => \N__41768\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\
        );

    \I__9331\ : InMux
    port map (
            O => \N__41765\,
            I => \N__41761\
        );

    \I__9330\ : InMux
    port map (
            O => \N__41764\,
            I => \N__41758\
        );

    \I__9329\ : LocalMux
    port map (
            O => \N__41761\,
            I => \N__41755\
        );

    \I__9328\ : LocalMux
    port map (
            O => \N__41758\,
            I => \N__41749\
        );

    \I__9327\ : Span4Mux_v
    port map (
            O => \N__41755\,
            I => \N__41749\
        );

    \I__9326\ : InMux
    port map (
            O => \N__41754\,
            I => \N__41746\
        );

    \I__9325\ : Odrv4
    port map (
            O => \N__41749\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17\
        );

    \I__9324\ : LocalMux
    port map (
            O => \N__41746\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17\
        );

    \I__9323\ : CascadeMux
    port map (
            O => \N__41741\,
            I => \N__41735\
        );

    \I__9322\ : CascadeMux
    port map (
            O => \N__41740\,
            I => \N__41732\
        );

    \I__9321\ : InMux
    port map (
            O => \N__41739\,
            I => \N__41729\
        );

    \I__9320\ : InMux
    port map (
            O => \N__41738\,
            I => \N__41726\
        );

    \I__9319\ : InMux
    port map (
            O => \N__41735\,
            I => \N__41723\
        );

    \I__9318\ : InMux
    port map (
            O => \N__41732\,
            I => \N__41720\
        );

    \I__9317\ : LocalMux
    port map (
            O => \N__41729\,
            I => \N__41717\
        );

    \I__9316\ : LocalMux
    port map (
            O => \N__41726\,
            I => \N__41712\
        );

    \I__9315\ : LocalMux
    port map (
            O => \N__41723\,
            I => \N__41712\
        );

    \I__9314\ : LocalMux
    port map (
            O => \N__41720\,
            I => \N__41707\
        );

    \I__9313\ : Span4Mux_h
    port map (
            O => \N__41717\,
            I => \N__41707\
        );

    \I__9312\ : Span4Mux_h
    port map (
            O => \N__41712\,
            I => \N__41704\
        );

    \I__9311\ : Span4Mux_v
    port map (
            O => \N__41707\,
            I => \N__41701\
        );

    \I__9310\ : Span4Mux_v
    port map (
            O => \N__41704\,
            I => \N__41698\
        );

    \I__9309\ : Odrv4
    port map (
            O => \N__41701\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__9308\ : Odrv4
    port map (
            O => \N__41698\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__9307\ : InMux
    port map (
            O => \N__41693\,
            I => \N__41688\
        );

    \I__9306\ : InMux
    port map (
            O => \N__41692\,
            I => \N__41685\
        );

    \I__9305\ : InMux
    port map (
            O => \N__41691\,
            I => \N__41682\
        );

    \I__9304\ : LocalMux
    port map (
            O => \N__41688\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23\
        );

    \I__9303\ : LocalMux
    port map (
            O => \N__41685\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23\
        );

    \I__9302\ : LocalMux
    port map (
            O => \N__41682\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23\
        );

    \I__9301\ : InMux
    port map (
            O => \N__41675\,
            I => \N__41669\
        );

    \I__9300\ : InMux
    port map (
            O => \N__41674\,
            I => \N__41666\
        );

    \I__9299\ : InMux
    port map (
            O => \N__41673\,
            I => \N__41663\
        );

    \I__9298\ : InMux
    port map (
            O => \N__41672\,
            I => \N__41660\
        );

    \I__9297\ : LocalMux
    port map (
            O => \N__41669\,
            I => \N__41657\
        );

    \I__9296\ : LocalMux
    port map (
            O => \N__41666\,
            I => \N__41652\
        );

    \I__9295\ : LocalMux
    port map (
            O => \N__41663\,
            I => \N__41652\
        );

    \I__9294\ : LocalMux
    port map (
            O => \N__41660\,
            I => \N__41649\
        );

    \I__9293\ : Span4Mux_h
    port map (
            O => \N__41657\,
            I => \N__41644\
        );

    \I__9292\ : Span4Mux_v
    port map (
            O => \N__41652\,
            I => \N__41644\
        );

    \I__9291\ : Span4Mux_h
    port map (
            O => \N__41649\,
            I => \N__41641\
        );

    \I__9290\ : Span4Mux_v
    port map (
            O => \N__41644\,
            I => \N__41638\
        );

    \I__9289\ : Span4Mux_v
    port map (
            O => \N__41641\,
            I => \N__41635\
        );

    \I__9288\ : Odrv4
    port map (
            O => \N__41638\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__9287\ : Odrv4
    port map (
            O => \N__41635\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__9286\ : InMux
    port map (
            O => \N__41630\,
            I => \N__41626\
        );

    \I__9285\ : InMux
    port map (
            O => \N__41629\,
            I => \N__41623\
        );

    \I__9284\ : LocalMux
    port map (
            O => \N__41626\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_23\
        );

    \I__9283\ : LocalMux
    port map (
            O => \N__41623\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_23\
        );

    \I__9282\ : CascadeMux
    port map (
            O => \N__41618\,
            I => \N__41615\
        );

    \I__9281\ : InMux
    port map (
            O => \N__41615\,
            I => \N__41612\
        );

    \I__9280\ : LocalMux
    port map (
            O => \N__41612\,
            I => \N__41609\
        );

    \I__9279\ : Span4Mux_v
    port map (
            O => \N__41609\,
            I => \N__41606\
        );

    \I__9278\ : Odrv4
    port map (
            O => \N__41606\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt16\
        );

    \I__9277\ : InMux
    port map (
            O => \N__41603\,
            I => \N__41597\
        );

    \I__9276\ : InMux
    port map (
            O => \N__41602\,
            I => \N__41597\
        );

    \I__9275\ : LocalMux
    port map (
            O => \N__41597\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\
        );

    \I__9274\ : InMux
    port map (
            O => \N__41594\,
            I => \N__41588\
        );

    \I__9273\ : InMux
    port map (
            O => \N__41593\,
            I => \N__41588\
        );

    \I__9272\ : LocalMux
    port map (
            O => \N__41588\,
            I => \N__41584\
        );

    \I__9271\ : InMux
    port map (
            O => \N__41587\,
            I => \N__41581\
        );

    \I__9270\ : Span4Mux_v
    port map (
            O => \N__41584\,
            I => \N__41578\
        );

    \I__9269\ : LocalMux
    port map (
            O => \N__41581\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__9268\ : Odrv4
    port map (
            O => \N__41578\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__9267\ : CascadeMux
    port map (
            O => \N__41573\,
            I => \N__41569\
        );

    \I__9266\ : InMux
    port map (
            O => \N__41572\,
            I => \N__41563\
        );

    \I__9265\ : InMux
    port map (
            O => \N__41569\,
            I => \N__41563\
        );

    \I__9264\ : InMux
    port map (
            O => \N__41568\,
            I => \N__41560\
        );

    \I__9263\ : LocalMux
    port map (
            O => \N__41563\,
            I => \N__41557\
        );

    \I__9262\ : LocalMux
    port map (
            O => \N__41560\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__9261\ : Odrv4
    port map (
            O => \N__41557\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__9260\ : CascadeMux
    port map (
            O => \N__41552\,
            I => \N__41548\
        );

    \I__9259\ : InMux
    port map (
            O => \N__41551\,
            I => \N__41543\
        );

    \I__9258\ : InMux
    port map (
            O => \N__41548\,
            I => \N__41543\
        );

    \I__9257\ : LocalMux
    port map (
            O => \N__41543\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\
        );

    \I__9256\ : InMux
    port map (
            O => \N__41540\,
            I => \N__41537\
        );

    \I__9255\ : LocalMux
    port map (
            O => \N__41537\,
            I => \N__41534\
        );

    \I__9254\ : Span4Mux_v
    port map (
            O => \N__41534\,
            I => \N__41531\
        );

    \I__9253\ : Odrv4
    port map (
            O => \N__41531\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\
        );

    \I__9252\ : InMux
    port map (
            O => \N__41528\,
            I => \N__41525\
        );

    \I__9251\ : LocalMux
    port map (
            O => \N__41525\,
            I => \N__41521\
        );

    \I__9250\ : InMux
    port map (
            O => \N__41524\,
            I => \N__41517\
        );

    \I__9249\ : Span12Mux_h
    port map (
            O => \N__41521\,
            I => \N__41514\
        );

    \I__9248\ : InMux
    port map (
            O => \N__41520\,
            I => \N__41511\
        );

    \I__9247\ : LocalMux
    port map (
            O => \N__41517\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14\
        );

    \I__9246\ : Odrv12
    port map (
            O => \N__41514\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14\
        );

    \I__9245\ : LocalMux
    port map (
            O => \N__41511\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14\
        );

    \I__9244\ : InMux
    port map (
            O => \N__41504\,
            I => \N__41498\
        );

    \I__9243\ : InMux
    port map (
            O => \N__41503\,
            I => \N__41495\
        );

    \I__9242\ : InMux
    port map (
            O => \N__41502\,
            I => \N__41492\
        );

    \I__9241\ : InMux
    port map (
            O => \N__41501\,
            I => \N__41489\
        );

    \I__9240\ : LocalMux
    port map (
            O => \N__41498\,
            I => \N__41484\
        );

    \I__9239\ : LocalMux
    port map (
            O => \N__41495\,
            I => \N__41484\
        );

    \I__9238\ : LocalMux
    port map (
            O => \N__41492\,
            I => \N__41479\
        );

    \I__9237\ : LocalMux
    port map (
            O => \N__41489\,
            I => \N__41479\
        );

    \I__9236\ : Span4Mux_v
    port map (
            O => \N__41484\,
            I => \N__41474\
        );

    \I__9235\ : Span4Mux_v
    port map (
            O => \N__41479\,
            I => \N__41474\
        );

    \I__9234\ : Odrv4
    port map (
            O => \N__41474\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\
        );

    \I__9233\ : InMux
    port map (
            O => \N__41471\,
            I => \N__41468\
        );

    \I__9232\ : LocalMux
    port map (
            O => \N__41468\,
            I => \N__41465\
        );

    \I__9231\ : Span4Mux_h
    port map (
            O => \N__41465\,
            I => \N__41462\
        );

    \I__9230\ : Odrv4
    port map (
            O => \N__41462\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\
        );

    \I__9229\ : InMux
    port map (
            O => \N__41459\,
            I => \N__41456\
        );

    \I__9228\ : LocalMux
    port map (
            O => \N__41456\,
            I => \N__41451\
        );

    \I__9227\ : InMux
    port map (
            O => \N__41455\,
            I => \N__41448\
        );

    \I__9226\ : InMux
    port map (
            O => \N__41454\,
            I => \N__41444\
        );

    \I__9225\ : Span4Mux_v
    port map (
            O => \N__41451\,
            I => \N__41439\
        );

    \I__9224\ : LocalMux
    port map (
            O => \N__41448\,
            I => \N__41439\
        );

    \I__9223\ : InMux
    port map (
            O => \N__41447\,
            I => \N__41436\
        );

    \I__9222\ : LocalMux
    port map (
            O => \N__41444\,
            I => \N__41433\
        );

    \I__9221\ : Span4Mux_v
    port map (
            O => \N__41439\,
            I => \N__41428\
        );

    \I__9220\ : LocalMux
    port map (
            O => \N__41436\,
            I => \N__41428\
        );

    \I__9219\ : Span4Mux_v
    port map (
            O => \N__41433\,
            I => \N__41423\
        );

    \I__9218\ : Span4Mux_h
    port map (
            O => \N__41428\,
            I => \N__41423\
        );

    \I__9217\ : Odrv4
    port map (
            O => \N__41423\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__9216\ : InMux
    port map (
            O => \N__41420\,
            I => \N__41417\
        );

    \I__9215\ : LocalMux
    port map (
            O => \N__41417\,
            I => \N__41412\
        );

    \I__9214\ : InMux
    port map (
            O => \N__41416\,
            I => \N__41409\
        );

    \I__9213\ : InMux
    port map (
            O => \N__41415\,
            I => \N__41406\
        );

    \I__9212\ : Span4Mux_h
    port map (
            O => \N__41412\,
            I => \N__41401\
        );

    \I__9211\ : LocalMux
    port map (
            O => \N__41409\,
            I => \N__41401\
        );

    \I__9210\ : LocalMux
    port map (
            O => \N__41406\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16\
        );

    \I__9209\ : Odrv4
    port map (
            O => \N__41401\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16\
        );

    \I__9208\ : InMux
    port map (
            O => \N__41396\,
            I => \N__41389\
        );

    \I__9207\ : InMux
    port map (
            O => \N__41395\,
            I => \N__41389\
        );

    \I__9206\ : InMux
    port map (
            O => \N__41394\,
            I => \N__41386\
        );

    \I__9205\ : LocalMux
    port map (
            O => \N__41389\,
            I => \N__41383\
        );

    \I__9204\ : LocalMux
    port map (
            O => \N__41386\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__9203\ : Odrv4
    port map (
            O => \N__41383\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__9202\ : InMux
    port map (
            O => \N__41378\,
            I => \current_shift_inst.timer_s1.counter_cry_26\
        );

    \I__9201\ : CascadeMux
    port map (
            O => \N__41375\,
            I => \N__41372\
        );

    \I__9200\ : InMux
    port map (
            O => \N__41372\,
            I => \N__41368\
        );

    \I__9199\ : InMux
    port map (
            O => \N__41371\,
            I => \N__41365\
        );

    \I__9198\ : LocalMux
    port map (
            O => \N__41368\,
            I => \N__41362\
        );

    \I__9197\ : LocalMux
    port map (
            O => \N__41365\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__9196\ : Odrv4
    port map (
            O => \N__41362\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__9195\ : InMux
    port map (
            O => \N__41357\,
            I => \current_shift_inst.timer_s1.counter_cry_27\
        );

    \I__9194\ : InMux
    port map (
            O => \N__41354\,
            I => \N__41316\
        );

    \I__9193\ : InMux
    port map (
            O => \N__41353\,
            I => \N__41316\
        );

    \I__9192\ : InMux
    port map (
            O => \N__41352\,
            I => \N__41316\
        );

    \I__9191\ : InMux
    port map (
            O => \N__41351\,
            I => \N__41316\
        );

    \I__9190\ : InMux
    port map (
            O => \N__41350\,
            I => \N__41307\
        );

    \I__9189\ : InMux
    port map (
            O => \N__41349\,
            I => \N__41307\
        );

    \I__9188\ : InMux
    port map (
            O => \N__41348\,
            I => \N__41307\
        );

    \I__9187\ : InMux
    port map (
            O => \N__41347\,
            I => \N__41307\
        );

    \I__9186\ : InMux
    port map (
            O => \N__41346\,
            I => \N__41302\
        );

    \I__9185\ : InMux
    port map (
            O => \N__41345\,
            I => \N__41302\
        );

    \I__9184\ : InMux
    port map (
            O => \N__41344\,
            I => \N__41293\
        );

    \I__9183\ : InMux
    port map (
            O => \N__41343\,
            I => \N__41293\
        );

    \I__9182\ : InMux
    port map (
            O => \N__41342\,
            I => \N__41293\
        );

    \I__9181\ : InMux
    port map (
            O => \N__41341\,
            I => \N__41293\
        );

    \I__9180\ : InMux
    port map (
            O => \N__41340\,
            I => \N__41284\
        );

    \I__9179\ : InMux
    port map (
            O => \N__41339\,
            I => \N__41284\
        );

    \I__9178\ : InMux
    port map (
            O => \N__41338\,
            I => \N__41284\
        );

    \I__9177\ : InMux
    port map (
            O => \N__41337\,
            I => \N__41284\
        );

    \I__9176\ : InMux
    port map (
            O => \N__41336\,
            I => \N__41275\
        );

    \I__9175\ : InMux
    port map (
            O => \N__41335\,
            I => \N__41275\
        );

    \I__9174\ : InMux
    port map (
            O => \N__41334\,
            I => \N__41275\
        );

    \I__9173\ : InMux
    port map (
            O => \N__41333\,
            I => \N__41275\
        );

    \I__9172\ : InMux
    port map (
            O => \N__41332\,
            I => \N__41266\
        );

    \I__9171\ : InMux
    port map (
            O => \N__41331\,
            I => \N__41266\
        );

    \I__9170\ : InMux
    port map (
            O => \N__41330\,
            I => \N__41266\
        );

    \I__9169\ : InMux
    port map (
            O => \N__41329\,
            I => \N__41266\
        );

    \I__9168\ : InMux
    port map (
            O => \N__41328\,
            I => \N__41257\
        );

    \I__9167\ : InMux
    port map (
            O => \N__41327\,
            I => \N__41257\
        );

    \I__9166\ : InMux
    port map (
            O => \N__41326\,
            I => \N__41257\
        );

    \I__9165\ : InMux
    port map (
            O => \N__41325\,
            I => \N__41257\
        );

    \I__9164\ : LocalMux
    port map (
            O => \N__41316\,
            I => \N__41254\
        );

    \I__9163\ : LocalMux
    port map (
            O => \N__41307\,
            I => \N__41247\
        );

    \I__9162\ : LocalMux
    port map (
            O => \N__41302\,
            I => \N__41247\
        );

    \I__9161\ : LocalMux
    port map (
            O => \N__41293\,
            I => \N__41247\
        );

    \I__9160\ : LocalMux
    port map (
            O => \N__41284\,
            I => \N__41240\
        );

    \I__9159\ : LocalMux
    port map (
            O => \N__41275\,
            I => \N__41240\
        );

    \I__9158\ : LocalMux
    port map (
            O => \N__41266\,
            I => \N__41240\
        );

    \I__9157\ : LocalMux
    port map (
            O => \N__41257\,
            I => \N__41237\
        );

    \I__9156\ : Span4Mux_h
    port map (
            O => \N__41254\,
            I => \N__41234\
        );

    \I__9155\ : Span4Mux_v
    port map (
            O => \N__41247\,
            I => \N__41229\
        );

    \I__9154\ : Span4Mux_v
    port map (
            O => \N__41240\,
            I => \N__41229\
        );

    \I__9153\ : Span4Mux_h
    port map (
            O => \N__41237\,
            I => \N__41224\
        );

    \I__9152\ : Span4Mux_h
    port map (
            O => \N__41234\,
            I => \N__41224\
        );

    \I__9151\ : Odrv4
    port map (
            O => \N__41229\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__9150\ : Odrv4
    port map (
            O => \N__41224\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__9149\ : InMux
    port map (
            O => \N__41219\,
            I => \current_shift_inst.timer_s1.counter_cry_28\
        );

    \I__9148\ : CascadeMux
    port map (
            O => \N__41216\,
            I => \N__41213\
        );

    \I__9147\ : InMux
    port map (
            O => \N__41213\,
            I => \N__41209\
        );

    \I__9146\ : InMux
    port map (
            O => \N__41212\,
            I => \N__41206\
        );

    \I__9145\ : LocalMux
    port map (
            O => \N__41209\,
            I => \N__41203\
        );

    \I__9144\ : LocalMux
    port map (
            O => \N__41206\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__9143\ : Odrv4
    port map (
            O => \N__41203\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__9142\ : CEMux
    port map (
            O => \N__41198\,
            I => \N__41194\
        );

    \I__9141\ : CEMux
    port map (
            O => \N__41197\,
            I => \N__41190\
        );

    \I__9140\ : LocalMux
    port map (
            O => \N__41194\,
            I => \N__41187\
        );

    \I__9139\ : CEMux
    port map (
            O => \N__41193\,
            I => \N__41183\
        );

    \I__9138\ : LocalMux
    port map (
            O => \N__41190\,
            I => \N__41180\
        );

    \I__9137\ : Span4Mux_v
    port map (
            O => \N__41187\,
            I => \N__41177\
        );

    \I__9136\ : CEMux
    port map (
            O => \N__41186\,
            I => \N__41174\
        );

    \I__9135\ : LocalMux
    port map (
            O => \N__41183\,
            I => \N__41171\
        );

    \I__9134\ : Span4Mux_v
    port map (
            O => \N__41180\,
            I => \N__41168\
        );

    \I__9133\ : Span4Mux_h
    port map (
            O => \N__41177\,
            I => \N__41163\
        );

    \I__9132\ : LocalMux
    port map (
            O => \N__41174\,
            I => \N__41163\
        );

    \I__9131\ : Span4Mux_h
    port map (
            O => \N__41171\,
            I => \N__41160\
        );

    \I__9130\ : Span4Mux_h
    port map (
            O => \N__41168\,
            I => \N__41155\
        );

    \I__9129\ : Span4Mux_h
    port map (
            O => \N__41163\,
            I => \N__41155\
        );

    \I__9128\ : Odrv4
    port map (
            O => \N__41160\,
            I => \current_shift_inst.timer_s1.N_163_i\
        );

    \I__9127\ : Odrv4
    port map (
            O => \N__41155\,
            I => \current_shift_inst.timer_s1.N_163_i\
        );

    \I__9126\ : InMux
    port map (
            O => \N__41150\,
            I => \N__41144\
        );

    \I__9125\ : InMux
    port map (
            O => \N__41149\,
            I => \N__41141\
        );

    \I__9124\ : InMux
    port map (
            O => \N__41148\,
            I => \N__41136\
        );

    \I__9123\ : InMux
    port map (
            O => \N__41147\,
            I => \N__41136\
        );

    \I__9122\ : LocalMux
    port map (
            O => \N__41144\,
            I => \N__41133\
        );

    \I__9121\ : LocalMux
    port map (
            O => \N__41141\,
            I => \N__41128\
        );

    \I__9120\ : LocalMux
    port map (
            O => \N__41136\,
            I => \N__41128\
        );

    \I__9119\ : Span4Mux_v
    port map (
            O => \N__41133\,
            I => \N__41125\
        );

    \I__9118\ : Span4Mux_h
    port map (
            O => \N__41128\,
            I => \N__41122\
        );

    \I__9117\ : Span4Mux_h
    port map (
            O => \N__41125\,
            I => \N__41119\
        );

    \I__9116\ : Odrv4
    port map (
            O => \N__41122\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__9115\ : Odrv4
    port map (
            O => \N__41119\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__9114\ : InMux
    port map (
            O => \N__41114\,
            I => \N__41106\
        );

    \I__9113\ : InMux
    port map (
            O => \N__41113\,
            I => \N__41106\
        );

    \I__9112\ : InMux
    port map (
            O => \N__41112\,
            I => \N__41103\
        );

    \I__9111\ : InMux
    port map (
            O => \N__41111\,
            I => \N__41100\
        );

    \I__9110\ : LocalMux
    port map (
            O => \N__41106\,
            I => \N__41097\
        );

    \I__9109\ : LocalMux
    port map (
            O => \N__41103\,
            I => \N__41094\
        );

    \I__9108\ : LocalMux
    port map (
            O => \N__41100\,
            I => \N__41091\
        );

    \I__9107\ : Span4Mux_v
    port map (
            O => \N__41097\,
            I => \N__41088\
        );

    \I__9106\ : Span4Mux_v
    port map (
            O => \N__41094\,
            I => \N__41085\
        );

    \I__9105\ : Span4Mux_v
    port map (
            O => \N__41091\,
            I => \N__41082\
        );

    \I__9104\ : Span4Mux_v
    port map (
            O => \N__41088\,
            I => \N__41079\
        );

    \I__9103\ : Span4Mux_h
    port map (
            O => \N__41085\,
            I => \N__41076\
        );

    \I__9102\ : Odrv4
    port map (
            O => \N__41082\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__9101\ : Odrv4
    port map (
            O => \N__41079\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__9100\ : Odrv4
    port map (
            O => \N__41076\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__9099\ : InMux
    port map (
            O => \N__41069\,
            I => \N__41066\
        );

    \I__9098\ : LocalMux
    port map (
            O => \N__41066\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20\
        );

    \I__9097\ : InMux
    port map (
            O => \N__41063\,
            I => \N__41059\
        );

    \I__9096\ : InMux
    port map (
            O => \N__41062\,
            I => \N__41056\
        );

    \I__9095\ : LocalMux
    port map (
            O => \N__41059\,
            I => \N__41053\
        );

    \I__9094\ : LocalMux
    port map (
            O => \N__41056\,
            I => \N__41050\
        );

    \I__9093\ : Span4Mux_h
    port map (
            O => \N__41053\,
            I => \N__41047\
        );

    \I__9092\ : Span4Mux_v
    port map (
            O => \N__41050\,
            I => \N__41042\
        );

    \I__9091\ : Span4Mux_h
    port map (
            O => \N__41047\,
            I => \N__41039\
        );

    \I__9090\ : InMux
    port map (
            O => \N__41046\,
            I => \N__41034\
        );

    \I__9089\ : InMux
    port map (
            O => \N__41045\,
            I => \N__41034\
        );

    \I__9088\ : Span4Mux_h
    port map (
            O => \N__41042\,
            I => \N__41031\
        );

    \I__9087\ : Odrv4
    port map (
            O => \N__41039\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__9086\ : LocalMux
    port map (
            O => \N__41034\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__9085\ : Odrv4
    port map (
            O => \N__41031\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__9084\ : InMux
    port map (
            O => \N__41024\,
            I => \N__41021\
        );

    \I__9083\ : LocalMux
    port map (
            O => \N__41021\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21\
        );

    \I__9082\ : InMux
    port map (
            O => \N__41018\,
            I => \N__41011\
        );

    \I__9081\ : InMux
    port map (
            O => \N__41017\,
            I => \N__41011\
        );

    \I__9080\ : InMux
    port map (
            O => \N__41016\,
            I => \N__41008\
        );

    \I__9079\ : LocalMux
    port map (
            O => \N__41011\,
            I => \N__41005\
        );

    \I__9078\ : LocalMux
    port map (
            O => \N__41008\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__9077\ : Odrv12
    port map (
            O => \N__41005\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__9076\ : InMux
    port map (
            O => \N__41000\,
            I => \current_shift_inst.timer_s1.counter_cry_17\
        );

    \I__9075\ : CascadeMux
    port map (
            O => \N__40997\,
            I => \N__40994\
        );

    \I__9074\ : InMux
    port map (
            O => \N__40994\,
            I => \N__40989\
        );

    \I__9073\ : InMux
    port map (
            O => \N__40993\,
            I => \N__40986\
        );

    \I__9072\ : InMux
    port map (
            O => \N__40992\,
            I => \N__40983\
        );

    \I__9071\ : LocalMux
    port map (
            O => \N__40989\,
            I => \N__40978\
        );

    \I__9070\ : LocalMux
    port map (
            O => \N__40986\,
            I => \N__40978\
        );

    \I__9069\ : LocalMux
    port map (
            O => \N__40983\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__9068\ : Odrv12
    port map (
            O => \N__40978\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__9067\ : InMux
    port map (
            O => \N__40973\,
            I => \current_shift_inst.timer_s1.counter_cry_18\
        );

    \I__9066\ : CascadeMux
    port map (
            O => \N__40970\,
            I => \N__40966\
        );

    \I__9065\ : CascadeMux
    port map (
            O => \N__40969\,
            I => \N__40963\
        );

    \I__9064\ : InMux
    port map (
            O => \N__40966\,
            I => \N__40957\
        );

    \I__9063\ : InMux
    port map (
            O => \N__40963\,
            I => \N__40957\
        );

    \I__9062\ : InMux
    port map (
            O => \N__40962\,
            I => \N__40954\
        );

    \I__9061\ : LocalMux
    port map (
            O => \N__40957\,
            I => \N__40951\
        );

    \I__9060\ : LocalMux
    port map (
            O => \N__40954\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__9059\ : Odrv4
    port map (
            O => \N__40951\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__9058\ : InMux
    port map (
            O => \N__40946\,
            I => \current_shift_inst.timer_s1.counter_cry_19\
        );

    \I__9057\ : InMux
    port map (
            O => \N__40943\,
            I => \N__40936\
        );

    \I__9056\ : InMux
    port map (
            O => \N__40942\,
            I => \N__40936\
        );

    \I__9055\ : InMux
    port map (
            O => \N__40941\,
            I => \N__40933\
        );

    \I__9054\ : LocalMux
    port map (
            O => \N__40936\,
            I => \N__40930\
        );

    \I__9053\ : LocalMux
    port map (
            O => \N__40933\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__9052\ : Odrv12
    port map (
            O => \N__40930\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__9051\ : InMux
    port map (
            O => \N__40925\,
            I => \current_shift_inst.timer_s1.counter_cry_20\
        );

    \I__9050\ : InMux
    port map (
            O => \N__40922\,
            I => \N__40915\
        );

    \I__9049\ : InMux
    port map (
            O => \N__40921\,
            I => \N__40915\
        );

    \I__9048\ : InMux
    port map (
            O => \N__40920\,
            I => \N__40912\
        );

    \I__9047\ : LocalMux
    port map (
            O => \N__40915\,
            I => \N__40909\
        );

    \I__9046\ : LocalMux
    port map (
            O => \N__40912\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__9045\ : Odrv4
    port map (
            O => \N__40909\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__9044\ : InMux
    port map (
            O => \N__40904\,
            I => \current_shift_inst.timer_s1.counter_cry_21\
        );

    \I__9043\ : CascadeMux
    port map (
            O => \N__40901\,
            I => \N__40897\
        );

    \I__9042\ : CascadeMux
    port map (
            O => \N__40900\,
            I => \N__40894\
        );

    \I__9041\ : InMux
    port map (
            O => \N__40897\,
            I => \N__40888\
        );

    \I__9040\ : InMux
    port map (
            O => \N__40894\,
            I => \N__40888\
        );

    \I__9039\ : InMux
    port map (
            O => \N__40893\,
            I => \N__40885\
        );

    \I__9038\ : LocalMux
    port map (
            O => \N__40888\,
            I => \N__40882\
        );

    \I__9037\ : LocalMux
    port map (
            O => \N__40885\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__9036\ : Odrv4
    port map (
            O => \N__40882\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__9035\ : InMux
    port map (
            O => \N__40877\,
            I => \current_shift_inst.timer_s1.counter_cry_22\
        );

    \I__9034\ : CascadeMux
    port map (
            O => \N__40874\,
            I => \N__40870\
        );

    \I__9033\ : CascadeMux
    port map (
            O => \N__40873\,
            I => \N__40867\
        );

    \I__9032\ : InMux
    port map (
            O => \N__40870\,
            I => \N__40864\
        );

    \I__9031\ : InMux
    port map (
            O => \N__40867\,
            I => \N__40860\
        );

    \I__9030\ : LocalMux
    port map (
            O => \N__40864\,
            I => \N__40857\
        );

    \I__9029\ : InMux
    port map (
            O => \N__40863\,
            I => \N__40854\
        );

    \I__9028\ : LocalMux
    port map (
            O => \N__40860\,
            I => \N__40851\
        );

    \I__9027\ : Span4Mux_v
    port map (
            O => \N__40857\,
            I => \N__40848\
        );

    \I__9026\ : LocalMux
    port map (
            O => \N__40854\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__9025\ : Odrv12
    port map (
            O => \N__40851\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__9024\ : Odrv4
    port map (
            O => \N__40848\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__9023\ : InMux
    port map (
            O => \N__40841\,
            I => \bfn_17_21_0_\
        );

    \I__9022\ : CascadeMux
    port map (
            O => \N__40838\,
            I => \N__40834\
        );

    \I__9021\ : InMux
    port map (
            O => \N__40837\,
            I => \N__40831\
        );

    \I__9020\ : InMux
    port map (
            O => \N__40834\,
            I => \N__40827\
        );

    \I__9019\ : LocalMux
    port map (
            O => \N__40831\,
            I => \N__40824\
        );

    \I__9018\ : InMux
    port map (
            O => \N__40830\,
            I => \N__40821\
        );

    \I__9017\ : LocalMux
    port map (
            O => \N__40827\,
            I => \N__40818\
        );

    \I__9016\ : Span4Mux_v
    port map (
            O => \N__40824\,
            I => \N__40815\
        );

    \I__9015\ : LocalMux
    port map (
            O => \N__40821\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__9014\ : Odrv12
    port map (
            O => \N__40818\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__9013\ : Odrv4
    port map (
            O => \N__40815\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__9012\ : InMux
    port map (
            O => \N__40808\,
            I => \current_shift_inst.timer_s1.counter_cry_24\
        );

    \I__9011\ : InMux
    port map (
            O => \N__40805\,
            I => \N__40798\
        );

    \I__9010\ : InMux
    port map (
            O => \N__40804\,
            I => \N__40798\
        );

    \I__9009\ : InMux
    port map (
            O => \N__40803\,
            I => \N__40795\
        );

    \I__9008\ : LocalMux
    port map (
            O => \N__40798\,
            I => \N__40792\
        );

    \I__9007\ : LocalMux
    port map (
            O => \N__40795\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__9006\ : Odrv4
    port map (
            O => \N__40792\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__9005\ : InMux
    port map (
            O => \N__40787\,
            I => \current_shift_inst.timer_s1.counter_cry_25\
        );

    \I__9004\ : InMux
    port map (
            O => \N__40784\,
            I => \N__40777\
        );

    \I__9003\ : InMux
    port map (
            O => \N__40783\,
            I => \N__40777\
        );

    \I__9002\ : InMux
    port map (
            O => \N__40782\,
            I => \N__40774\
        );

    \I__9001\ : LocalMux
    port map (
            O => \N__40777\,
            I => \N__40771\
        );

    \I__9000\ : LocalMux
    port map (
            O => \N__40774\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__8999\ : Odrv4
    port map (
            O => \N__40771\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__8998\ : InMux
    port map (
            O => \N__40766\,
            I => \current_shift_inst.timer_s1.counter_cry_9\
        );

    \I__8997\ : InMux
    port map (
            O => \N__40763\,
            I => \N__40756\
        );

    \I__8996\ : InMux
    port map (
            O => \N__40762\,
            I => \N__40756\
        );

    \I__8995\ : InMux
    port map (
            O => \N__40761\,
            I => \N__40753\
        );

    \I__8994\ : LocalMux
    port map (
            O => \N__40756\,
            I => \N__40750\
        );

    \I__8993\ : LocalMux
    port map (
            O => \N__40753\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__8992\ : Odrv4
    port map (
            O => \N__40750\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__8991\ : InMux
    port map (
            O => \N__40745\,
            I => \current_shift_inst.timer_s1.counter_cry_10\
        );

    \I__8990\ : CascadeMux
    port map (
            O => \N__40742\,
            I => \N__40738\
        );

    \I__8989\ : InMux
    port map (
            O => \N__40741\,
            I => \N__40734\
        );

    \I__8988\ : InMux
    port map (
            O => \N__40738\,
            I => \N__40731\
        );

    \I__8987\ : InMux
    port map (
            O => \N__40737\,
            I => \N__40728\
        );

    \I__8986\ : LocalMux
    port map (
            O => \N__40734\,
            I => \N__40723\
        );

    \I__8985\ : LocalMux
    port map (
            O => \N__40731\,
            I => \N__40723\
        );

    \I__8984\ : LocalMux
    port map (
            O => \N__40728\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__8983\ : Odrv4
    port map (
            O => \N__40723\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__8982\ : InMux
    port map (
            O => \N__40718\,
            I => \current_shift_inst.timer_s1.counter_cry_11\
        );

    \I__8981\ : CascadeMux
    port map (
            O => \N__40715\,
            I => \N__40711\
        );

    \I__8980\ : InMux
    port map (
            O => \N__40714\,
            I => \N__40707\
        );

    \I__8979\ : InMux
    port map (
            O => \N__40711\,
            I => \N__40704\
        );

    \I__8978\ : InMux
    port map (
            O => \N__40710\,
            I => \N__40701\
        );

    \I__8977\ : LocalMux
    port map (
            O => \N__40707\,
            I => \N__40696\
        );

    \I__8976\ : LocalMux
    port map (
            O => \N__40704\,
            I => \N__40696\
        );

    \I__8975\ : LocalMux
    port map (
            O => \N__40701\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__8974\ : Odrv4
    port map (
            O => \N__40696\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__8973\ : InMux
    port map (
            O => \N__40691\,
            I => \current_shift_inst.timer_s1.counter_cry_12\
        );

    \I__8972\ : CascadeMux
    port map (
            O => \N__40688\,
            I => \N__40684\
        );

    \I__8971\ : CascadeMux
    port map (
            O => \N__40687\,
            I => \N__40681\
        );

    \I__8970\ : InMux
    port map (
            O => \N__40684\,
            I => \N__40675\
        );

    \I__8969\ : InMux
    port map (
            O => \N__40681\,
            I => \N__40675\
        );

    \I__8968\ : InMux
    port map (
            O => \N__40680\,
            I => \N__40672\
        );

    \I__8967\ : LocalMux
    port map (
            O => \N__40675\,
            I => \N__40669\
        );

    \I__8966\ : LocalMux
    port map (
            O => \N__40672\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__8965\ : Odrv4
    port map (
            O => \N__40669\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__8964\ : InMux
    port map (
            O => \N__40664\,
            I => \current_shift_inst.timer_s1.counter_cry_13\
        );

    \I__8963\ : CascadeMux
    port map (
            O => \N__40661\,
            I => \N__40657\
        );

    \I__8962\ : CascadeMux
    port map (
            O => \N__40660\,
            I => \N__40654\
        );

    \I__8961\ : InMux
    port map (
            O => \N__40657\,
            I => \N__40648\
        );

    \I__8960\ : InMux
    port map (
            O => \N__40654\,
            I => \N__40648\
        );

    \I__8959\ : InMux
    port map (
            O => \N__40653\,
            I => \N__40645\
        );

    \I__8958\ : LocalMux
    port map (
            O => \N__40648\,
            I => \N__40642\
        );

    \I__8957\ : LocalMux
    port map (
            O => \N__40645\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__8956\ : Odrv4
    port map (
            O => \N__40642\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__8955\ : InMux
    port map (
            O => \N__40637\,
            I => \current_shift_inst.timer_s1.counter_cry_14\
        );

    \I__8954\ : CascadeMux
    port map (
            O => \N__40634\,
            I => \N__40630\
        );

    \I__8953\ : InMux
    port map (
            O => \N__40633\,
            I => \N__40627\
        );

    \I__8952\ : InMux
    port map (
            O => \N__40630\,
            I => \N__40623\
        );

    \I__8951\ : LocalMux
    port map (
            O => \N__40627\,
            I => \N__40620\
        );

    \I__8950\ : InMux
    port map (
            O => \N__40626\,
            I => \N__40617\
        );

    \I__8949\ : LocalMux
    port map (
            O => \N__40623\,
            I => \N__40614\
        );

    \I__8948\ : Span4Mux_v
    port map (
            O => \N__40620\,
            I => \N__40611\
        );

    \I__8947\ : LocalMux
    port map (
            O => \N__40617\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__8946\ : Odrv12
    port map (
            O => \N__40614\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__8945\ : Odrv4
    port map (
            O => \N__40611\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__8944\ : InMux
    port map (
            O => \N__40604\,
            I => \bfn_17_20_0_\
        );

    \I__8943\ : CascadeMux
    port map (
            O => \N__40601\,
            I => \N__40597\
        );

    \I__8942\ : InMux
    port map (
            O => \N__40600\,
            I => \N__40594\
        );

    \I__8941\ : InMux
    port map (
            O => \N__40597\,
            I => \N__40591\
        );

    \I__8940\ : LocalMux
    port map (
            O => \N__40594\,
            I => \N__40588\
        );

    \I__8939\ : LocalMux
    port map (
            O => \N__40591\,
            I => \N__40582\
        );

    \I__8938\ : Span4Mux_v
    port map (
            O => \N__40588\,
            I => \N__40582\
        );

    \I__8937\ : InMux
    port map (
            O => \N__40587\,
            I => \N__40579\
        );

    \I__8936\ : Span4Mux_h
    port map (
            O => \N__40582\,
            I => \N__40576\
        );

    \I__8935\ : LocalMux
    port map (
            O => \N__40579\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__8934\ : Odrv4
    port map (
            O => \N__40576\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__8933\ : InMux
    port map (
            O => \N__40571\,
            I => \current_shift_inst.timer_s1.counter_cry_16\
        );

    \I__8932\ : InMux
    port map (
            O => \N__40568\,
            I => \N__40561\
        );

    \I__8931\ : InMux
    port map (
            O => \N__40567\,
            I => \N__40561\
        );

    \I__8930\ : InMux
    port map (
            O => \N__40566\,
            I => \N__40558\
        );

    \I__8929\ : LocalMux
    port map (
            O => \N__40561\,
            I => \N__40555\
        );

    \I__8928\ : LocalMux
    port map (
            O => \N__40558\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__8927\ : Odrv12
    port map (
            O => \N__40555\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__8926\ : InMux
    port map (
            O => \N__40550\,
            I => \current_shift_inst.timer_s1.counter_cry_1\
        );

    \I__8925\ : CascadeMux
    port map (
            O => \N__40547\,
            I => \N__40543\
        );

    \I__8924\ : InMux
    port map (
            O => \N__40546\,
            I => \N__40540\
        );

    \I__8923\ : InMux
    port map (
            O => \N__40543\,
            I => \N__40537\
        );

    \I__8922\ : LocalMux
    port map (
            O => \N__40540\,
            I => \N__40531\
        );

    \I__8921\ : LocalMux
    port map (
            O => \N__40537\,
            I => \N__40531\
        );

    \I__8920\ : InMux
    port map (
            O => \N__40536\,
            I => \N__40528\
        );

    \I__8919\ : Span4Mux_h
    port map (
            O => \N__40531\,
            I => \N__40525\
        );

    \I__8918\ : LocalMux
    port map (
            O => \N__40528\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__8917\ : Odrv4
    port map (
            O => \N__40525\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__8916\ : InMux
    port map (
            O => \N__40520\,
            I => \current_shift_inst.timer_s1.counter_cry_2\
        );

    \I__8915\ : CascadeMux
    port map (
            O => \N__40517\,
            I => \N__40513\
        );

    \I__8914\ : CascadeMux
    port map (
            O => \N__40516\,
            I => \N__40510\
        );

    \I__8913\ : InMux
    port map (
            O => \N__40513\,
            I => \N__40504\
        );

    \I__8912\ : InMux
    port map (
            O => \N__40510\,
            I => \N__40504\
        );

    \I__8911\ : InMux
    port map (
            O => \N__40509\,
            I => \N__40501\
        );

    \I__8910\ : LocalMux
    port map (
            O => \N__40504\,
            I => \N__40498\
        );

    \I__8909\ : LocalMux
    port map (
            O => \N__40501\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__8908\ : Odrv4
    port map (
            O => \N__40498\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__8907\ : InMux
    port map (
            O => \N__40493\,
            I => \current_shift_inst.timer_s1.counter_cry_3\
        );

    \I__8906\ : CascadeMux
    port map (
            O => \N__40490\,
            I => \N__40486\
        );

    \I__8905\ : CascadeMux
    port map (
            O => \N__40489\,
            I => \N__40483\
        );

    \I__8904\ : InMux
    port map (
            O => \N__40486\,
            I => \N__40477\
        );

    \I__8903\ : InMux
    port map (
            O => \N__40483\,
            I => \N__40477\
        );

    \I__8902\ : InMux
    port map (
            O => \N__40482\,
            I => \N__40474\
        );

    \I__8901\ : LocalMux
    port map (
            O => \N__40477\,
            I => \N__40471\
        );

    \I__8900\ : LocalMux
    port map (
            O => \N__40474\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__8899\ : Odrv4
    port map (
            O => \N__40471\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__8898\ : InMux
    port map (
            O => \N__40466\,
            I => \current_shift_inst.timer_s1.counter_cry_4\
        );

    \I__8897\ : InMux
    port map (
            O => \N__40463\,
            I => \N__40456\
        );

    \I__8896\ : InMux
    port map (
            O => \N__40462\,
            I => \N__40456\
        );

    \I__8895\ : InMux
    port map (
            O => \N__40461\,
            I => \N__40453\
        );

    \I__8894\ : LocalMux
    port map (
            O => \N__40456\,
            I => \N__40450\
        );

    \I__8893\ : LocalMux
    port map (
            O => \N__40453\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__8892\ : Odrv4
    port map (
            O => \N__40450\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__8891\ : InMux
    port map (
            O => \N__40445\,
            I => \current_shift_inst.timer_s1.counter_cry_5\
        );

    \I__8890\ : InMux
    port map (
            O => \N__40442\,
            I => \N__40435\
        );

    \I__8889\ : InMux
    port map (
            O => \N__40441\,
            I => \N__40435\
        );

    \I__8888\ : InMux
    port map (
            O => \N__40440\,
            I => \N__40432\
        );

    \I__8887\ : LocalMux
    port map (
            O => \N__40435\,
            I => \N__40429\
        );

    \I__8886\ : LocalMux
    port map (
            O => \N__40432\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__8885\ : Odrv4
    port map (
            O => \N__40429\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__8884\ : InMux
    port map (
            O => \N__40424\,
            I => \current_shift_inst.timer_s1.counter_cry_6\
        );

    \I__8883\ : CascadeMux
    port map (
            O => \N__40421\,
            I => \N__40417\
        );

    \I__8882\ : CascadeMux
    port map (
            O => \N__40420\,
            I => \N__40414\
        );

    \I__8881\ : InMux
    port map (
            O => \N__40417\,
            I => \N__40410\
        );

    \I__8880\ : InMux
    port map (
            O => \N__40414\,
            I => \N__40407\
        );

    \I__8879\ : InMux
    port map (
            O => \N__40413\,
            I => \N__40404\
        );

    \I__8878\ : LocalMux
    port map (
            O => \N__40410\,
            I => \N__40399\
        );

    \I__8877\ : LocalMux
    port map (
            O => \N__40407\,
            I => \N__40399\
        );

    \I__8876\ : LocalMux
    port map (
            O => \N__40404\,
            I => \N__40394\
        );

    \I__8875\ : Span4Mux_v
    port map (
            O => \N__40399\,
            I => \N__40394\
        );

    \I__8874\ : Odrv4
    port map (
            O => \N__40394\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__8873\ : InMux
    port map (
            O => \N__40391\,
            I => \bfn_17_19_0_\
        );

    \I__8872\ : CascadeMux
    port map (
            O => \N__40388\,
            I => \N__40384\
        );

    \I__8871\ : CascadeMux
    port map (
            O => \N__40387\,
            I => \N__40381\
        );

    \I__8870\ : InMux
    port map (
            O => \N__40384\,
            I => \N__40378\
        );

    \I__8869\ : InMux
    port map (
            O => \N__40381\,
            I => \N__40375\
        );

    \I__8868\ : LocalMux
    port map (
            O => \N__40378\,
            I => \N__40371\
        );

    \I__8867\ : LocalMux
    port map (
            O => \N__40375\,
            I => \N__40368\
        );

    \I__8866\ : InMux
    port map (
            O => \N__40374\,
            I => \N__40365\
        );

    \I__8865\ : Span4Mux_h
    port map (
            O => \N__40371\,
            I => \N__40360\
        );

    \I__8864\ : Span4Mux_v
    port map (
            O => \N__40368\,
            I => \N__40360\
        );

    \I__8863\ : LocalMux
    port map (
            O => \N__40365\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__8862\ : Odrv4
    port map (
            O => \N__40360\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__8861\ : InMux
    port map (
            O => \N__40355\,
            I => \current_shift_inst.timer_s1.counter_cry_8\
        );

    \I__8860\ : CascadeMux
    port map (
            O => \N__40352\,
            I => \N__40349\
        );

    \I__8859\ : InMux
    port map (
            O => \N__40349\,
            I => \N__40344\
        );

    \I__8858\ : InMux
    port map (
            O => \N__40348\,
            I => \N__40341\
        );

    \I__8857\ : InMux
    port map (
            O => \N__40347\,
            I => \N__40338\
        );

    \I__8856\ : LocalMux
    port map (
            O => \N__40344\,
            I => \N__40335\
        );

    \I__8855\ : LocalMux
    port map (
            O => \N__40341\,
            I => \N__40332\
        );

    \I__8854\ : LocalMux
    port map (
            O => \N__40338\,
            I => \N__40329\
        );

    \I__8853\ : Span4Mux_v
    port map (
            O => \N__40335\,
            I => \N__40323\
        );

    \I__8852\ : Span4Mux_h
    port map (
            O => \N__40332\,
            I => \N__40323\
        );

    \I__8851\ : Span4Mux_h
    port map (
            O => \N__40329\,
            I => \N__40320\
        );

    \I__8850\ : InMux
    port map (
            O => \N__40328\,
            I => \N__40317\
        );

    \I__8849\ : Odrv4
    port map (
            O => \N__40323\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__8848\ : Odrv4
    port map (
            O => \N__40320\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__8847\ : LocalMux
    port map (
            O => \N__40317\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__8846\ : InMux
    port map (
            O => \N__40310\,
            I => \N__40307\
        );

    \I__8845\ : LocalMux
    port map (
            O => \N__40307\,
            I => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\
        );

    \I__8844\ : InMux
    port map (
            O => \N__40304\,
            I => \N__40297\
        );

    \I__8843\ : InMux
    port map (
            O => \N__40303\,
            I => \N__40297\
        );

    \I__8842\ : InMux
    port map (
            O => \N__40302\,
            I => \N__40294\
        );

    \I__8841\ : LocalMux
    port map (
            O => \N__40297\,
            I => \N__40289\
        );

    \I__8840\ : LocalMux
    port map (
            O => \N__40294\,
            I => \N__40289\
        );

    \I__8839\ : Span4Mux_h
    port map (
            O => \N__40289\,
            I => \N__40285\
        );

    \I__8838\ : InMux
    port map (
            O => \N__40288\,
            I => \N__40282\
        );

    \I__8837\ : Odrv4
    port map (
            O => \N__40285\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__8836\ : LocalMux
    port map (
            O => \N__40282\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__8835\ : CascadeMux
    port map (
            O => \N__40277\,
            I => \N__40274\
        );

    \I__8834\ : InMux
    port map (
            O => \N__40274\,
            I => \N__40271\
        );

    \I__8833\ : LocalMux
    port map (
            O => \N__40271\,
            I => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\
        );

    \I__8832\ : InMux
    port map (
            O => \N__40268\,
            I => \N__40265\
        );

    \I__8831\ : LocalMux
    port map (
            O => \N__40265\,
            I => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\
        );

    \I__8830\ : InMux
    port map (
            O => \N__40262\,
            I => \N__40255\
        );

    \I__8829\ : InMux
    port map (
            O => \N__40261\,
            I => \N__40255\
        );

    \I__8828\ : InMux
    port map (
            O => \N__40260\,
            I => \N__40252\
        );

    \I__8827\ : LocalMux
    port map (
            O => \N__40255\,
            I => \N__40249\
        );

    \I__8826\ : LocalMux
    port map (
            O => \N__40252\,
            I => \N__40245\
        );

    \I__8825\ : Span4Mux_h
    port map (
            O => \N__40249\,
            I => \N__40242\
        );

    \I__8824\ : InMux
    port map (
            O => \N__40248\,
            I => \N__40239\
        );

    \I__8823\ : Odrv12
    port map (
            O => \N__40245\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__8822\ : Odrv4
    port map (
            O => \N__40242\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__8821\ : LocalMux
    port map (
            O => \N__40239\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__8820\ : CascadeMux
    port map (
            O => \N__40232\,
            I => \N__40229\
        );

    \I__8819\ : InMux
    port map (
            O => \N__40229\,
            I => \N__40226\
        );

    \I__8818\ : LocalMux
    port map (
            O => \N__40226\,
            I => \N__40223\
        );

    \I__8817\ : Span4Mux_v
    port map (
            O => \N__40223\,
            I => \N__40220\
        );

    \I__8816\ : Span4Mux_h
    port map (
            O => \N__40220\,
            I => \N__40217\
        );

    \I__8815\ : Odrv4
    port map (
            O => \N__40217\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\
        );

    \I__8814\ : InMux
    port map (
            O => \N__40214\,
            I => \N__40211\
        );

    \I__8813\ : LocalMux
    port map (
            O => \N__40211\,
            I => \N__40208\
        );

    \I__8812\ : Odrv12
    port map (
            O => \N__40208\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\
        );

    \I__8811\ : InMux
    port map (
            O => \N__40205\,
            I => \N__40202\
        );

    \I__8810\ : LocalMux
    port map (
            O => \N__40202\,
            I => \N__40199\
        );

    \I__8809\ : Span4Mux_h
    port map (
            O => \N__40199\,
            I => \N__40196\
        );

    \I__8808\ : Odrv4
    port map (
            O => \N__40196\,
            I => \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0\
        );

    \I__8807\ : InMux
    port map (
            O => \N__40193\,
            I => \N__40188\
        );

    \I__8806\ : InMux
    port map (
            O => \N__40192\,
            I => \N__40185\
        );

    \I__8805\ : InMux
    port map (
            O => \N__40191\,
            I => \N__40182\
        );

    \I__8804\ : LocalMux
    port map (
            O => \N__40188\,
            I => \N__40179\
        );

    \I__8803\ : LocalMux
    port map (
            O => \N__40185\,
            I => \N__40175\
        );

    \I__8802\ : LocalMux
    port map (
            O => \N__40182\,
            I => \N__40170\
        );

    \I__8801\ : Span4Mux_h
    port map (
            O => \N__40179\,
            I => \N__40170\
        );

    \I__8800\ : InMux
    port map (
            O => \N__40178\,
            I => \N__40167\
        );

    \I__8799\ : Odrv12
    port map (
            O => \N__40175\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__8798\ : Odrv4
    port map (
            O => \N__40170\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__8797\ : LocalMux
    port map (
            O => \N__40167\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__8796\ : InMux
    port map (
            O => \N__40160\,
            I => \N__40157\
        );

    \I__8795\ : LocalMux
    port map (
            O => \N__40157\,
            I => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\
        );

    \I__8794\ : InMux
    port map (
            O => \N__40154\,
            I => \N__40150\
        );

    \I__8793\ : CascadeMux
    port map (
            O => \N__40153\,
            I => \N__40147\
        );

    \I__8792\ : LocalMux
    port map (
            O => \N__40150\,
            I => \N__40143\
        );

    \I__8791\ : InMux
    port map (
            O => \N__40147\,
            I => \N__40140\
        );

    \I__8790\ : InMux
    port map (
            O => \N__40146\,
            I => \N__40137\
        );

    \I__8789\ : Span12Mux_v
    port map (
            O => \N__40143\,
            I => \N__40132\
        );

    \I__8788\ : LocalMux
    port map (
            O => \N__40140\,
            I => \N__40132\
        );

    \I__8787\ : LocalMux
    port map (
            O => \N__40137\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__8786\ : Odrv12
    port map (
            O => \N__40132\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__8785\ : InMux
    port map (
            O => \N__40127\,
            I => \bfn_17_18_0_\
        );

    \I__8784\ : InMux
    port map (
            O => \N__40124\,
            I => \current_shift_inst.timer_s1.counter_cry_0\
        );

    \I__8783\ : CascadeMux
    port map (
            O => \N__40121\,
            I => \N__40117\
        );

    \I__8782\ : InMux
    port map (
            O => \N__40120\,
            I => \N__40114\
        );

    \I__8781\ : InMux
    port map (
            O => \N__40117\,
            I => \N__40110\
        );

    \I__8780\ : LocalMux
    port map (
            O => \N__40114\,
            I => \N__40107\
        );

    \I__8779\ : InMux
    port map (
            O => \N__40113\,
            I => \N__40104\
        );

    \I__8778\ : LocalMux
    port map (
            O => \N__40110\,
            I => \N__40101\
        );

    \I__8777\ : Span4Mux_v
    port map (
            O => \N__40107\,
            I => \N__40096\
        );

    \I__8776\ : LocalMux
    port map (
            O => \N__40104\,
            I => \N__40096\
        );

    \I__8775\ : Span4Mux_h
    port map (
            O => \N__40101\,
            I => \N__40090\
        );

    \I__8774\ : Span4Mux_h
    port map (
            O => \N__40096\,
            I => \N__40090\
        );

    \I__8773\ : InMux
    port map (
            O => \N__40095\,
            I => \N__40087\
        );

    \I__8772\ : Odrv4
    port map (
            O => \N__40090\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__8771\ : LocalMux
    port map (
            O => \N__40087\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__8770\ : CascadeMux
    port map (
            O => \N__40082\,
            I => \N__40079\
        );

    \I__8769\ : InMux
    port map (
            O => \N__40079\,
            I => \N__40076\
        );

    \I__8768\ : LocalMux
    port map (
            O => \N__40076\,
            I => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\
        );

    \I__8767\ : InMux
    port map (
            O => \N__40073\,
            I => \N__40069\
        );

    \I__8766\ : InMux
    port map (
            O => \N__40072\,
            I => \N__40066\
        );

    \I__8765\ : LocalMux
    port map (
            O => \N__40069\,
            I => \N__40062\
        );

    \I__8764\ : LocalMux
    port map (
            O => \N__40066\,
            I => \N__40059\
        );

    \I__8763\ : InMux
    port map (
            O => \N__40065\,
            I => \N__40056\
        );

    \I__8762\ : Span4Mux_h
    port map (
            O => \N__40062\,
            I => \N__40053\
        );

    \I__8761\ : Span4Mux_h
    port map (
            O => \N__40059\,
            I => \N__40049\
        );

    \I__8760\ : LocalMux
    port map (
            O => \N__40056\,
            I => \N__40046\
        );

    \I__8759\ : Span4Mux_v
    port map (
            O => \N__40053\,
            I => \N__40043\
        );

    \I__8758\ : InMux
    port map (
            O => \N__40052\,
            I => \N__40040\
        );

    \I__8757\ : Odrv4
    port map (
            O => \N__40049\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__8756\ : Odrv12
    port map (
            O => \N__40046\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__8755\ : Odrv4
    port map (
            O => \N__40043\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__8754\ : LocalMux
    port map (
            O => \N__40040\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__8753\ : CascadeMux
    port map (
            O => \N__40031\,
            I => \N__40028\
        );

    \I__8752\ : InMux
    port map (
            O => \N__40028\,
            I => \N__40025\
        );

    \I__8751\ : LocalMux
    port map (
            O => \N__40025\,
            I => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\
        );

    \I__8750\ : InMux
    port map (
            O => \N__40022\,
            I => \N__40019\
        );

    \I__8749\ : LocalMux
    port map (
            O => \N__40019\,
            I => \N__40014\
        );

    \I__8748\ : InMux
    port map (
            O => \N__40018\,
            I => \N__40011\
        );

    \I__8747\ : InMux
    port map (
            O => \N__40017\,
            I => \N__40008\
        );

    \I__8746\ : Span4Mux_v
    port map (
            O => \N__40014\,
            I => \N__40003\
        );

    \I__8745\ : LocalMux
    port map (
            O => \N__40011\,
            I => \N__40003\
        );

    \I__8744\ : LocalMux
    port map (
            O => \N__40008\,
            I => \N__40000\
        );

    \I__8743\ : Span4Mux_h
    port map (
            O => \N__40003\,
            I => \N__39994\
        );

    \I__8742\ : Span4Mux_h
    port map (
            O => \N__40000\,
            I => \N__39994\
        );

    \I__8741\ : InMux
    port map (
            O => \N__39999\,
            I => \N__39991\
        );

    \I__8740\ : Odrv4
    port map (
            O => \N__39994\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__8739\ : LocalMux
    port map (
            O => \N__39991\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__8738\ : CascadeMux
    port map (
            O => \N__39986\,
            I => \N__39983\
        );

    \I__8737\ : InMux
    port map (
            O => \N__39983\,
            I => \N__39980\
        );

    \I__8736\ : LocalMux
    port map (
            O => \N__39980\,
            I => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\
        );

    \I__8735\ : InMux
    port map (
            O => \N__39977\,
            I => \N__39974\
        );

    \I__8734\ : LocalMux
    port map (
            O => \N__39974\,
            I => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\
        );

    \I__8733\ : InMux
    port map (
            O => \N__39971\,
            I => \N__39966\
        );

    \I__8732\ : InMux
    port map (
            O => \N__39970\,
            I => \N__39963\
        );

    \I__8731\ : InMux
    port map (
            O => \N__39969\,
            I => \N__39960\
        );

    \I__8730\ : LocalMux
    port map (
            O => \N__39966\,
            I => \N__39957\
        );

    \I__8729\ : LocalMux
    port map (
            O => \N__39963\,
            I => \N__39952\
        );

    \I__8728\ : LocalMux
    port map (
            O => \N__39960\,
            I => \N__39952\
        );

    \I__8727\ : Span4Mux_h
    port map (
            O => \N__39957\,
            I => \N__39946\
        );

    \I__8726\ : Span4Mux_h
    port map (
            O => \N__39952\,
            I => \N__39946\
        );

    \I__8725\ : InMux
    port map (
            O => \N__39951\,
            I => \N__39943\
        );

    \I__8724\ : Odrv4
    port map (
            O => \N__39946\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__8723\ : LocalMux
    port map (
            O => \N__39943\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__8722\ : InMux
    port map (
            O => \N__39938\,
            I => \N__39935\
        );

    \I__8721\ : LocalMux
    port map (
            O => \N__39935\,
            I => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\
        );

    \I__8720\ : InMux
    port map (
            O => \N__39932\,
            I => \N__39929\
        );

    \I__8719\ : LocalMux
    port map (
            O => \N__39929\,
            I => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\
        );

    \I__8718\ : CascadeMux
    port map (
            O => \N__39926\,
            I => \N__39922\
        );

    \I__8717\ : CascadeMux
    port map (
            O => \N__39925\,
            I => \N__39919\
        );

    \I__8716\ : InMux
    port map (
            O => \N__39922\,
            I => \N__39915\
        );

    \I__8715\ : InMux
    port map (
            O => \N__39919\,
            I => \N__39912\
        );

    \I__8714\ : InMux
    port map (
            O => \N__39918\,
            I => \N__39909\
        );

    \I__8713\ : LocalMux
    port map (
            O => \N__39915\,
            I => \N__39904\
        );

    \I__8712\ : LocalMux
    port map (
            O => \N__39912\,
            I => \N__39904\
        );

    \I__8711\ : LocalMux
    port map (
            O => \N__39909\,
            I => \N__39901\
        );

    \I__8710\ : Span4Mux_h
    port map (
            O => \N__39904\,
            I => \N__39895\
        );

    \I__8709\ : Span4Mux_h
    port map (
            O => \N__39901\,
            I => \N__39895\
        );

    \I__8708\ : InMux
    port map (
            O => \N__39900\,
            I => \N__39892\
        );

    \I__8707\ : Odrv4
    port map (
            O => \N__39895\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__8706\ : LocalMux
    port map (
            O => \N__39892\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__8705\ : CascadeMux
    port map (
            O => \N__39887\,
            I => \N__39884\
        );

    \I__8704\ : InMux
    port map (
            O => \N__39884\,
            I => \N__39881\
        );

    \I__8703\ : LocalMux
    port map (
            O => \N__39881\,
            I => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\
        );

    \I__8702\ : InMux
    port map (
            O => \N__39878\,
            I => \N__39873\
        );

    \I__8701\ : InMux
    port map (
            O => \N__39877\,
            I => \N__39870\
        );

    \I__8700\ : InMux
    port map (
            O => \N__39876\,
            I => \N__39867\
        );

    \I__8699\ : LocalMux
    port map (
            O => \N__39873\,
            I => \N__39864\
        );

    \I__8698\ : LocalMux
    port map (
            O => \N__39870\,
            I => \N__39861\
        );

    \I__8697\ : LocalMux
    port map (
            O => \N__39867\,
            I => \N__39857\
        );

    \I__8696\ : Span4Mux_h
    port map (
            O => \N__39864\,
            I => \N__39852\
        );

    \I__8695\ : Span4Mux_h
    port map (
            O => \N__39861\,
            I => \N__39852\
        );

    \I__8694\ : InMux
    port map (
            O => \N__39860\,
            I => \N__39849\
        );

    \I__8693\ : Odrv12
    port map (
            O => \N__39857\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__8692\ : Odrv4
    port map (
            O => \N__39852\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__8691\ : LocalMux
    port map (
            O => \N__39849\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__8690\ : CascadeMux
    port map (
            O => \N__39842\,
            I => \N__39839\
        );

    \I__8689\ : InMux
    port map (
            O => \N__39839\,
            I => \N__39836\
        );

    \I__8688\ : LocalMux
    port map (
            O => \N__39836\,
            I => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\
        );

    \I__8687\ : CascadeMux
    port map (
            O => \N__39833\,
            I => \N__39830\
        );

    \I__8686\ : InMux
    port map (
            O => \N__39830\,
            I => \N__39827\
        );

    \I__8685\ : LocalMux
    port map (
            O => \N__39827\,
            I => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\
        );

    \I__8684\ : CascadeMux
    port map (
            O => \N__39824\,
            I => \N__39819\
        );

    \I__8683\ : CascadeMux
    port map (
            O => \N__39823\,
            I => \N__39816\
        );

    \I__8682\ : InMux
    port map (
            O => \N__39822\,
            I => \N__39813\
        );

    \I__8681\ : InMux
    port map (
            O => \N__39819\,
            I => \N__39808\
        );

    \I__8680\ : InMux
    port map (
            O => \N__39816\,
            I => \N__39808\
        );

    \I__8679\ : LocalMux
    port map (
            O => \N__39813\,
            I => \N__39805\
        );

    \I__8678\ : LocalMux
    port map (
            O => \N__39808\,
            I => \N__39801\
        );

    \I__8677\ : Span4Mux_h
    port map (
            O => \N__39805\,
            I => \N__39798\
        );

    \I__8676\ : InMux
    port map (
            O => \N__39804\,
            I => \N__39795\
        );

    \I__8675\ : Odrv12
    port map (
            O => \N__39801\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__8674\ : Odrv4
    port map (
            O => \N__39798\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__8673\ : LocalMux
    port map (
            O => \N__39795\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__8672\ : CascadeMux
    port map (
            O => \N__39788\,
            I => \N__39785\
        );

    \I__8671\ : InMux
    port map (
            O => \N__39785\,
            I => \N__39782\
        );

    \I__8670\ : LocalMux
    port map (
            O => \N__39782\,
            I => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\
        );

    \I__8669\ : CascadeMux
    port map (
            O => \N__39779\,
            I => \N__39776\
        );

    \I__8668\ : InMux
    port map (
            O => \N__39776\,
            I => \N__39773\
        );

    \I__8667\ : LocalMux
    port map (
            O => \N__39773\,
            I => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\
        );

    \I__8666\ : CascadeMux
    port map (
            O => \N__39770\,
            I => \N__39767\
        );

    \I__8665\ : InMux
    port map (
            O => \N__39767\,
            I => \N__39764\
        );

    \I__8664\ : LocalMux
    port map (
            O => \N__39764\,
            I => \N__39761\
        );

    \I__8663\ : Odrv12
    port map (
            O => \N__39761\,
            I => \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0\
        );

    \I__8662\ : CascadeMux
    port map (
            O => \N__39758\,
            I => \N__39754\
        );

    \I__8661\ : CascadeMux
    port map (
            O => \N__39757\,
            I => \N__39751\
        );

    \I__8660\ : InMux
    port map (
            O => \N__39754\,
            I => \N__39747\
        );

    \I__8659\ : InMux
    port map (
            O => \N__39751\,
            I => \N__39744\
        );

    \I__8658\ : InMux
    port map (
            O => \N__39750\,
            I => \N__39741\
        );

    \I__8657\ : LocalMux
    port map (
            O => \N__39747\,
            I => \N__39736\
        );

    \I__8656\ : LocalMux
    port map (
            O => \N__39744\,
            I => \N__39736\
        );

    \I__8655\ : LocalMux
    port map (
            O => \N__39741\,
            I => \N__39733\
        );

    \I__8654\ : Span4Mux_h
    port map (
            O => \N__39736\,
            I => \N__39728\
        );

    \I__8653\ : Span4Mux_h
    port map (
            O => \N__39733\,
            I => \N__39728\
        );

    \I__8652\ : Span4Mux_v
    port map (
            O => \N__39728\,
            I => \N__39724\
        );

    \I__8651\ : InMux
    port map (
            O => \N__39727\,
            I => \N__39721\
        );

    \I__8650\ : Odrv4
    port map (
            O => \N__39724\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__8649\ : LocalMux
    port map (
            O => \N__39721\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__8648\ : InMux
    port map (
            O => \N__39716\,
            I => \N__39713\
        );

    \I__8647\ : LocalMux
    port map (
            O => \N__39713\,
            I => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\
        );

    \I__8646\ : CascadeMux
    port map (
            O => \N__39710\,
            I => \N__39706\
        );

    \I__8645\ : CascadeMux
    port map (
            O => \N__39709\,
            I => \N__39703\
        );

    \I__8644\ : InMux
    port map (
            O => \N__39706\,
            I => \N__39697\
        );

    \I__8643\ : InMux
    port map (
            O => \N__39703\,
            I => \N__39697\
        );

    \I__8642\ : InMux
    port map (
            O => \N__39702\,
            I => \N__39694\
        );

    \I__8641\ : LocalMux
    port map (
            O => \N__39697\,
            I => \N__39691\
        );

    \I__8640\ : LocalMux
    port map (
            O => \N__39694\,
            I => \N__39688\
        );

    \I__8639\ : Span4Mux_h
    port map (
            O => \N__39691\,
            I => \N__39682\
        );

    \I__8638\ : Span4Mux_h
    port map (
            O => \N__39688\,
            I => \N__39682\
        );

    \I__8637\ : InMux
    port map (
            O => \N__39687\,
            I => \N__39679\
        );

    \I__8636\ : Odrv4
    port map (
            O => \N__39682\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__8635\ : LocalMux
    port map (
            O => \N__39679\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__8634\ : CascadeMux
    port map (
            O => \N__39674\,
            I => \N__39671\
        );

    \I__8633\ : InMux
    port map (
            O => \N__39671\,
            I => \N__39668\
        );

    \I__8632\ : LocalMux
    port map (
            O => \N__39668\,
            I => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\
        );

    \I__8631\ : CascadeMux
    port map (
            O => \N__39665\,
            I => \N__39661\
        );

    \I__8630\ : InMux
    port map (
            O => \N__39664\,
            I => \N__39657\
        );

    \I__8629\ : InMux
    port map (
            O => \N__39661\,
            I => \N__39654\
        );

    \I__8628\ : InMux
    port map (
            O => \N__39660\,
            I => \N__39651\
        );

    \I__8627\ : LocalMux
    port map (
            O => \N__39657\,
            I => \N__39648\
        );

    \I__8626\ : LocalMux
    port map (
            O => \N__39654\,
            I => \N__39643\
        );

    \I__8625\ : LocalMux
    port map (
            O => \N__39651\,
            I => \N__39643\
        );

    \I__8624\ : Span4Mux_h
    port map (
            O => \N__39648\,
            I => \N__39637\
        );

    \I__8623\ : Span4Mux_h
    port map (
            O => \N__39643\,
            I => \N__39637\
        );

    \I__8622\ : InMux
    port map (
            O => \N__39642\,
            I => \N__39634\
        );

    \I__8621\ : Odrv4
    port map (
            O => \N__39637\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__8620\ : LocalMux
    port map (
            O => \N__39634\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__8619\ : CascadeMux
    port map (
            O => \N__39629\,
            I => \N__39626\
        );

    \I__8618\ : InMux
    port map (
            O => \N__39626\,
            I => \N__39623\
        );

    \I__8617\ : LocalMux
    port map (
            O => \N__39623\,
            I => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\
        );

    \I__8616\ : CascadeMux
    port map (
            O => \N__39620\,
            I => \N__39616\
        );

    \I__8615\ : CascadeMux
    port map (
            O => \N__39619\,
            I => \N__39612\
        );

    \I__8614\ : InMux
    port map (
            O => \N__39616\,
            I => \N__39609\
        );

    \I__8613\ : InMux
    port map (
            O => \N__39615\,
            I => \N__39606\
        );

    \I__8612\ : InMux
    port map (
            O => \N__39612\,
            I => \N__39603\
        );

    \I__8611\ : LocalMux
    port map (
            O => \N__39609\,
            I => \N__39600\
        );

    \I__8610\ : LocalMux
    port map (
            O => \N__39606\,
            I => \N__39597\
        );

    \I__8609\ : LocalMux
    port map (
            O => \N__39603\,
            I => \N__39593\
        );

    \I__8608\ : Span4Mux_h
    port map (
            O => \N__39600\,
            I => \N__39588\
        );

    \I__8607\ : Span4Mux_h
    port map (
            O => \N__39597\,
            I => \N__39588\
        );

    \I__8606\ : InMux
    port map (
            O => \N__39596\,
            I => \N__39585\
        );

    \I__8605\ : Odrv12
    port map (
            O => \N__39593\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__8604\ : Odrv4
    port map (
            O => \N__39588\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__8603\ : LocalMux
    port map (
            O => \N__39585\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__8602\ : InMux
    port map (
            O => \N__39578\,
            I => \N__39575\
        );

    \I__8601\ : LocalMux
    port map (
            O => \N__39575\,
            I => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\
        );

    \I__8600\ : InMux
    port map (
            O => \N__39572\,
            I => \N__39568\
        );

    \I__8599\ : InMux
    port map (
            O => \N__39571\,
            I => \N__39564\
        );

    \I__8598\ : LocalMux
    port map (
            O => \N__39568\,
            I => \N__39561\
        );

    \I__8597\ : InMux
    port map (
            O => \N__39567\,
            I => \N__39558\
        );

    \I__8596\ : LocalMux
    port map (
            O => \N__39564\,
            I => \N__39553\
        );

    \I__8595\ : Span4Mux_h
    port map (
            O => \N__39561\,
            I => \N__39553\
        );

    \I__8594\ : LocalMux
    port map (
            O => \N__39558\,
            I => \N__39549\
        );

    \I__8593\ : Span4Mux_h
    port map (
            O => \N__39553\,
            I => \N__39546\
        );

    \I__8592\ : InMux
    port map (
            O => \N__39552\,
            I => \N__39543\
        );

    \I__8591\ : Odrv12
    port map (
            O => \N__39549\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__8590\ : Odrv4
    port map (
            O => \N__39546\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__8589\ : LocalMux
    port map (
            O => \N__39543\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__8588\ : InMux
    port map (
            O => \N__39536\,
            I => \N__39533\
        );

    \I__8587\ : LocalMux
    port map (
            O => \N__39533\,
            I => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\
        );

    \I__8586\ : InMux
    port map (
            O => \N__39530\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\
        );

    \I__8585\ : CascadeMux
    port map (
            O => \N__39527\,
            I => \N__39522\
        );

    \I__8584\ : InMux
    port map (
            O => \N__39526\,
            I => \N__39517\
        );

    \I__8583\ : InMux
    port map (
            O => \N__39525\,
            I => \N__39517\
        );

    \I__8582\ : InMux
    port map (
            O => \N__39522\,
            I => \N__39513\
        );

    \I__8581\ : LocalMux
    port map (
            O => \N__39517\,
            I => \N__39510\
        );

    \I__8580\ : InMux
    port map (
            O => \N__39516\,
            I => \N__39507\
        );

    \I__8579\ : LocalMux
    port map (
            O => \N__39513\,
            I => \N__39504\
        );

    \I__8578\ : Span4Mux_h
    port map (
            O => \N__39510\,
            I => \N__39501\
        );

    \I__8577\ : LocalMux
    port map (
            O => \N__39507\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__8576\ : Odrv12
    port map (
            O => \N__39504\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__8575\ : Odrv4
    port map (
            O => \N__39501\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__8574\ : InMux
    port map (
            O => \N__39494\,
            I => \N__39490\
        );

    \I__8573\ : InMux
    port map (
            O => \N__39493\,
            I => \N__39486\
        );

    \I__8572\ : LocalMux
    port map (
            O => \N__39490\,
            I => \N__39483\
        );

    \I__8571\ : InMux
    port map (
            O => \N__39489\,
            I => \N__39480\
        );

    \I__8570\ : LocalMux
    port map (
            O => \N__39486\,
            I => \N__39475\
        );

    \I__8569\ : Span4Mux_h
    port map (
            O => \N__39483\,
            I => \N__39475\
        );

    \I__8568\ : LocalMux
    port map (
            O => \N__39480\,
            I => \N__39471\
        );

    \I__8567\ : Span4Mux_v
    port map (
            O => \N__39475\,
            I => \N__39468\
        );

    \I__8566\ : InMux
    port map (
            O => \N__39474\,
            I => \N__39465\
        );

    \I__8565\ : Odrv12
    port map (
            O => \N__39471\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__8564\ : Odrv4
    port map (
            O => \N__39468\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__8563\ : LocalMux
    port map (
            O => \N__39465\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__8562\ : InMux
    port map (
            O => \N__39458\,
            I => \N__39455\
        );

    \I__8561\ : LocalMux
    port map (
            O => \N__39455\,
            I => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\
        );

    \I__8560\ : InMux
    port map (
            O => \N__39452\,
            I => \N__39449\
        );

    \I__8559\ : LocalMux
    port map (
            O => \N__39449\,
            I => \N__39444\
        );

    \I__8558\ : InMux
    port map (
            O => \N__39448\,
            I => \N__39441\
        );

    \I__8557\ : InMux
    port map (
            O => \N__39447\,
            I => \N__39438\
        );

    \I__8556\ : Span4Mux_h
    port map (
            O => \N__39444\,
            I => \N__39435\
        );

    \I__8555\ : LocalMux
    port map (
            O => \N__39441\,
            I => \N__39429\
        );

    \I__8554\ : LocalMux
    port map (
            O => \N__39438\,
            I => \N__39429\
        );

    \I__8553\ : Span4Mux_v
    port map (
            O => \N__39435\,
            I => \N__39426\
        );

    \I__8552\ : InMux
    port map (
            O => \N__39434\,
            I => \N__39423\
        );

    \I__8551\ : Odrv12
    port map (
            O => \N__39429\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__8550\ : Odrv4
    port map (
            O => \N__39426\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__8549\ : LocalMux
    port map (
            O => \N__39423\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__8548\ : CascadeMux
    port map (
            O => \N__39416\,
            I => \N__39413\
        );

    \I__8547\ : InMux
    port map (
            O => \N__39413\,
            I => \N__39410\
        );

    \I__8546\ : LocalMux
    port map (
            O => \N__39410\,
            I => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\
        );

    \I__8545\ : InMux
    port map (
            O => \N__39407\,
            I => \N__39400\
        );

    \I__8544\ : InMux
    port map (
            O => \N__39406\,
            I => \N__39400\
        );

    \I__8543\ : InMux
    port map (
            O => \N__39405\,
            I => \N__39397\
        );

    \I__8542\ : LocalMux
    port map (
            O => \N__39400\,
            I => \N__39392\
        );

    \I__8541\ : LocalMux
    port map (
            O => \N__39397\,
            I => \N__39392\
        );

    \I__8540\ : Span4Mux_h
    port map (
            O => \N__39392\,
            I => \N__39388\
        );

    \I__8539\ : InMux
    port map (
            O => \N__39391\,
            I => \N__39385\
        );

    \I__8538\ : Odrv4
    port map (
            O => \N__39388\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__8537\ : LocalMux
    port map (
            O => \N__39385\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__8536\ : InMux
    port map (
            O => \N__39380\,
            I => \N__39377\
        );

    \I__8535\ : LocalMux
    port map (
            O => \N__39377\,
            I => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\
        );

    \I__8534\ : CascadeMux
    port map (
            O => \N__39374\,
            I => \N__39370\
        );

    \I__8533\ : CascadeMux
    port map (
            O => \N__39373\,
            I => \N__39366\
        );

    \I__8532\ : InMux
    port map (
            O => \N__39370\,
            I => \N__39363\
        );

    \I__8531\ : InMux
    port map (
            O => \N__39369\,
            I => \N__39360\
        );

    \I__8530\ : InMux
    port map (
            O => \N__39366\,
            I => \N__39357\
        );

    \I__8529\ : LocalMux
    port map (
            O => \N__39363\,
            I => \N__39354\
        );

    \I__8528\ : LocalMux
    port map (
            O => \N__39360\,
            I => \N__39351\
        );

    \I__8527\ : LocalMux
    port map (
            O => \N__39357\,
            I => \N__39343\
        );

    \I__8526\ : Span4Mux_h
    port map (
            O => \N__39354\,
            I => \N__39343\
        );

    \I__8525\ : Span4Mux_h
    port map (
            O => \N__39351\,
            I => \N__39343\
        );

    \I__8524\ : InMux
    port map (
            O => \N__39350\,
            I => \N__39340\
        );

    \I__8523\ : Odrv4
    port map (
            O => \N__39343\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__8522\ : LocalMux
    port map (
            O => \N__39340\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__8521\ : CascadeMux
    port map (
            O => \N__39335\,
            I => \N__39332\
        );

    \I__8520\ : InMux
    port map (
            O => \N__39332\,
            I => \N__39329\
        );

    \I__8519\ : LocalMux
    port map (
            O => \N__39329\,
            I => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\
        );

    \I__8518\ : CascadeMux
    port map (
            O => \N__39326\,
            I => \N__39322\
        );

    \I__8517\ : InMux
    port map (
            O => \N__39325\,
            I => \N__39316\
        );

    \I__8516\ : InMux
    port map (
            O => \N__39322\,
            I => \N__39316\
        );

    \I__8515\ : InMux
    port map (
            O => \N__39321\,
            I => \N__39313\
        );

    \I__8514\ : LocalMux
    port map (
            O => \N__39316\,
            I => \N__39310\
        );

    \I__8513\ : LocalMux
    port map (
            O => \N__39313\,
            I => \N__39307\
        );

    \I__8512\ : Span4Mux_h
    port map (
            O => \N__39310\,
            I => \N__39301\
        );

    \I__8511\ : Span4Mux_h
    port map (
            O => \N__39307\,
            I => \N__39301\
        );

    \I__8510\ : InMux
    port map (
            O => \N__39306\,
            I => \N__39298\
        );

    \I__8509\ : Odrv4
    port map (
            O => \N__39301\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__8508\ : LocalMux
    port map (
            O => \N__39298\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__8507\ : InMux
    port map (
            O => \N__39293\,
            I => \N__39290\
        );

    \I__8506\ : LocalMux
    port map (
            O => \N__39290\,
            I => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\
        );

    \I__8505\ : InMux
    port map (
            O => \N__39287\,
            I => \N__39284\
        );

    \I__8504\ : LocalMux
    port map (
            O => \N__39284\,
            I => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\
        );

    \I__8503\ : InMux
    port map (
            O => \N__39281\,
            I => \N__39277\
        );

    \I__8502\ : InMux
    port map (
            O => \N__39280\,
            I => \N__39274\
        );

    \I__8501\ : LocalMux
    port map (
            O => \N__39277\,
            I => \N__39270\
        );

    \I__8500\ : LocalMux
    port map (
            O => \N__39274\,
            I => \N__39267\
        );

    \I__8499\ : InMux
    port map (
            O => \N__39273\,
            I => \N__39263\
        );

    \I__8498\ : Span4Mux_h
    port map (
            O => \N__39270\,
            I => \N__39258\
        );

    \I__8497\ : Span4Mux_h
    port map (
            O => \N__39267\,
            I => \N__39258\
        );

    \I__8496\ : InMux
    port map (
            O => \N__39266\,
            I => \N__39255\
        );

    \I__8495\ : LocalMux
    port map (
            O => \N__39263\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__8494\ : Odrv4
    port map (
            O => \N__39258\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__8493\ : LocalMux
    port map (
            O => \N__39255\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__8492\ : CascadeMux
    port map (
            O => \N__39248\,
            I => \N__39245\
        );

    \I__8491\ : InMux
    port map (
            O => \N__39245\,
            I => \N__39242\
        );

    \I__8490\ : LocalMux
    port map (
            O => \N__39242\,
            I => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\
        );

    \I__8489\ : CascadeMux
    port map (
            O => \N__39239\,
            I => \N__39236\
        );

    \I__8488\ : InMux
    port map (
            O => \N__39236\,
            I => \N__39231\
        );

    \I__8487\ : InMux
    port map (
            O => \N__39235\,
            I => \N__39228\
        );

    \I__8486\ : InMux
    port map (
            O => \N__39234\,
            I => \N__39225\
        );

    \I__8485\ : LocalMux
    port map (
            O => \N__39231\,
            I => \N__39220\
        );

    \I__8484\ : LocalMux
    port map (
            O => \N__39228\,
            I => \N__39220\
        );

    \I__8483\ : LocalMux
    port map (
            O => \N__39225\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__8482\ : Odrv12
    port map (
            O => \N__39220\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__8481\ : InMux
    port map (
            O => \N__39215\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\
        );

    \I__8480\ : CascadeMux
    port map (
            O => \N__39212\,
            I => \N__39209\
        );

    \I__8479\ : InMux
    port map (
            O => \N__39209\,
            I => \N__39202\
        );

    \I__8478\ : InMux
    port map (
            O => \N__39208\,
            I => \N__39202\
        );

    \I__8477\ : InMux
    port map (
            O => \N__39207\,
            I => \N__39199\
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__39202\,
            I => \N__39196\
        );

    \I__8475\ : LocalMux
    port map (
            O => \N__39199\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__8474\ : Odrv12
    port map (
            O => \N__39196\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__8473\ : InMux
    port map (
            O => \N__39191\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\
        );

    \I__8472\ : InMux
    port map (
            O => \N__39188\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\
        );

    \I__8471\ : InMux
    port map (
            O => \N__39185\,
            I => \bfn_17_13_0_\
        );

    \I__8470\ : InMux
    port map (
            O => \N__39182\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\
        );

    \I__8469\ : InMux
    port map (
            O => \N__39179\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\
        );

    \I__8468\ : InMux
    port map (
            O => \N__39176\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\
        );

    \I__8467\ : InMux
    port map (
            O => \N__39173\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\
        );

    \I__8466\ : CascadeMux
    port map (
            O => \N__39170\,
            I => \N__39166\
        );

    \I__8465\ : InMux
    port map (
            O => \N__39169\,
            I => \N__39160\
        );

    \I__8464\ : InMux
    port map (
            O => \N__39166\,
            I => \N__39160\
        );

    \I__8463\ : InMux
    port map (
            O => \N__39165\,
            I => \N__39156\
        );

    \I__8462\ : LocalMux
    port map (
            O => \N__39160\,
            I => \N__39153\
        );

    \I__8461\ : InMux
    port map (
            O => \N__39159\,
            I => \N__39150\
        );

    \I__8460\ : LocalMux
    port map (
            O => \N__39156\,
            I => \N__39147\
        );

    \I__8459\ : Span4Mux_h
    port map (
            O => \N__39153\,
            I => \N__39144\
        );

    \I__8458\ : LocalMux
    port map (
            O => \N__39150\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__8457\ : Odrv12
    port map (
            O => \N__39147\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__8456\ : Odrv4
    port map (
            O => \N__39144\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__8455\ : InMux
    port map (
            O => \N__39137\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\
        );

    \I__8454\ : InMux
    port map (
            O => \N__39134\,
            I => \N__39130\
        );

    \I__8453\ : InMux
    port map (
            O => \N__39133\,
            I => \N__39127\
        );

    \I__8452\ : LocalMux
    port map (
            O => \N__39130\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__8451\ : LocalMux
    port map (
            O => \N__39127\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__8450\ : InMux
    port map (
            O => \N__39122\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\
        );

    \I__8449\ : InMux
    port map (
            O => \N__39119\,
            I => \N__39115\
        );

    \I__8448\ : InMux
    port map (
            O => \N__39118\,
            I => \N__39112\
        );

    \I__8447\ : LocalMux
    port map (
            O => \N__39115\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__8446\ : LocalMux
    port map (
            O => \N__39112\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__8445\ : InMux
    port map (
            O => \N__39107\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\
        );

    \I__8444\ : InMux
    port map (
            O => \N__39104\,
            I => \N__39100\
        );

    \I__8443\ : InMux
    port map (
            O => \N__39103\,
            I => \N__39097\
        );

    \I__8442\ : LocalMux
    port map (
            O => \N__39100\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__8441\ : LocalMux
    port map (
            O => \N__39097\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__8440\ : InMux
    port map (
            O => \N__39092\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\
        );

    \I__8439\ : InMux
    port map (
            O => \N__39089\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\
        );

    \I__8438\ : InMux
    port map (
            O => \N__39086\,
            I => \bfn_17_12_0_\
        );

    \I__8437\ : InMux
    port map (
            O => \N__39083\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\
        );

    \I__8436\ : InMux
    port map (
            O => \N__39080\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\
        );

    \I__8435\ : CascadeMux
    port map (
            O => \N__39077\,
            I => \N__39073\
        );

    \I__8434\ : InMux
    port map (
            O => \N__39076\,
            I => \N__39067\
        );

    \I__8433\ : InMux
    port map (
            O => \N__39073\,
            I => \N__39067\
        );

    \I__8432\ : InMux
    port map (
            O => \N__39072\,
            I => \N__39064\
        );

    \I__8431\ : LocalMux
    port map (
            O => \N__39067\,
            I => \N__39061\
        );

    \I__8430\ : LocalMux
    port map (
            O => \N__39064\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__8429\ : Odrv4
    port map (
            O => \N__39061\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__8428\ : InMux
    port map (
            O => \N__39056\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\
        );

    \I__8427\ : InMux
    port map (
            O => \N__39053\,
            I => \N__39046\
        );

    \I__8426\ : InMux
    port map (
            O => \N__39052\,
            I => \N__39046\
        );

    \I__8425\ : InMux
    port map (
            O => \N__39051\,
            I => \N__39043\
        );

    \I__8424\ : LocalMux
    port map (
            O => \N__39046\,
            I => \N__39040\
        );

    \I__8423\ : LocalMux
    port map (
            O => \N__39043\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__8422\ : Odrv4
    port map (
            O => \N__39040\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__8421\ : InMux
    port map (
            O => \N__39035\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__8420\ : InMux
    port map (
            O => \N__39032\,
            I => \N__39028\
        );

    \I__8419\ : InMux
    port map (
            O => \N__39031\,
            I => \N__39025\
        );

    \I__8418\ : LocalMux
    port map (
            O => \N__39028\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__8417\ : LocalMux
    port map (
            O => \N__39025\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__8416\ : InMux
    port map (
            O => \N__39020\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\
        );

    \I__8415\ : InMux
    port map (
            O => \N__39017\,
            I => \N__39013\
        );

    \I__8414\ : InMux
    port map (
            O => \N__39016\,
            I => \N__39010\
        );

    \I__8413\ : LocalMux
    port map (
            O => \N__39013\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__8412\ : LocalMux
    port map (
            O => \N__39010\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__8411\ : InMux
    port map (
            O => \N__39005\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\
        );

    \I__8410\ : InMux
    port map (
            O => \N__39002\,
            I => \N__38998\
        );

    \I__8409\ : InMux
    port map (
            O => \N__39001\,
            I => \N__38995\
        );

    \I__8408\ : LocalMux
    port map (
            O => \N__38998\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__8407\ : LocalMux
    port map (
            O => \N__38995\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__8406\ : InMux
    port map (
            O => \N__38990\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\
        );

    \I__8405\ : InMux
    port map (
            O => \N__38987\,
            I => \N__38983\
        );

    \I__8404\ : InMux
    port map (
            O => \N__38986\,
            I => \N__38980\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__38983\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__8402\ : LocalMux
    port map (
            O => \N__38980\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__8401\ : InMux
    port map (
            O => \N__38975\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\
        );

    \I__8400\ : InMux
    port map (
            O => \N__38972\,
            I => \N__38968\
        );

    \I__8399\ : InMux
    port map (
            O => \N__38971\,
            I => \N__38965\
        );

    \I__8398\ : LocalMux
    port map (
            O => \N__38968\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__8397\ : LocalMux
    port map (
            O => \N__38965\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__8396\ : InMux
    port map (
            O => \N__38960\,
            I => \bfn_17_11_0_\
        );

    \I__8395\ : InMux
    port map (
            O => \N__38957\,
            I => \N__38953\
        );

    \I__8394\ : InMux
    port map (
            O => \N__38956\,
            I => \N__38950\
        );

    \I__8393\ : LocalMux
    port map (
            O => \N__38953\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__8392\ : LocalMux
    port map (
            O => \N__38950\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__8391\ : InMux
    port map (
            O => \N__38945\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\
        );

    \I__8390\ : InMux
    port map (
            O => \N__38942\,
            I => \N__38938\
        );

    \I__8389\ : InMux
    port map (
            O => \N__38941\,
            I => \N__38935\
        );

    \I__8388\ : LocalMux
    port map (
            O => \N__38938\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__8387\ : LocalMux
    port map (
            O => \N__38935\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__8386\ : InMux
    port map (
            O => \N__38930\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\
        );

    \I__8385\ : InMux
    port map (
            O => \N__38927\,
            I => \N__38923\
        );

    \I__8384\ : InMux
    port map (
            O => \N__38926\,
            I => \N__38920\
        );

    \I__8383\ : LocalMux
    port map (
            O => \N__38923\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__8382\ : LocalMux
    port map (
            O => \N__38920\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__8381\ : InMux
    port map (
            O => \N__38915\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\
        );

    \I__8380\ : InMux
    port map (
            O => \N__38912\,
            I => \N__38907\
        );

    \I__8379\ : InMux
    port map (
            O => \N__38911\,
            I => \N__38904\
        );

    \I__8378\ : InMux
    port map (
            O => \N__38910\,
            I => \N__38900\
        );

    \I__8377\ : LocalMux
    port map (
            O => \N__38907\,
            I => \N__38897\
        );

    \I__8376\ : LocalMux
    port map (
            O => \N__38904\,
            I => \N__38894\
        );

    \I__8375\ : InMux
    port map (
            O => \N__38903\,
            I => \N__38891\
        );

    \I__8374\ : LocalMux
    port map (
            O => \N__38900\,
            I => \N__38888\
        );

    \I__8373\ : Span4Mux_h
    port map (
            O => \N__38897\,
            I => \N__38885\
        );

    \I__8372\ : Span4Mux_v
    port map (
            O => \N__38894\,
            I => \N__38880\
        );

    \I__8371\ : LocalMux
    port map (
            O => \N__38891\,
            I => \N__38880\
        );

    \I__8370\ : Span4Mux_h
    port map (
            O => \N__38888\,
            I => \N__38877\
        );

    \I__8369\ : Span4Mux_v
    port map (
            O => \N__38885\,
            I => \N__38874\
        );

    \I__8368\ : Odrv4
    port map (
            O => \N__38880\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__8367\ : Odrv4
    port map (
            O => \N__38877\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__8366\ : Odrv4
    port map (
            O => \N__38874\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__8365\ : InMux
    port map (
            O => \N__38867\,
            I => \N__38862\
        );

    \I__8364\ : InMux
    port map (
            O => \N__38866\,
            I => \N__38859\
        );

    \I__8363\ : InMux
    port map (
            O => \N__38865\,
            I => \N__38856\
        );

    \I__8362\ : LocalMux
    port map (
            O => \N__38862\,
            I => \N__38851\
        );

    \I__8361\ : LocalMux
    port map (
            O => \N__38859\,
            I => \N__38851\
        );

    \I__8360\ : LocalMux
    port map (
            O => \N__38856\,
            I => \elapsed_time_ns_1_RNIU8PBB_0_20\
        );

    \I__8359\ : Odrv4
    port map (
            O => \N__38851\,
            I => \elapsed_time_ns_1_RNIU8PBB_0_20\
        );

    \I__8358\ : InMux
    port map (
            O => \N__38846\,
            I => \N__38843\
        );

    \I__8357\ : LocalMux
    port map (
            O => \N__38843\,
            I => \N__38838\
        );

    \I__8356\ : InMux
    port map (
            O => \N__38842\,
            I => \N__38833\
        );

    \I__8355\ : InMux
    port map (
            O => \N__38841\,
            I => \N__38833\
        );

    \I__8354\ : Span4Mux_h
    port map (
            O => \N__38838\,
            I => \N__38830\
        );

    \I__8353\ : LocalMux
    port map (
            O => \N__38833\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\
        );

    \I__8352\ : Odrv4
    port map (
            O => \N__38830\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\
        );

    \I__8351\ : InMux
    port map (
            O => \N__38825\,
            I => \N__38821\
        );

    \I__8350\ : CascadeMux
    port map (
            O => \N__38824\,
            I => \N__38818\
        );

    \I__8349\ : LocalMux
    port map (
            O => \N__38821\,
            I => \N__38814\
        );

    \I__8348\ : InMux
    port map (
            O => \N__38818\,
            I => \N__38809\
        );

    \I__8347\ : InMux
    port map (
            O => \N__38817\,
            I => \N__38809\
        );

    \I__8346\ : Span4Mux_v
    port map (
            O => \N__38814\,
            I => \N__38806\
        );

    \I__8345\ : LocalMux
    port map (
            O => \N__38809\,
            I => \N__38801\
        );

    \I__8344\ : Span4Mux_h
    port map (
            O => \N__38806\,
            I => \N__38801\
        );

    \I__8343\ : Odrv4
    port map (
            O => \N__38801\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\
        );

    \I__8342\ : InMux
    port map (
            O => \N__38798\,
            I => \N__38792\
        );

    \I__8341\ : InMux
    port map (
            O => \N__38797\,
            I => \N__38789\
        );

    \I__8340\ : InMux
    port map (
            O => \N__38796\,
            I => \N__38786\
        );

    \I__8339\ : InMux
    port map (
            O => \N__38795\,
            I => \N__38783\
        );

    \I__8338\ : LocalMux
    port map (
            O => \N__38792\,
            I => \N__38780\
        );

    \I__8337\ : LocalMux
    port map (
            O => \N__38789\,
            I => \N__38773\
        );

    \I__8336\ : LocalMux
    port map (
            O => \N__38786\,
            I => \N__38773\
        );

    \I__8335\ : LocalMux
    port map (
            O => \N__38783\,
            I => \N__38773\
        );

    \I__8334\ : Span4Mux_v
    port map (
            O => \N__38780\,
            I => \N__38770\
        );

    \I__8333\ : Span4Mux_v
    port map (
            O => \N__38773\,
            I => \N__38767\
        );

    \I__8332\ : Odrv4
    port map (
            O => \N__38770\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__8331\ : Odrv4
    port map (
            O => \N__38767\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__8330\ : InMux
    port map (
            O => \N__38762\,
            I => \N__38759\
        );

    \I__8329\ : LocalMux
    port map (
            O => \N__38759\,
            I => \N__38755\
        );

    \I__8328\ : InMux
    port map (
            O => \N__38758\,
            I => \N__38751\
        );

    \I__8327\ : Span4Mux_v
    port map (
            O => \N__38755\,
            I => \N__38748\
        );

    \I__8326\ : InMux
    port map (
            O => \N__38754\,
            I => \N__38745\
        );

    \I__8325\ : LocalMux
    port map (
            O => \N__38751\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7\
        );

    \I__8324\ : Odrv4
    port map (
            O => \N__38748\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7\
        );

    \I__8323\ : LocalMux
    port map (
            O => \N__38745\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7\
        );

    \I__8322\ : InMux
    port map (
            O => \N__38738\,
            I => \N__38732\
        );

    \I__8321\ : InMux
    port map (
            O => \N__38737\,
            I => \N__38729\
        );

    \I__8320\ : CascadeMux
    port map (
            O => \N__38736\,
            I => \N__38726\
        );

    \I__8319\ : InMux
    port map (
            O => \N__38735\,
            I => \N__38723\
        );

    \I__8318\ : LocalMux
    port map (
            O => \N__38732\,
            I => \N__38718\
        );

    \I__8317\ : LocalMux
    port map (
            O => \N__38729\,
            I => \N__38718\
        );

    \I__8316\ : InMux
    port map (
            O => \N__38726\,
            I => \N__38715\
        );

    \I__8315\ : LocalMux
    port map (
            O => \N__38723\,
            I => \N__38712\
        );

    \I__8314\ : Span4Mux_h
    port map (
            O => \N__38718\,
            I => \N__38709\
        );

    \I__8313\ : LocalMux
    port map (
            O => \N__38715\,
            I => \N__38706\
        );

    \I__8312\ : Odrv4
    port map (
            O => \N__38712\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__8311\ : Odrv4
    port map (
            O => \N__38709\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__8310\ : Odrv4
    port map (
            O => \N__38706\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__8309\ : InMux
    port map (
            O => \N__38699\,
            I => \N__38694\
        );

    \I__8308\ : InMux
    port map (
            O => \N__38698\,
            I => \N__38691\
        );

    \I__8307\ : InMux
    port map (
            O => \N__38697\,
            I => \N__38688\
        );

    \I__8306\ : LocalMux
    port map (
            O => \N__38694\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12\
        );

    \I__8305\ : LocalMux
    port map (
            O => \N__38691\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12\
        );

    \I__8304\ : LocalMux
    port map (
            O => \N__38688\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12\
        );

    \I__8303\ : CascadeMux
    port map (
            O => \N__38681\,
            I => \N__38678\
        );

    \I__8302\ : InMux
    port map (
            O => \N__38678\,
            I => \N__38675\
        );

    \I__8301\ : LocalMux
    port map (
            O => \N__38675\,
            I => \N__38671\
        );

    \I__8300\ : CascadeMux
    port map (
            O => \N__38674\,
            I => \N__38667\
        );

    \I__8299\ : Span4Mux_v
    port map (
            O => \N__38671\,
            I => \N__38664\
        );

    \I__8298\ : InMux
    port map (
            O => \N__38670\,
            I => \N__38661\
        );

    \I__8297\ : InMux
    port map (
            O => \N__38667\,
            I => \N__38658\
        );

    \I__8296\ : Sp12to4
    port map (
            O => \N__38664\,
            I => \N__38653\
        );

    \I__8295\ : LocalMux
    port map (
            O => \N__38661\,
            I => \N__38653\
        );

    \I__8294\ : LocalMux
    port map (
            O => \N__38658\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__8293\ : Odrv12
    port map (
            O => \N__38653\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__8292\ : InMux
    port map (
            O => \N__38648\,
            I => \N__38644\
        );

    \I__8291\ : InMux
    port map (
            O => \N__38647\,
            I => \N__38641\
        );

    \I__8290\ : LocalMux
    port map (
            O => \N__38644\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__8289\ : LocalMux
    port map (
            O => \N__38641\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__8288\ : InMux
    port map (
            O => \N__38636\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\
        );

    \I__8287\ : InMux
    port map (
            O => \N__38633\,
            I => \N__38629\
        );

    \I__8286\ : InMux
    port map (
            O => \N__38632\,
            I => \N__38626\
        );

    \I__8285\ : LocalMux
    port map (
            O => \N__38629\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__8284\ : LocalMux
    port map (
            O => \N__38626\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__8283\ : InMux
    port map (
            O => \N__38621\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\
        );

    \I__8282\ : InMux
    port map (
            O => \N__38618\,
            I => \N__38614\
        );

    \I__8281\ : InMux
    port map (
            O => \N__38617\,
            I => \N__38611\
        );

    \I__8280\ : LocalMux
    port map (
            O => \N__38614\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__38611\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__8278\ : InMux
    port map (
            O => \N__38606\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\
        );

    \I__8277\ : InMux
    port map (
            O => \N__38603\,
            I => \N__38600\
        );

    \I__8276\ : LocalMux
    port map (
            O => \N__38600\,
            I => \N__38597\
        );

    \I__8275\ : Odrv4
    port map (
            O => \N__38597\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17\
        );

    \I__8274\ : InMux
    port map (
            O => \N__38594\,
            I => \N__38591\
        );

    \I__8273\ : LocalMux
    port map (
            O => \N__38591\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23\
        );

    \I__8272\ : InMux
    port map (
            O => \N__38588\,
            I => \N__38585\
        );

    \I__8271\ : LocalMux
    port map (
            O => \N__38585\,
            I => \N__38582\
        );

    \I__8270\ : Span4Mux_h
    port map (
            O => \N__38582\,
            I => \N__38579\
        );

    \I__8269\ : Span4Mux_v
    port map (
            O => \N__38579\,
            I => \N__38576\
        );

    \I__8268\ : Odrv4
    port map (
            O => \N__38576\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt22\
        );

    \I__8267\ : CascadeMux
    port map (
            O => \N__38573\,
            I => \N__38570\
        );

    \I__8266\ : InMux
    port map (
            O => \N__38570\,
            I => \N__38567\
        );

    \I__8265\ : LocalMux
    port map (
            O => \N__38567\,
            I => \N__38564\
        );

    \I__8264\ : Span4Mux_v
    port map (
            O => \N__38564\,
            I => \N__38561\
        );

    \I__8263\ : Odrv4
    port map (
            O => \N__38561\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22\
        );

    \I__8262\ : InMux
    port map (
            O => \N__38558\,
            I => \N__38554\
        );

    \I__8261\ : InMux
    port map (
            O => \N__38557\,
            I => \N__38551\
        );

    \I__8260\ : LocalMux
    port map (
            O => \N__38554\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22\
        );

    \I__8259\ : LocalMux
    port map (
            O => \N__38551\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22\
        );

    \I__8258\ : CascadeMux
    port map (
            O => \N__38546\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22_cascade_\
        );

    \I__8257\ : InMux
    port map (
            O => \N__38543\,
            I => \N__38537\
        );

    \I__8256\ : InMux
    port map (
            O => \N__38542\,
            I => \N__38537\
        );

    \I__8255\ : LocalMux
    port map (
            O => \N__38537\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_22\
        );

    \I__8254\ : InMux
    port map (
            O => \N__38534\,
            I => \N__38531\
        );

    \I__8253\ : LocalMux
    port map (
            O => \N__38531\,
            I => \N__38528\
        );

    \I__8252\ : Span4Mux_h
    port map (
            O => \N__38528\,
            I => \N__38525\
        );

    \I__8251\ : Odrv4
    port map (
            O => \N__38525\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\
        );

    \I__8250\ : CascadeMux
    port map (
            O => \N__38522\,
            I => \N__38517\
        );

    \I__8249\ : InMux
    port map (
            O => \N__38521\,
            I => \N__38514\
        );

    \I__8248\ : InMux
    port map (
            O => \N__38520\,
            I => \N__38511\
        );

    \I__8247\ : InMux
    port map (
            O => \N__38517\,
            I => \N__38508\
        );

    \I__8246\ : LocalMux
    port map (
            O => \N__38514\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8\
        );

    \I__8245\ : LocalMux
    port map (
            O => \N__38511\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8\
        );

    \I__8244\ : LocalMux
    port map (
            O => \N__38508\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8\
        );

    \I__8243\ : InMux
    port map (
            O => \N__38501\,
            I => \N__38495\
        );

    \I__8242\ : InMux
    port map (
            O => \N__38500\,
            I => \N__38490\
        );

    \I__8241\ : InMux
    port map (
            O => \N__38499\,
            I => \N__38490\
        );

    \I__8240\ : InMux
    port map (
            O => \N__38498\,
            I => \N__38487\
        );

    \I__8239\ : LocalMux
    port map (
            O => \N__38495\,
            I => \N__38482\
        );

    \I__8238\ : LocalMux
    port map (
            O => \N__38490\,
            I => \N__38482\
        );

    \I__8237\ : LocalMux
    port map (
            O => \N__38487\,
            I => \N__38479\
        );

    \I__8236\ : Span4Mux_v
    port map (
            O => \N__38482\,
            I => \N__38476\
        );

    \I__8235\ : Odrv4
    port map (
            O => \N__38479\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__8234\ : Odrv4
    port map (
            O => \N__38476\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__8233\ : CascadeMux
    port map (
            O => \N__38471\,
            I => \N__38468\
        );

    \I__8232\ : InMux
    port map (
            O => \N__38468\,
            I => \N__38465\
        );

    \I__8231\ : LocalMux
    port map (
            O => \N__38465\,
            I => \N__38462\
        );

    \I__8230\ : Odrv4
    port map (
            O => \N__38462\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\
        );

    \I__8229\ : CascadeMux
    port map (
            O => \N__38459\,
            I => \N__38454\
        );

    \I__8228\ : InMux
    port map (
            O => \N__38458\,
            I => \N__38451\
        );

    \I__8227\ : InMux
    port map (
            O => \N__38457\,
            I => \N__38448\
        );

    \I__8226\ : InMux
    port map (
            O => \N__38454\,
            I => \N__38445\
        );

    \I__8225\ : LocalMux
    port map (
            O => \N__38451\,
            I => \N__38439\
        );

    \I__8224\ : LocalMux
    port map (
            O => \N__38448\,
            I => \N__38439\
        );

    \I__8223\ : LocalMux
    port map (
            O => \N__38445\,
            I => \N__38436\
        );

    \I__8222\ : InMux
    port map (
            O => \N__38444\,
            I => \N__38433\
        );

    \I__8221\ : Span4Mux_v
    port map (
            O => \N__38439\,
            I => \N__38428\
        );

    \I__8220\ : Span4Mux_v
    port map (
            O => \N__38436\,
            I => \N__38428\
        );

    \I__8219\ : LocalMux
    port map (
            O => \N__38433\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__8218\ : Odrv4
    port map (
            O => \N__38428\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__8217\ : InMux
    port map (
            O => \N__38423\,
            I => \N__38420\
        );

    \I__8216\ : LocalMux
    port map (
            O => \N__38420\,
            I => \N__38417\
        );

    \I__8215\ : Odrv4
    port map (
            O => \N__38417\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\
        );

    \I__8214\ : InMux
    port map (
            O => \N__38414\,
            I => \N__38410\
        );

    \I__8213\ : InMux
    port map (
            O => \N__38413\,
            I => \N__38407\
        );

    \I__8212\ : LocalMux
    port map (
            O => \N__38410\,
            I => \elapsed_time_ns_1_RNIV9PBB_0_21\
        );

    \I__8211\ : LocalMux
    port map (
            O => \N__38407\,
            I => \elapsed_time_ns_1_RNIV9PBB_0_21\
        );

    \I__8210\ : CascadeMux
    port map (
            O => \N__38402\,
            I => \elapsed_time_ns_1_RNIV9PBB_0_21_cascade_\
        );

    \I__8209\ : CascadeMux
    port map (
            O => \N__38399\,
            I => \N__38396\
        );

    \I__8208\ : InMux
    port map (
            O => \N__38396\,
            I => \N__38390\
        );

    \I__8207\ : InMux
    port map (
            O => \N__38395\,
            I => \N__38390\
        );

    \I__8206\ : LocalMux
    port map (
            O => \N__38390\,
            I => \N__38387\
        );

    \I__8205\ : Span4Mux_v
    port map (
            O => \N__38387\,
            I => \N__38384\
        );

    \I__8204\ : Odrv4
    port map (
            O => \N__38384\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_21\
        );

    \I__8203\ : CascadeMux
    port map (
            O => \N__38381\,
            I => \N__38378\
        );

    \I__8202\ : InMux
    port map (
            O => \N__38378\,
            I => \N__38375\
        );

    \I__8201\ : LocalMux
    port map (
            O => \N__38375\,
            I => \N__38372\
        );

    \I__8200\ : Odrv4
    port map (
            O => \N__38372\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\
        );

    \I__8199\ : InMux
    port map (
            O => \N__38369\,
            I => \N__38366\
        );

    \I__8198\ : LocalMux
    port map (
            O => \N__38366\,
            I => \N__38363\
        );

    \I__8197\ : Span4Mux_h
    port map (
            O => \N__38363\,
            I => \N__38360\
        );

    \I__8196\ : Odrv4
    port map (
            O => \N__38360\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15\
        );

    \I__8195\ : InMux
    port map (
            O => \N__38357\,
            I => \N__38353\
        );

    \I__8194\ : InMux
    port map (
            O => \N__38356\,
            I => \N__38350\
        );

    \I__8193\ : LocalMux
    port map (
            O => \N__38353\,
            I => \N__38347\
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__38350\,
            I => \N__38344\
        );

    \I__8191\ : Span4Mux_h
    port map (
            O => \N__38347\,
            I => \N__38339\
        );

    \I__8190\ : Span4Mux_h
    port map (
            O => \N__38344\,
            I => \N__38336\
        );

    \I__8189\ : InMux
    port map (
            O => \N__38343\,
            I => \N__38331\
        );

    \I__8188\ : InMux
    port map (
            O => \N__38342\,
            I => \N__38331\
        );

    \I__8187\ : Span4Mux_v
    port map (
            O => \N__38339\,
            I => \N__38328\
        );

    \I__8186\ : Odrv4
    port map (
            O => \N__38336\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__8185\ : LocalMux
    port map (
            O => \N__38331\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__8184\ : Odrv4
    port map (
            O => \N__38328\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__8183\ : CascadeMux
    port map (
            O => \N__38321\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22_cascade_\
        );

    \I__8182\ : InMux
    port map (
            O => \N__38318\,
            I => \N__38315\
        );

    \I__8181\ : LocalMux
    port map (
            O => \N__38315\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\
        );

    \I__8180\ : CascadeMux
    port map (
            O => \N__38312\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\
        );

    \I__8179\ : InMux
    port map (
            O => \N__38309\,
            I => \N__38305\
        );

    \I__8178\ : InMux
    port map (
            O => \N__38308\,
            I => \N__38302\
        );

    \I__8177\ : LocalMux
    port map (
            O => \N__38305\,
            I => \N__38295\
        );

    \I__8176\ : LocalMux
    port map (
            O => \N__38302\,
            I => \N__38295\
        );

    \I__8175\ : InMux
    port map (
            O => \N__38301\,
            I => \N__38292\
        );

    \I__8174\ : InMux
    port map (
            O => \N__38300\,
            I => \N__38289\
        );

    \I__8173\ : Span4Mux_h
    port map (
            O => \N__38295\,
            I => \N__38286\
        );

    \I__8172\ : LocalMux
    port map (
            O => \N__38292\,
            I => \N__38283\
        );

    \I__8171\ : LocalMux
    port map (
            O => \N__38289\,
            I => \N__38280\
        );

    \I__8170\ : Span4Mux_v
    port map (
            O => \N__38286\,
            I => \N__38277\
        );

    \I__8169\ : Span4Mux_v
    port map (
            O => \N__38283\,
            I => \N__38272\
        );

    \I__8168\ : Span4Mux_h
    port map (
            O => \N__38280\,
            I => \N__38272\
        );

    \I__8167\ : Odrv4
    port map (
            O => \N__38277\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\
        );

    \I__8166\ : Odrv4
    port map (
            O => \N__38272\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\
        );

    \I__8165\ : InMux
    port map (
            O => \N__38267\,
            I => \N__38259\
        );

    \I__8164\ : InMux
    port map (
            O => \N__38266\,
            I => \N__38259\
        );

    \I__8163\ : InMux
    port map (
            O => \N__38265\,
            I => \N__38256\
        );

    \I__8162\ : InMux
    port map (
            O => \N__38264\,
            I => \N__38253\
        );

    \I__8161\ : LocalMux
    port map (
            O => \N__38259\,
            I => \N__38250\
        );

    \I__8160\ : LocalMux
    port map (
            O => \N__38256\,
            I => \N__38247\
        );

    \I__8159\ : LocalMux
    port map (
            O => \N__38253\,
            I => \N__38244\
        );

    \I__8158\ : Span4Mux_v
    port map (
            O => \N__38250\,
            I => \N__38241\
        );

    \I__8157\ : Span4Mux_v
    port map (
            O => \N__38247\,
            I => \N__38236\
        );

    \I__8156\ : Span4Mux_h
    port map (
            O => \N__38244\,
            I => \N__38236\
        );

    \I__8155\ : Odrv4
    port map (
            O => \N__38241\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__8154\ : Odrv4
    port map (
            O => \N__38236\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__8153\ : CascadeMux
    port map (
            O => \N__38231\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3_cascade_\
        );

    \I__8152\ : InMux
    port map (
            O => \N__38228\,
            I => \N__38224\
        );

    \I__8151\ : InMux
    port map (
            O => \N__38227\,
            I => \N__38221\
        );

    \I__8150\ : LocalMux
    port map (
            O => \N__38224\,
            I => \N__38218\
        );

    \I__8149\ : LocalMux
    port map (
            O => \N__38221\,
            I => \N__38214\
        );

    \I__8148\ : Span4Mux_v
    port map (
            O => \N__38218\,
            I => \N__38210\
        );

    \I__8147\ : InMux
    port map (
            O => \N__38217\,
            I => \N__38207\
        );

    \I__8146\ : Span4Mux_h
    port map (
            O => \N__38214\,
            I => \N__38204\
        );

    \I__8145\ : InMux
    port map (
            O => \N__38213\,
            I => \N__38201\
        );

    \I__8144\ : Odrv4
    port map (
            O => \N__38210\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__8143\ : LocalMux
    port map (
            O => \N__38207\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__8142\ : Odrv4
    port map (
            O => \N__38204\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__8141\ : LocalMux
    port map (
            O => \N__38201\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__8140\ : InMux
    port map (
            O => \N__38192\,
            I => \N__38188\
        );

    \I__8139\ : InMux
    port map (
            O => \N__38191\,
            I => \N__38185\
        );

    \I__8138\ : LocalMux
    port map (
            O => \N__38188\,
            I => \N__38181\
        );

    \I__8137\ : LocalMux
    port map (
            O => \N__38185\,
            I => \N__38178\
        );

    \I__8136\ : InMux
    port map (
            O => \N__38184\,
            I => \N__38175\
        );

    \I__8135\ : Span4Mux_v
    port map (
            O => \N__38181\,
            I => \N__38170\
        );

    \I__8134\ : Span4Mux_h
    port map (
            O => \N__38178\,
            I => \N__38170\
        );

    \I__8133\ : LocalMux
    port map (
            O => \N__38175\,
            I => \elapsed_time_ns_1_RNIED91B_0_2\
        );

    \I__8132\ : Odrv4
    port map (
            O => \N__38170\,
            I => \elapsed_time_ns_1_RNIED91B_0_2\
        );

    \I__8131\ : InMux
    port map (
            O => \N__38165\,
            I => \N__38162\
        );

    \I__8130\ : LocalMux
    port map (
            O => \N__38162\,
            I => \N__38156\
        );

    \I__8129\ : InMux
    port map (
            O => \N__38161\,
            I => \N__38153\
        );

    \I__8128\ : InMux
    port map (
            O => \N__38160\,
            I => \N__38150\
        );

    \I__8127\ : InMux
    port map (
            O => \N__38159\,
            I => \N__38147\
        );

    \I__8126\ : Span4Mux_v
    port map (
            O => \N__38156\,
            I => \N__38144\
        );

    \I__8125\ : LocalMux
    port map (
            O => \N__38153\,
            I => \N__38141\
        );

    \I__8124\ : LocalMux
    port map (
            O => \N__38150\,
            I => \N__38138\
        );

    \I__8123\ : LocalMux
    port map (
            O => \N__38147\,
            I => \N__38135\
        );

    \I__8122\ : Span4Mux_v
    port map (
            O => \N__38144\,
            I => \N__38132\
        );

    \I__8121\ : Span4Mux_h
    port map (
            O => \N__38141\,
            I => \N__38127\
        );

    \I__8120\ : Span4Mux_h
    port map (
            O => \N__38138\,
            I => \N__38127\
        );

    \I__8119\ : Odrv12
    port map (
            O => \N__38135\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__8118\ : Odrv4
    port map (
            O => \N__38132\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__8117\ : Odrv4
    port map (
            O => \N__38127\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__8116\ : InMux
    port map (
            O => \N__38120\,
            I => \N__38115\
        );

    \I__8115\ : InMux
    port map (
            O => \N__38119\,
            I => \N__38112\
        );

    \I__8114\ : InMux
    port map (
            O => \N__38118\,
            I => \N__38109\
        );

    \I__8113\ : LocalMux
    port map (
            O => \N__38115\,
            I => \N__38106\
        );

    \I__8112\ : LocalMux
    port map (
            O => \N__38112\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3\
        );

    \I__8111\ : LocalMux
    port map (
            O => \N__38109\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3\
        );

    \I__8110\ : Odrv4
    port map (
            O => \N__38106\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3\
        );

    \I__8109\ : InMux
    port map (
            O => \N__38099\,
            I => \N__38094\
        );

    \I__8108\ : InMux
    port map (
            O => \N__38098\,
            I => \N__38091\
        );

    \I__8107\ : InMux
    port map (
            O => \N__38097\,
            I => \N__38088\
        );

    \I__8106\ : LocalMux
    port map (
            O => \N__38094\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6\
        );

    \I__8105\ : LocalMux
    port map (
            O => \N__38091\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6\
        );

    \I__8104\ : LocalMux
    port map (
            O => \N__38088\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6\
        );

    \I__8103\ : InMux
    port map (
            O => \N__38081\,
            I => \N__38076\
        );

    \I__8102\ : InMux
    port map (
            O => \N__38080\,
            I => \N__38073\
        );

    \I__8101\ : InMux
    port map (
            O => \N__38079\,
            I => \N__38070\
        );

    \I__8100\ : LocalMux
    port map (
            O => \N__38076\,
            I => \N__38067\
        );

    \I__8099\ : LocalMux
    port map (
            O => \N__38073\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__8098\ : LocalMux
    port map (
            O => \N__38070\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__8097\ : Odrv4
    port map (
            O => \N__38067\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__8096\ : CascadeMux
    port map (
            O => \N__38060\,
            I => \N__38057\
        );

    \I__8095\ : InMux
    port map (
            O => \N__38057\,
            I => \N__38050\
        );

    \I__8094\ : InMux
    port map (
            O => \N__38056\,
            I => \N__38050\
        );

    \I__8093\ : InMux
    port map (
            O => \N__38055\,
            I => \N__38047\
        );

    \I__8092\ : LocalMux
    port map (
            O => \N__38050\,
            I => \N__38043\
        );

    \I__8091\ : LocalMux
    port map (
            O => \N__38047\,
            I => \N__38040\
        );

    \I__8090\ : InMux
    port map (
            O => \N__38046\,
            I => \N__38037\
        );

    \I__8089\ : Span4Mux_v
    port map (
            O => \N__38043\,
            I => \N__38034\
        );

    \I__8088\ : Span4Mux_h
    port map (
            O => \N__38040\,
            I => \N__38031\
        );

    \I__8087\ : LocalMux
    port map (
            O => \N__38037\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__8086\ : Odrv4
    port map (
            O => \N__38034\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__8085\ : Odrv4
    port map (
            O => \N__38031\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__8084\ : InMux
    port map (
            O => \N__38024\,
            I => \N__38021\
        );

    \I__8083\ : LocalMux
    port map (
            O => \N__38021\,
            I => \N__38017\
        );

    \I__8082\ : InMux
    port map (
            O => \N__38020\,
            I => \N__38014\
        );

    \I__8081\ : Span4Mux_v
    port map (
            O => \N__38017\,
            I => \N__38011\
        );

    \I__8080\ : LocalMux
    port map (
            O => \N__38014\,
            I => \N__38008\
        );

    \I__8079\ : Odrv4
    port map (
            O => \N__38011\,
            I => \phase_controller_inst1.time_passed_RNI7NN7\
        );

    \I__8078\ : Odrv4
    port map (
            O => \N__38008\,
            I => \phase_controller_inst1.time_passed_RNI7NN7\
        );

    \I__8077\ : InMux
    port map (
            O => \N__38003\,
            I => \N__37987\
        );

    \I__8076\ : InMux
    port map (
            O => \N__38002\,
            I => \N__37984\
        );

    \I__8075\ : InMux
    port map (
            O => \N__38001\,
            I => \N__37981\
        );

    \I__8074\ : CascadeMux
    port map (
            O => \N__38000\,
            I => \N__37972\
        );

    \I__8073\ : CascadeMux
    port map (
            O => \N__37999\,
            I => \N__37968\
        );

    \I__8072\ : CascadeMux
    port map (
            O => \N__37998\,
            I => \N__37964\
        );

    \I__8071\ : CascadeMux
    port map (
            O => \N__37997\,
            I => \N__37960\
        );

    \I__8070\ : CascadeMux
    port map (
            O => \N__37996\,
            I => \N__37956\
        );

    \I__8069\ : CascadeMux
    port map (
            O => \N__37995\,
            I => \N__37952\
        );

    \I__8068\ : CascadeMux
    port map (
            O => \N__37994\,
            I => \N__37948\
        );

    \I__8067\ : CascadeMux
    port map (
            O => \N__37993\,
            I => \N__37944\
        );

    \I__8066\ : CascadeMux
    port map (
            O => \N__37992\,
            I => \N__37940\
        );

    \I__8065\ : CascadeMux
    port map (
            O => \N__37991\,
            I => \N__37936\
        );

    \I__8064\ : CascadeMux
    port map (
            O => \N__37990\,
            I => \N__37932\
        );

    \I__8063\ : LocalMux
    port map (
            O => \N__37987\,
            I => \N__37921\
        );

    \I__8062\ : LocalMux
    port map (
            O => \N__37984\,
            I => \N__37921\
        );

    \I__8061\ : LocalMux
    port map (
            O => \N__37981\,
            I => \N__37921\
        );

    \I__8060\ : InMux
    port map (
            O => \N__37980\,
            I => \N__37918\
        );

    \I__8059\ : InMux
    port map (
            O => \N__37979\,
            I => \N__37914\
        );

    \I__8058\ : InMux
    port map (
            O => \N__37978\,
            I => \N__37909\
        );

    \I__8057\ : InMux
    port map (
            O => \N__37977\,
            I => \N__37909\
        );

    \I__8056\ : InMux
    port map (
            O => \N__37976\,
            I => \N__37906\
        );

    \I__8055\ : InMux
    port map (
            O => \N__37975\,
            I => \N__37894\
        );

    \I__8054\ : InMux
    port map (
            O => \N__37972\,
            I => \N__37879\
        );

    \I__8053\ : InMux
    port map (
            O => \N__37971\,
            I => \N__37879\
        );

    \I__8052\ : InMux
    port map (
            O => \N__37968\,
            I => \N__37879\
        );

    \I__8051\ : InMux
    port map (
            O => \N__37967\,
            I => \N__37879\
        );

    \I__8050\ : InMux
    port map (
            O => \N__37964\,
            I => \N__37879\
        );

    \I__8049\ : InMux
    port map (
            O => \N__37963\,
            I => \N__37879\
        );

    \I__8048\ : InMux
    port map (
            O => \N__37960\,
            I => \N__37879\
        );

    \I__8047\ : InMux
    port map (
            O => \N__37959\,
            I => \N__37864\
        );

    \I__8046\ : InMux
    port map (
            O => \N__37956\,
            I => \N__37864\
        );

    \I__8045\ : InMux
    port map (
            O => \N__37955\,
            I => \N__37864\
        );

    \I__8044\ : InMux
    port map (
            O => \N__37952\,
            I => \N__37864\
        );

    \I__8043\ : InMux
    port map (
            O => \N__37951\,
            I => \N__37864\
        );

    \I__8042\ : InMux
    port map (
            O => \N__37948\,
            I => \N__37864\
        );

    \I__8041\ : InMux
    port map (
            O => \N__37947\,
            I => \N__37864\
        );

    \I__8040\ : InMux
    port map (
            O => \N__37944\,
            I => \N__37847\
        );

    \I__8039\ : InMux
    port map (
            O => \N__37943\,
            I => \N__37847\
        );

    \I__8038\ : InMux
    port map (
            O => \N__37940\,
            I => \N__37847\
        );

    \I__8037\ : InMux
    port map (
            O => \N__37939\,
            I => \N__37847\
        );

    \I__8036\ : InMux
    port map (
            O => \N__37936\,
            I => \N__37847\
        );

    \I__8035\ : InMux
    port map (
            O => \N__37935\,
            I => \N__37847\
        );

    \I__8034\ : InMux
    port map (
            O => \N__37932\,
            I => \N__37847\
        );

    \I__8033\ : InMux
    port map (
            O => \N__37931\,
            I => \N__37847\
        );

    \I__8032\ : InMux
    port map (
            O => \N__37930\,
            I => \N__37840\
        );

    \I__8031\ : InMux
    port map (
            O => \N__37929\,
            I => \N__37835\
        );

    \I__8030\ : InMux
    port map (
            O => \N__37928\,
            I => \N__37835\
        );

    \I__8029\ : Span4Mux_s2_v
    port map (
            O => \N__37921\,
            I => \N__37830\
        );

    \I__8028\ : LocalMux
    port map (
            O => \N__37918\,
            I => \N__37830\
        );

    \I__8027\ : CascadeMux
    port map (
            O => \N__37917\,
            I => \N__37819\
        );

    \I__8026\ : LocalMux
    port map (
            O => \N__37914\,
            I => \N__37815\
        );

    \I__8025\ : LocalMux
    port map (
            O => \N__37909\,
            I => \N__37810\
        );

    \I__8024\ : LocalMux
    port map (
            O => \N__37906\,
            I => \N__37810\
        );

    \I__8023\ : InMux
    port map (
            O => \N__37905\,
            I => \N__37807\
        );

    \I__8022\ : InMux
    port map (
            O => \N__37904\,
            I => \N__37804\
        );

    \I__8021\ : InMux
    port map (
            O => \N__37903\,
            I => \N__37797\
        );

    \I__8020\ : InMux
    port map (
            O => \N__37902\,
            I => \N__37797\
        );

    \I__8019\ : InMux
    port map (
            O => \N__37901\,
            I => \N__37797\
        );

    \I__8018\ : InMux
    port map (
            O => \N__37900\,
            I => \N__37788\
        );

    \I__8017\ : InMux
    port map (
            O => \N__37899\,
            I => \N__37788\
        );

    \I__8016\ : InMux
    port map (
            O => \N__37898\,
            I => \N__37788\
        );

    \I__8015\ : InMux
    port map (
            O => \N__37897\,
            I => \N__37788\
        );

    \I__8014\ : LocalMux
    port map (
            O => \N__37894\,
            I => \N__37785\
        );

    \I__8013\ : LocalMux
    port map (
            O => \N__37879\,
            I => \N__37782\
        );

    \I__8012\ : LocalMux
    port map (
            O => \N__37864\,
            I => \N__37777\
        );

    \I__8011\ : LocalMux
    port map (
            O => \N__37847\,
            I => \N__37777\
        );

    \I__8010\ : CascadeMux
    port map (
            O => \N__37846\,
            I => \N__37774\
        );

    \I__8009\ : CascadeMux
    port map (
            O => \N__37845\,
            I => \N__37770\
        );

    \I__8008\ : CascadeMux
    port map (
            O => \N__37844\,
            I => \N__37766\
        );

    \I__8007\ : CascadeMux
    port map (
            O => \N__37843\,
            I => \N__37762\
        );

    \I__8006\ : LocalMux
    port map (
            O => \N__37840\,
            I => \N__37756\
        );

    \I__8005\ : LocalMux
    port map (
            O => \N__37835\,
            I => \N__37753\
        );

    \I__8004\ : Span4Mux_v
    port map (
            O => \N__37830\,
            I => \N__37750\
        );

    \I__8003\ : InMux
    port map (
            O => \N__37829\,
            I => \N__37743\
        );

    \I__8002\ : InMux
    port map (
            O => \N__37828\,
            I => \N__37743\
        );

    \I__8001\ : InMux
    port map (
            O => \N__37827\,
            I => \N__37743\
        );

    \I__8000\ : InMux
    port map (
            O => \N__37826\,
            I => \N__37734\
        );

    \I__7999\ : InMux
    port map (
            O => \N__37825\,
            I => \N__37734\
        );

    \I__7998\ : InMux
    port map (
            O => \N__37824\,
            I => \N__37734\
        );

    \I__7997\ : InMux
    port map (
            O => \N__37823\,
            I => \N__37734\
        );

    \I__7996\ : InMux
    port map (
            O => \N__37822\,
            I => \N__37727\
        );

    \I__7995\ : InMux
    port map (
            O => \N__37819\,
            I => \N__37727\
        );

    \I__7994\ : InMux
    port map (
            O => \N__37818\,
            I => \N__37727\
        );

    \I__7993\ : Span4Mux_v
    port map (
            O => \N__37815\,
            I => \N__37720\
        );

    \I__7992\ : Span4Mux_v
    port map (
            O => \N__37810\,
            I => \N__37720\
        );

    \I__7991\ : LocalMux
    port map (
            O => \N__37807\,
            I => \N__37720\
        );

    \I__7990\ : LocalMux
    port map (
            O => \N__37804\,
            I => \N__37711\
        );

    \I__7989\ : LocalMux
    port map (
            O => \N__37797\,
            I => \N__37711\
        );

    \I__7988\ : LocalMux
    port map (
            O => \N__37788\,
            I => \N__37711\
        );

    \I__7987\ : Span12Mux_s2_v
    port map (
            O => \N__37785\,
            I => \N__37711\
        );

    \I__7986\ : Span4Mux_v
    port map (
            O => \N__37782\,
            I => \N__37706\
        );

    \I__7985\ : Span4Mux_v
    port map (
            O => \N__37777\,
            I => \N__37706\
        );

    \I__7984\ : InMux
    port map (
            O => \N__37774\,
            I => \N__37689\
        );

    \I__7983\ : InMux
    port map (
            O => \N__37773\,
            I => \N__37689\
        );

    \I__7982\ : InMux
    port map (
            O => \N__37770\,
            I => \N__37689\
        );

    \I__7981\ : InMux
    port map (
            O => \N__37769\,
            I => \N__37689\
        );

    \I__7980\ : InMux
    port map (
            O => \N__37766\,
            I => \N__37689\
        );

    \I__7979\ : InMux
    port map (
            O => \N__37765\,
            I => \N__37689\
        );

    \I__7978\ : InMux
    port map (
            O => \N__37762\,
            I => \N__37689\
        );

    \I__7977\ : InMux
    port map (
            O => \N__37761\,
            I => \N__37689\
        );

    \I__7976\ : InMux
    port map (
            O => \N__37760\,
            I => \N__37684\
        );

    \I__7975\ : InMux
    port map (
            O => \N__37759\,
            I => \N__37684\
        );

    \I__7974\ : Span4Mux_s1_h
    port map (
            O => \N__37756\,
            I => \N__37679\
        );

    \I__7973\ : Span4Mux_v
    port map (
            O => \N__37753\,
            I => \N__37679\
        );

    \I__7972\ : Sp12to4
    port map (
            O => \N__37750\,
            I => \N__37670\
        );

    \I__7971\ : LocalMux
    port map (
            O => \N__37743\,
            I => \N__37670\
        );

    \I__7970\ : LocalMux
    port map (
            O => \N__37734\,
            I => \N__37670\
        );

    \I__7969\ : LocalMux
    port map (
            O => \N__37727\,
            I => \N__37670\
        );

    \I__7968\ : Sp12to4
    port map (
            O => \N__37720\,
            I => \N__37667\
        );

    \I__7967\ : Span12Mux_v
    port map (
            O => \N__37711\,
            I => \N__37660\
        );

    \I__7966\ : Sp12to4
    port map (
            O => \N__37706\,
            I => \N__37660\
        );

    \I__7965\ : LocalMux
    port map (
            O => \N__37689\,
            I => \N__37660\
        );

    \I__7964\ : LocalMux
    port map (
            O => \N__37684\,
            I => \N__37657\
        );

    \I__7963\ : Span4Mux_h
    port map (
            O => \N__37679\,
            I => \N__37654\
        );

    \I__7962\ : Span12Mux_s5_h
    port map (
            O => \N__37670\,
            I => \N__37651\
        );

    \I__7961\ : Span12Mux_v
    port map (
            O => \N__37667\,
            I => \N__37644\
        );

    \I__7960\ : Span12Mux_h
    port map (
            O => \N__37660\,
            I => \N__37644\
        );

    \I__7959\ : Span12Mux_v
    port map (
            O => \N__37657\,
            I => \N__37644\
        );

    \I__7958\ : Odrv4
    port map (
            O => \N__37654\,
            I => \CONSTANT_ONE_NET\
        );

    \I__7957\ : Odrv12
    port map (
            O => \N__37651\,
            I => \CONSTANT_ONE_NET\
        );

    \I__7956\ : Odrv12
    port map (
            O => \N__37644\,
            I => \CONSTANT_ONE_NET\
        );

    \I__7955\ : InMux
    port map (
            O => \N__37637\,
            I => \current_shift_inst.un10_control_input_cry_30\
        );

    \I__7954\ : InMux
    port map (
            O => \N__37634\,
            I => \N__37628\
        );

    \I__7953\ : CascadeMux
    port map (
            O => \N__37633\,
            I => \N__37625\
        );

    \I__7952\ : InMux
    port map (
            O => \N__37632\,
            I => \N__37616\
        );

    \I__7951\ : InMux
    port map (
            O => \N__37631\,
            I => \N__37616\
        );

    \I__7950\ : LocalMux
    port map (
            O => \N__37628\,
            I => \N__37613\
        );

    \I__7949\ : InMux
    port map (
            O => \N__37625\,
            I => \N__37610\
        );

    \I__7948\ : InMux
    port map (
            O => \N__37624\,
            I => \N__37607\
        );

    \I__7947\ : InMux
    port map (
            O => \N__37623\,
            I => \N__37602\
        );

    \I__7946\ : InMux
    port map (
            O => \N__37622\,
            I => \N__37602\
        );

    \I__7945\ : CascadeMux
    port map (
            O => \N__37621\,
            I => \N__37595\
        );

    \I__7944\ : LocalMux
    port map (
            O => \N__37616\,
            I => \N__37590\
        );

    \I__7943\ : Span4Mux_v
    port map (
            O => \N__37613\,
            I => \N__37586\
        );

    \I__7942\ : LocalMux
    port map (
            O => \N__37610\,
            I => \N__37583\
        );

    \I__7941\ : LocalMux
    port map (
            O => \N__37607\,
            I => \N__37578\
        );

    \I__7940\ : LocalMux
    port map (
            O => \N__37602\,
            I => \N__37578\
        );

    \I__7939\ : InMux
    port map (
            O => \N__37601\,
            I => \N__37563\
        );

    \I__7938\ : InMux
    port map (
            O => \N__37600\,
            I => \N__37563\
        );

    \I__7937\ : InMux
    port map (
            O => \N__37599\,
            I => \N__37563\
        );

    \I__7936\ : InMux
    port map (
            O => \N__37598\,
            I => \N__37563\
        );

    \I__7935\ : InMux
    port map (
            O => \N__37595\,
            I => \N__37563\
        );

    \I__7934\ : InMux
    port map (
            O => \N__37594\,
            I => \N__37563\
        );

    \I__7933\ : InMux
    port map (
            O => \N__37593\,
            I => \N__37563\
        );

    \I__7932\ : Span4Mux_h
    port map (
            O => \N__37590\,
            I => \N__37560\
        );

    \I__7931\ : InMux
    port map (
            O => \N__37589\,
            I => \N__37557\
        );

    \I__7930\ : Span4Mux_h
    port map (
            O => \N__37586\,
            I => \N__37552\
        );

    \I__7929\ : Span4Mux_v
    port map (
            O => \N__37583\,
            I => \N__37552\
        );

    \I__7928\ : Span4Mux_v
    port map (
            O => \N__37578\,
            I => \N__37547\
        );

    \I__7927\ : LocalMux
    port map (
            O => \N__37563\,
            I => \N__37547\
        );

    \I__7926\ : Span4Mux_h
    port map (
            O => \N__37560\,
            I => \N__37544\
        );

    \I__7925\ : LocalMux
    port map (
            O => \N__37557\,
            I => \N__37541\
        );

    \I__7924\ : Odrv4
    port map (
            O => \N__37552\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__7923\ : Odrv4
    port map (
            O => \N__37547\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__7922\ : Odrv4
    port map (
            O => \N__37544\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__7921\ : Odrv12
    port map (
            O => \N__37541\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__7920\ : InMux
    port map (
            O => \N__37532\,
            I => \N__37529\
        );

    \I__7919\ : LocalMux
    port map (
            O => \N__37529\,
            I => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\
        );

    \I__7918\ : CascadeMux
    port map (
            O => \N__37526\,
            I => \N__37523\
        );

    \I__7917\ : InMux
    port map (
            O => \N__37523\,
            I => \N__37520\
        );

    \I__7916\ : LocalMux
    port map (
            O => \N__37520\,
            I => \N__37517\
        );

    \I__7915\ : Span4Mux_v
    port map (
            O => \N__37517\,
            I => \N__37514\
        );

    \I__7914\ : Odrv4
    port map (
            O => \N__37514\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30\
        );

    \I__7913\ : InMux
    port map (
            O => \N__37511\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_28\
        );

    \I__7912\ : InMux
    port map (
            O => \N__37508\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_30\
        );

    \I__7911\ : CascadeMux
    port map (
            O => \N__37505\,
            I => \N__37502\
        );

    \I__7910\ : InMux
    port map (
            O => \N__37502\,
            I => \N__37498\
        );

    \I__7909\ : InMux
    port map (
            O => \N__37501\,
            I => \N__37495\
        );

    \I__7908\ : LocalMux
    port map (
            O => \N__37498\,
            I => \N__37492\
        );

    \I__7907\ : LocalMux
    port map (
            O => \N__37495\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__7906\ : Odrv12
    port map (
            O => \N__37492\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__7905\ : CascadeMux
    port map (
            O => \N__37487\,
            I => \N__37484\
        );

    \I__7904\ : InMux
    port map (
            O => \N__37484\,
            I => \N__37481\
        );

    \I__7903\ : LocalMux
    port map (
            O => \N__37481\,
            I => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\
        );

    \I__7902\ : CascadeMux
    port map (
            O => \N__37478\,
            I => \N__37475\
        );

    \I__7901\ : InMux
    port map (
            O => \N__37475\,
            I => \N__37472\
        );

    \I__7900\ : LocalMux
    port map (
            O => \N__37472\,
            I => \N__37469\
        );

    \I__7899\ : Odrv4
    port map (
            O => \N__37469\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\
        );

    \I__7898\ : CascadeMux
    port map (
            O => \N__37466\,
            I => \N__37463\
        );

    \I__7897\ : InMux
    port map (
            O => \N__37463\,
            I => \N__37460\
        );

    \I__7896\ : LocalMux
    port map (
            O => \N__37460\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\
        );

    \I__7895\ : InMux
    port map (
            O => \N__37457\,
            I => \N__37454\
        );

    \I__7894\ : LocalMux
    port map (
            O => \N__37454\,
            I => \N__37451\
        );

    \I__7893\ : Odrv4
    port map (
            O => \N__37451\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20\
        );

    \I__7892\ : CascadeMux
    port map (
            O => \N__37448\,
            I => \N__37445\
        );

    \I__7891\ : InMux
    port map (
            O => \N__37445\,
            I => \N__37442\
        );

    \I__7890\ : LocalMux
    port map (
            O => \N__37442\,
            I => \N__37439\
        );

    \I__7889\ : Span4Mux_v
    port map (
            O => \N__37439\,
            I => \N__37436\
        );

    \I__7888\ : Odrv4
    port map (
            O => \N__37436\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt20\
        );

    \I__7887\ : InMux
    port map (
            O => \N__37433\,
            I => \N__37430\
        );

    \I__7886\ : LocalMux
    port map (
            O => \N__37430\,
            I => \N__37427\
        );

    \I__7885\ : Odrv12
    port map (
            O => \N__37427\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\
        );

    \I__7884\ : CascadeMux
    port map (
            O => \N__37424\,
            I => \N__37421\
        );

    \I__7883\ : InMux
    port map (
            O => \N__37421\,
            I => \N__37418\
        );

    \I__7882\ : LocalMux
    port map (
            O => \N__37418\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\
        );

    \I__7881\ : CascadeMux
    port map (
            O => \N__37415\,
            I => \N__37412\
        );

    \I__7880\ : InMux
    port map (
            O => \N__37412\,
            I => \N__37409\
        );

    \I__7879\ : LocalMux
    port map (
            O => \N__37409\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\
        );

    \I__7878\ : InMux
    port map (
            O => \N__37406\,
            I => \N__37403\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__37403\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\
        );

    \I__7876\ : InMux
    port map (
            O => \N__37400\,
            I => \N__37397\
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__37397\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\
        );

    \I__7874\ : CascadeMux
    port map (
            O => \N__37394\,
            I => \N__37391\
        );

    \I__7873\ : InMux
    port map (
            O => \N__37391\,
            I => \N__37388\
        );

    \I__7872\ : LocalMux
    port map (
            O => \N__37388\,
            I => \N__37385\
        );

    \I__7871\ : Odrv4
    port map (
            O => \N__37385\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\
        );

    \I__7870\ : InMux
    port map (
            O => \N__37382\,
            I => \N__37379\
        );

    \I__7869\ : LocalMux
    port map (
            O => \N__37379\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\
        );

    \I__7868\ : InMux
    port map (
            O => \N__37376\,
            I => \N__37373\
        );

    \I__7867\ : LocalMux
    port map (
            O => \N__37373\,
            I => \N__37370\
        );

    \I__7866\ : Odrv12
    port map (
            O => \N__37370\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\
        );

    \I__7865\ : CascadeMux
    port map (
            O => \N__37367\,
            I => \N__37364\
        );

    \I__7864\ : InMux
    port map (
            O => \N__37364\,
            I => \N__37361\
        );

    \I__7863\ : LocalMux
    port map (
            O => \N__37361\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\
        );

    \I__7862\ : InMux
    port map (
            O => \N__37358\,
            I => \N__37355\
        );

    \I__7861\ : LocalMux
    port map (
            O => \N__37355\,
            I => \N__37352\
        );

    \I__7860\ : Odrv4
    port map (
            O => \N__37352\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\
        );

    \I__7859\ : CascadeMux
    port map (
            O => \N__37349\,
            I => \N__37346\
        );

    \I__7858\ : InMux
    port map (
            O => \N__37346\,
            I => \N__37343\
        );

    \I__7857\ : LocalMux
    port map (
            O => \N__37343\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\
        );

    \I__7856\ : CascadeMux
    port map (
            O => \N__37340\,
            I => \N__37337\
        );

    \I__7855\ : InMux
    port map (
            O => \N__37337\,
            I => \N__37334\
        );

    \I__7854\ : LocalMux
    port map (
            O => \N__37334\,
            I => \N__37331\
        );

    \I__7853\ : Odrv4
    port map (
            O => \N__37331\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\
        );

    \I__7852\ : InMux
    port map (
            O => \N__37328\,
            I => \N__37325\
        );

    \I__7851\ : LocalMux
    port map (
            O => \N__37325\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\
        );

    \I__7850\ : InMux
    port map (
            O => \N__37322\,
            I => \N__37316\
        );

    \I__7849\ : InMux
    port map (
            O => \N__37321\,
            I => \N__37316\
        );

    \I__7848\ : LocalMux
    port map (
            O => \N__37316\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_20\
        );

    \I__7847\ : InMux
    port map (
            O => \N__37313\,
            I => \N__37310\
        );

    \I__7846\ : LocalMux
    port map (
            O => \N__37310\,
            I => \N__37306\
        );

    \I__7845\ : InMux
    port map (
            O => \N__37309\,
            I => \N__37302\
        );

    \I__7844\ : Span4Mux_v
    port map (
            O => \N__37306\,
            I => \N__37299\
        );

    \I__7843\ : InMux
    port map (
            O => \N__37305\,
            I => \N__37296\
        );

    \I__7842\ : LocalMux
    port map (
            O => \N__37302\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__7841\ : Odrv4
    port map (
            O => \N__37299\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__7840\ : LocalMux
    port map (
            O => \N__37296\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__7839\ : InMux
    port map (
            O => \N__37289\,
            I => \N__37286\
        );

    \I__7838\ : LocalMux
    port map (
            O => \N__37286\,
            I => \N__37283\
        );

    \I__7837\ : Span4Mux_v
    port map (
            O => \N__37283\,
            I => \N__37277\
        );

    \I__7836\ : InMux
    port map (
            O => \N__37282\,
            I => \N__37274\
        );

    \I__7835\ : InMux
    port map (
            O => \N__37281\,
            I => \N__37269\
        );

    \I__7834\ : InMux
    port map (
            O => \N__37280\,
            I => \N__37269\
        );

    \I__7833\ : Odrv4
    port map (
            O => \N__37277\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__7832\ : LocalMux
    port map (
            O => \N__37274\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__7831\ : LocalMux
    port map (
            O => \N__37269\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__7830\ : CascadeMux
    port map (
            O => \N__37262\,
            I => \N__37257\
        );

    \I__7829\ : InMux
    port map (
            O => \N__37261\,
            I => \N__37254\
        );

    \I__7828\ : InMux
    port map (
            O => \N__37260\,
            I => \N__37251\
        );

    \I__7827\ : InMux
    port map (
            O => \N__37257\,
            I => \N__37248\
        );

    \I__7826\ : LocalMux
    port map (
            O => \N__37254\,
            I => \N__37244\
        );

    \I__7825\ : LocalMux
    port map (
            O => \N__37251\,
            I => \N__37241\
        );

    \I__7824\ : LocalMux
    port map (
            O => \N__37248\,
            I => \N__37238\
        );

    \I__7823\ : InMux
    port map (
            O => \N__37247\,
            I => \N__37235\
        );

    \I__7822\ : Span4Mux_v
    port map (
            O => \N__37244\,
            I => \N__37230\
        );

    \I__7821\ : Span4Mux_h
    port map (
            O => \N__37241\,
            I => \N__37230\
        );

    \I__7820\ : Span4Mux_h
    port map (
            O => \N__37238\,
            I => \N__37227\
        );

    \I__7819\ : LocalMux
    port map (
            O => \N__37235\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__7818\ : Odrv4
    port map (
            O => \N__37230\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__7817\ : Odrv4
    port map (
            O => \N__37227\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__7816\ : InMux
    port map (
            O => \N__37220\,
            I => \N__37217\
        );

    \I__7815\ : LocalMux
    port map (
            O => \N__37217\,
            I => \N__37213\
        );

    \I__7814\ : InMux
    port map (
            O => \N__37216\,
            I => \N__37209\
        );

    \I__7813\ : Span4Mux_h
    port map (
            O => \N__37213\,
            I => \N__37206\
        );

    \I__7812\ : InMux
    port map (
            O => \N__37212\,
            I => \N__37203\
        );

    \I__7811\ : LocalMux
    port map (
            O => \N__37209\,
            I => \N__37198\
        );

    \I__7810\ : Span4Mux_h
    port map (
            O => \N__37206\,
            I => \N__37198\
        );

    \I__7809\ : LocalMux
    port map (
            O => \N__37203\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4\
        );

    \I__7808\ : Odrv4
    port map (
            O => \N__37198\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4\
        );

    \I__7807\ : CascadeMux
    port map (
            O => \N__37193\,
            I => \N__37190\
        );

    \I__7806\ : InMux
    port map (
            O => \N__37190\,
            I => \N__37187\
        );

    \I__7805\ : LocalMux
    port map (
            O => \N__37187\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\
        );

    \I__7804\ : InMux
    port map (
            O => \N__37184\,
            I => \N__37181\
        );

    \I__7803\ : LocalMux
    port map (
            O => \N__37181\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\
        );

    \I__7802\ : InMux
    port map (
            O => \N__37178\,
            I => \N__37175\
        );

    \I__7801\ : LocalMux
    port map (
            O => \N__37175\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\
        );

    \I__7800\ : CascadeMux
    port map (
            O => \N__37172\,
            I => \N__37169\
        );

    \I__7799\ : InMux
    port map (
            O => \N__37169\,
            I => \N__37166\
        );

    \I__7798\ : LocalMux
    port map (
            O => \N__37166\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\
        );

    \I__7797\ : InMux
    port map (
            O => \N__37163\,
            I => \N__37160\
        );

    \I__7796\ : LocalMux
    port map (
            O => \N__37160\,
            I => \N__37157\
        );

    \I__7795\ : Span4Mux_v
    port map (
            O => \N__37157\,
            I => \N__37154\
        );

    \I__7794\ : Odrv4
    port map (
            O => \N__37154\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\
        );

    \I__7793\ : CascadeMux
    port map (
            O => \N__37151\,
            I => \N__37148\
        );

    \I__7792\ : InMux
    port map (
            O => \N__37148\,
            I => \N__37145\
        );

    \I__7791\ : LocalMux
    port map (
            O => \N__37145\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\
        );

    \I__7790\ : CascadeMux
    port map (
            O => \N__37142\,
            I => \N__37139\
        );

    \I__7789\ : InMux
    port map (
            O => \N__37139\,
            I => \N__37136\
        );

    \I__7788\ : LocalMux
    port map (
            O => \N__37136\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\
        );

    \I__7787\ : InMux
    port map (
            O => \N__37133\,
            I => \N__37130\
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__37130\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\
        );

    \I__7785\ : InMux
    port map (
            O => \N__37127\,
            I => \N__37124\
        );

    \I__7784\ : LocalMux
    port map (
            O => \N__37124\,
            I => \N__37121\
        );

    \I__7783\ : Span4Mux_v
    port map (
            O => \N__37121\,
            I => \N__37118\
        );

    \I__7782\ : Odrv4
    port map (
            O => \N__37118\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\
        );

    \I__7781\ : CascadeMux
    port map (
            O => \N__37115\,
            I => \N__37112\
        );

    \I__7780\ : InMux
    port map (
            O => \N__37112\,
            I => \N__37109\
        );

    \I__7779\ : LocalMux
    port map (
            O => \N__37109\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\
        );

    \I__7778\ : CascadeMux
    port map (
            O => \N__37106\,
            I => \N__37103\
        );

    \I__7777\ : InMux
    port map (
            O => \N__37103\,
            I => \N__37100\
        );

    \I__7776\ : LocalMux
    port map (
            O => \N__37100\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\
        );

    \I__7775\ : InMux
    port map (
            O => \N__37097\,
            I => \N__37093\
        );

    \I__7774\ : InMux
    port map (
            O => \N__37096\,
            I => \N__37090\
        );

    \I__7773\ : LocalMux
    port map (
            O => \N__37093\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11\
        );

    \I__7772\ : LocalMux
    port map (
            O => \N__37090\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11\
        );

    \I__7771\ : CascadeMux
    port map (
            O => \N__37085\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11_cascade_\
        );

    \I__7770\ : InMux
    port map (
            O => \N__37082\,
            I => \N__37079\
        );

    \I__7769\ : LocalMux
    port map (
            O => \N__37079\,
            I => \N__37075\
        );

    \I__7768\ : InMux
    port map (
            O => \N__37078\,
            I => \N__37072\
        );

    \I__7767\ : Odrv4
    port map (
            O => \N__37075\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10\
        );

    \I__7766\ : LocalMux
    port map (
            O => \N__37072\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10\
        );

    \I__7765\ : CascadeMux
    port map (
            O => \N__37067\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10_cascade_\
        );

    \I__7764\ : InMux
    port map (
            O => \N__37064\,
            I => \N__37061\
        );

    \I__7763\ : LocalMux
    port map (
            O => \N__37061\,
            I => \N__37055\
        );

    \I__7762\ : InMux
    port map (
            O => \N__37060\,
            I => \N__37048\
        );

    \I__7761\ : InMux
    port map (
            O => \N__37059\,
            I => \N__37048\
        );

    \I__7760\ : InMux
    port map (
            O => \N__37058\,
            I => \N__37048\
        );

    \I__7759\ : Span4Mux_h
    port map (
            O => \N__37055\,
            I => \N__37043\
        );

    \I__7758\ : LocalMux
    port map (
            O => \N__37048\,
            I => \N__37043\
        );

    \I__7757\ : Odrv4
    port map (
            O => \N__37043\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__7756\ : InMux
    port map (
            O => \N__37040\,
            I => \N__37037\
        );

    \I__7755\ : LocalMux
    port map (
            O => \N__37037\,
            I => \N__37034\
        );

    \I__7754\ : Span4Mux_h
    port map (
            O => \N__37034\,
            I => \N__37028\
        );

    \I__7753\ : InMux
    port map (
            O => \N__37033\,
            I => \N__37021\
        );

    \I__7752\ : InMux
    port map (
            O => \N__37032\,
            I => \N__37021\
        );

    \I__7751\ : InMux
    port map (
            O => \N__37031\,
            I => \N__37021\
        );

    \I__7750\ : Odrv4
    port map (
            O => \N__37028\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__7749\ : LocalMux
    port map (
            O => \N__37021\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__7748\ : InMux
    port map (
            O => \N__37016\,
            I => \N__37010\
        );

    \I__7747\ : InMux
    port map (
            O => \N__37015\,
            I => \N__37010\
        );

    \I__7746\ : LocalMux
    port map (
            O => \N__37010\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_20\
        );

    \I__7745\ : InMux
    port map (
            O => \N__37007\,
            I => \N__37004\
        );

    \I__7744\ : LocalMux
    port map (
            O => \N__37004\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\
        );

    \I__7743\ : CascadeMux
    port map (
            O => \N__37001\,
            I => \N__36998\
        );

    \I__7742\ : InMux
    port map (
            O => \N__36998\,
            I => \N__36995\
        );

    \I__7741\ : LocalMux
    port map (
            O => \N__36995\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\
        );

    \I__7740\ : InMux
    port map (
            O => \N__36992\,
            I => \N__36989\
        );

    \I__7739\ : LocalMux
    port map (
            O => \N__36989\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\
        );

    \I__7738\ : CascadeMux
    port map (
            O => \N__36986\,
            I => \N__36983\
        );

    \I__7737\ : InMux
    port map (
            O => \N__36983\,
            I => \N__36980\
        );

    \I__7736\ : LocalMux
    port map (
            O => \N__36980\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt22\
        );

    \I__7735\ : InMux
    port map (
            O => \N__36977\,
            I => \N__36971\
        );

    \I__7734\ : InMux
    port map (
            O => \N__36976\,
            I => \N__36971\
        );

    \I__7733\ : LocalMux
    port map (
            O => \N__36971\,
            I => \N__36967\
        );

    \I__7732\ : InMux
    port map (
            O => \N__36970\,
            I => \N__36964\
        );

    \I__7731\ : Span4Mux_h
    port map (
            O => \N__36967\,
            I => \N__36961\
        );

    \I__7730\ : LocalMux
    port map (
            O => \N__36964\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__7729\ : Odrv4
    port map (
            O => \N__36961\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__7728\ : CascadeMux
    port map (
            O => \N__36956\,
            I => \N__36953\
        );

    \I__7727\ : InMux
    port map (
            O => \N__36953\,
            I => \N__36947\
        );

    \I__7726\ : InMux
    port map (
            O => \N__36952\,
            I => \N__36947\
        );

    \I__7725\ : LocalMux
    port map (
            O => \N__36947\,
            I => \N__36943\
        );

    \I__7724\ : InMux
    port map (
            O => \N__36946\,
            I => \N__36940\
        );

    \I__7723\ : Span4Mux_v
    port map (
            O => \N__36943\,
            I => \N__36937\
        );

    \I__7722\ : LocalMux
    port map (
            O => \N__36940\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__7721\ : Odrv4
    port map (
            O => \N__36937\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__7720\ : InMux
    port map (
            O => \N__36932\,
            I => \N__36929\
        );

    \I__7719\ : LocalMux
    port map (
            O => \N__36929\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22\
        );

    \I__7718\ : InMux
    port map (
            O => \N__36926\,
            I => \N__36920\
        );

    \I__7717\ : InMux
    port map (
            O => \N__36925\,
            I => \N__36920\
        );

    \I__7716\ : LocalMux
    port map (
            O => \N__36920\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_22\
        );

    \I__7715\ : CascadeMux
    port map (
            O => \N__36917\,
            I => \N__36914\
        );

    \I__7714\ : InMux
    port map (
            O => \N__36914\,
            I => \N__36908\
        );

    \I__7713\ : InMux
    port map (
            O => \N__36913\,
            I => \N__36908\
        );

    \I__7712\ : LocalMux
    port map (
            O => \N__36908\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_23\
        );

    \I__7711\ : CascadeMux
    port map (
            O => \N__36905\,
            I => \N__36902\
        );

    \I__7710\ : InMux
    port map (
            O => \N__36902\,
            I => \N__36899\
        );

    \I__7709\ : LocalMux
    port map (
            O => \N__36899\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\
        );

    \I__7708\ : InMux
    port map (
            O => \N__36896\,
            I => \N__36893\
        );

    \I__7707\ : LocalMux
    port map (
            O => \N__36893\,
            I => \N__36890\
        );

    \I__7706\ : Span4Mux_h
    port map (
            O => \N__36890\,
            I => \N__36885\
        );

    \I__7705\ : InMux
    port map (
            O => \N__36889\,
            I => \N__36880\
        );

    \I__7704\ : InMux
    port map (
            O => \N__36888\,
            I => \N__36880\
        );

    \I__7703\ : Odrv4
    port map (
            O => \N__36885\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5\
        );

    \I__7702\ : LocalMux
    port map (
            O => \N__36880\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5\
        );

    \I__7701\ : InMux
    port map (
            O => \N__36875\,
            I => \N__36872\
        );

    \I__7700\ : LocalMux
    port map (
            O => \N__36872\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\
        );

    \I__7699\ : InMux
    port map (
            O => \N__36869\,
            I => \N__36866\
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__36866\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\
        );

    \I__7697\ : InMux
    port map (
            O => \N__36863\,
            I => \N__36859\
        );

    \I__7696\ : InMux
    port map (
            O => \N__36862\,
            I => \N__36856\
        );

    \I__7695\ : LocalMux
    port map (
            O => \N__36859\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\
        );

    \I__7694\ : LocalMux
    port map (
            O => \N__36856\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\
        );

    \I__7693\ : CascadeMux
    port map (
            O => \N__36851\,
            I => \N__36848\
        );

    \I__7692\ : InMux
    port map (
            O => \N__36848\,
            I => \N__36845\
        );

    \I__7691\ : LocalMux
    port map (
            O => \N__36845\,
            I => \N__36842\
        );

    \I__7690\ : Span4Mux_h
    port map (
            O => \N__36842\,
            I => \N__36839\
        );

    \I__7689\ : Odrv4
    port map (
            O => \N__36839\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt20\
        );

    \I__7688\ : InMux
    port map (
            O => \N__36836\,
            I => \N__36830\
        );

    \I__7687\ : InMux
    port map (
            O => \N__36835\,
            I => \N__36830\
        );

    \I__7686\ : LocalMux
    port map (
            O => \N__36830\,
            I => \N__36826\
        );

    \I__7685\ : InMux
    port map (
            O => \N__36829\,
            I => \N__36823\
        );

    \I__7684\ : Span4Mux_h
    port map (
            O => \N__36826\,
            I => \N__36820\
        );

    \I__7683\ : LocalMux
    port map (
            O => \N__36823\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__7682\ : Odrv4
    port map (
            O => \N__36820\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__7681\ : CascadeMux
    port map (
            O => \N__36815\,
            I => \N__36811\
        );

    \I__7680\ : CascadeMux
    port map (
            O => \N__36814\,
            I => \N__36808\
        );

    \I__7679\ : InMux
    port map (
            O => \N__36811\,
            I => \N__36805\
        );

    \I__7678\ : InMux
    port map (
            O => \N__36808\,
            I => \N__36802\
        );

    \I__7677\ : LocalMux
    port map (
            O => \N__36805\,
            I => \N__36796\
        );

    \I__7676\ : LocalMux
    port map (
            O => \N__36802\,
            I => \N__36796\
        );

    \I__7675\ : InMux
    port map (
            O => \N__36801\,
            I => \N__36793\
        );

    \I__7674\ : Span4Mux_v
    port map (
            O => \N__36796\,
            I => \N__36790\
        );

    \I__7673\ : LocalMux
    port map (
            O => \N__36793\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__7672\ : Odrv4
    port map (
            O => \N__36790\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__7671\ : InMux
    port map (
            O => \N__36785\,
            I => \N__36781\
        );

    \I__7670\ : InMux
    port map (
            O => \N__36784\,
            I => \N__36778\
        );

    \I__7669\ : LocalMux
    port map (
            O => \N__36781\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_21\
        );

    \I__7668\ : LocalMux
    port map (
            O => \N__36778\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_21\
        );

    \I__7667\ : InMux
    port map (
            O => \N__36773\,
            I => \N__36770\
        );

    \I__7666\ : LocalMux
    port map (
            O => \N__36770\,
            I => \N__36767\
        );

    \I__7665\ : Odrv4
    port map (
            O => \N__36767\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20\
        );

    \I__7664\ : InMux
    port map (
            O => \N__36764\,
            I => \bfn_15_21_0_\
        );

    \I__7663\ : InMux
    port map (
            O => \N__36761\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\
        );

    \I__7662\ : InMux
    port map (
            O => \N__36758\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\
        );

    \I__7661\ : InMux
    port map (
            O => \N__36755\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\
        );

    \I__7660\ : InMux
    port map (
            O => \N__36752\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\
        );

    \I__7659\ : IoInMux
    port map (
            O => \N__36749\,
            I => \N__36746\
        );

    \I__7658\ : LocalMux
    port map (
            O => \N__36746\,
            I => \N__36743\
        );

    \I__7657\ : Span4Mux_s3_v
    port map (
            O => \N__36743\,
            I => \N__36740\
        );

    \I__7656\ : Span4Mux_v
    port map (
            O => \N__36740\,
            I => \N__36736\
        );

    \I__7655\ : InMux
    port map (
            O => \N__36739\,
            I => \N__36733\
        );

    \I__7654\ : Odrv4
    port map (
            O => \N__36736\,
            I => \T12_c\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__36733\,
            I => \T12_c\
        );

    \I__7652\ : IoInMux
    port map (
            O => \N__36728\,
            I => \N__36725\
        );

    \I__7651\ : LocalMux
    port map (
            O => \N__36725\,
            I => \N__36722\
        );

    \I__7650\ : Span4Mux_s3_v
    port map (
            O => \N__36722\,
            I => \N__36718\
        );

    \I__7649\ : InMux
    port map (
            O => \N__36721\,
            I => \N__36715\
        );

    \I__7648\ : Odrv4
    port map (
            O => \N__36718\,
            I => \T45_c\
        );

    \I__7647\ : LocalMux
    port map (
            O => \N__36715\,
            I => \T45_c\
        );

    \I__7646\ : InMux
    port map (
            O => \N__36710\,
            I => \N__36704\
        );

    \I__7645\ : InMux
    port map (
            O => \N__36709\,
            I => \N__36704\
        );

    \I__7644\ : LocalMux
    port map (
            O => \N__36704\,
            I => \N__36700\
        );

    \I__7643\ : InMux
    port map (
            O => \N__36703\,
            I => \N__36697\
        );

    \I__7642\ : Span4Mux_h
    port map (
            O => \N__36700\,
            I => \N__36690\
        );

    \I__7641\ : LocalMux
    port map (
            O => \N__36697\,
            I => \N__36687\
        );

    \I__7640\ : InMux
    port map (
            O => \N__36696\,
            I => \N__36684\
        );

    \I__7639\ : InMux
    port map (
            O => \N__36695\,
            I => \N__36679\
        );

    \I__7638\ : InMux
    port map (
            O => \N__36694\,
            I => \N__36679\
        );

    \I__7637\ : InMux
    port map (
            O => \N__36693\,
            I => \N__36675\
        );

    \I__7636\ : Span4Mux_v
    port map (
            O => \N__36690\,
            I => \N__36672\
        );

    \I__7635\ : Span4Mux_v
    port map (
            O => \N__36687\,
            I => \N__36669\
        );

    \I__7634\ : LocalMux
    port map (
            O => \N__36684\,
            I => \N__36664\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__36679\,
            I => \N__36664\
        );

    \I__7632\ : InMux
    port map (
            O => \N__36678\,
            I => \N__36661\
        );

    \I__7631\ : LocalMux
    port map (
            O => \N__36675\,
            I => state_3
        );

    \I__7630\ : Odrv4
    port map (
            O => \N__36672\,
            I => state_3
        );

    \I__7629\ : Odrv4
    port map (
            O => \N__36669\,
            I => state_3
        );

    \I__7628\ : Odrv12
    port map (
            O => \N__36664\,
            I => state_3
        );

    \I__7627\ : LocalMux
    port map (
            O => \N__36661\,
            I => state_3
        );

    \I__7626\ : InMux
    port map (
            O => \N__36650\,
            I => \N__36646\
        );

    \I__7625\ : InMux
    port map (
            O => \N__36649\,
            I => \N__36643\
        );

    \I__7624\ : LocalMux
    port map (
            O => \N__36646\,
            I => \N__36640\
        );

    \I__7623\ : LocalMux
    port map (
            O => \N__36643\,
            I => \N__36637\
        );

    \I__7622\ : Span4Mux_h
    port map (
            O => \N__36640\,
            I => \N__36631\
        );

    \I__7621\ : Span4Mux_h
    port map (
            O => \N__36637\,
            I => \N__36628\
        );

    \I__7620\ : InMux
    port map (
            O => \N__36636\,
            I => \N__36625\
        );

    \I__7619\ : InMux
    port map (
            O => \N__36635\,
            I => \N__36622\
        );

    \I__7618\ : InMux
    port map (
            O => \N__36634\,
            I => \N__36619\
        );

    \I__7617\ : Odrv4
    port map (
            O => \N__36631\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__7616\ : Odrv4
    port map (
            O => \N__36628\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__7615\ : LocalMux
    port map (
            O => \N__36625\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__7614\ : LocalMux
    port map (
            O => \N__36622\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__7613\ : LocalMux
    port map (
            O => \N__36619\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__7612\ : IoInMux
    port map (
            O => \N__36608\,
            I => \N__36605\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__36605\,
            I => \N__36602\
        );

    \I__7610\ : Span4Mux_s2_v
    port map (
            O => \N__36602\,
            I => \N__36599\
        );

    \I__7609\ : Span4Mux_v
    port map (
            O => \N__36599\,
            I => \N__36595\
        );

    \I__7608\ : InMux
    port map (
            O => \N__36598\,
            I => \N__36592\
        );

    \I__7607\ : Odrv4
    port map (
            O => \N__36595\,
            I => \T01_c\
        );

    \I__7606\ : LocalMux
    port map (
            O => \N__36592\,
            I => \T01_c\
        );

    \I__7605\ : InMux
    port map (
            O => \N__36587\,
            I => \N__36583\
        );

    \I__7604\ : InMux
    port map (
            O => \N__36586\,
            I => \N__36580\
        );

    \I__7603\ : LocalMux
    port map (
            O => \N__36583\,
            I => \N__36571\
        );

    \I__7602\ : LocalMux
    port map (
            O => \N__36580\,
            I => \N__36571\
        );

    \I__7601\ : InMux
    port map (
            O => \N__36579\,
            I => \N__36568\
        );

    \I__7600\ : InMux
    port map (
            O => \N__36578\,
            I => \N__36565\
        );

    \I__7599\ : InMux
    port map (
            O => \N__36577\,
            I => \N__36560\
        );

    \I__7598\ : InMux
    port map (
            O => \N__36576\,
            I => \N__36560\
        );

    \I__7597\ : Span4Mux_v
    port map (
            O => \N__36571\,
            I => \N__36555\
        );

    \I__7596\ : LocalMux
    port map (
            O => \N__36568\,
            I => \N__36555\
        );

    \I__7595\ : LocalMux
    port map (
            O => \N__36565\,
            I => \N__36552\
        );

    \I__7594\ : LocalMux
    port map (
            O => \N__36560\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__7593\ : Odrv4
    port map (
            O => \N__36555\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__7592\ : Odrv4
    port map (
            O => \N__36552\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__7591\ : IoInMux
    port map (
            O => \N__36545\,
            I => \N__36542\
        );

    \I__7590\ : LocalMux
    port map (
            O => \N__36542\,
            I => \N__36539\
        );

    \I__7589\ : Span4Mux_s2_v
    port map (
            O => \N__36539\,
            I => \N__36536\
        );

    \I__7588\ : Span4Mux_v
    port map (
            O => \N__36536\,
            I => \N__36532\
        );

    \I__7587\ : InMux
    port map (
            O => \N__36535\,
            I => \N__36529\
        );

    \I__7586\ : Odrv4
    port map (
            O => \N__36532\,
            I => \T23_c\
        );

    \I__7585\ : LocalMux
    port map (
            O => \N__36529\,
            I => \T23_c\
        );

    \I__7584\ : InMux
    port map (
            O => \N__36524\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\
        );

    \I__7583\ : InMux
    port map (
            O => \N__36521\,
            I => \bfn_15_20_0_\
        );

    \I__7582\ : InMux
    port map (
            O => \N__36518\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\
        );

    \I__7581\ : InMux
    port map (
            O => \N__36515\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\
        );

    \I__7580\ : InMux
    port map (
            O => \N__36512\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\
        );

    \I__7579\ : InMux
    port map (
            O => \N__36509\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\
        );

    \I__7578\ : InMux
    port map (
            O => \N__36506\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\
        );

    \I__7577\ : InMux
    port map (
            O => \N__36503\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\
        );

    \I__7576\ : InMux
    port map (
            O => \N__36500\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\
        );

    \I__7575\ : InMux
    port map (
            O => \N__36497\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\
        );

    \I__7574\ : InMux
    port map (
            O => \N__36494\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\
        );

    \I__7573\ : InMux
    port map (
            O => \N__36491\,
            I => \bfn_15_19_0_\
        );

    \I__7572\ : InMux
    port map (
            O => \N__36488\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\
        );

    \I__7571\ : InMux
    port map (
            O => \N__36485\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\
        );

    \I__7570\ : InMux
    port map (
            O => \N__36482\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\
        );

    \I__7569\ : InMux
    port map (
            O => \N__36479\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\
        );

    \I__7568\ : InMux
    port map (
            O => \N__36476\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\
        );

    \I__7567\ : InMux
    port map (
            O => \N__36473\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\
        );

    \I__7566\ : InMux
    port map (
            O => \N__36470\,
            I => \N__36467\
        );

    \I__7565\ : LocalMux
    port map (
            O => \N__36467\,
            I => \N__36464\
        );

    \I__7564\ : Span4Mux_v
    port map (
            O => \N__36464\,
            I => \N__36461\
        );

    \I__7563\ : Odrv4
    port map (
            O => \N__36461\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\
        );

    \I__7562\ : InMux
    port map (
            O => \N__36458\,
            I => \N__36455\
        );

    \I__7561\ : LocalMux
    port map (
            O => \N__36455\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\
        );

    \I__7560\ : InMux
    port map (
            O => \N__36452\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\
        );

    \I__7559\ : InMux
    port map (
            O => \N__36449\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\
        );

    \I__7558\ : InMux
    port map (
            O => \N__36446\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\
        );

    \I__7557\ : InMux
    port map (
            O => \N__36443\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\
        );

    \I__7556\ : InMux
    port map (
            O => \N__36440\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\
        );

    \I__7555\ : CascadeMux
    port map (
            O => \N__36437\,
            I => \N__36434\
        );

    \I__7554\ : InMux
    port map (
            O => \N__36434\,
            I => \N__36431\
        );

    \I__7553\ : LocalMux
    port map (
            O => \N__36431\,
            I => \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0\
        );

    \I__7552\ : InMux
    port map (
            O => \N__36428\,
            I => \N__36425\
        );

    \I__7551\ : LocalMux
    port map (
            O => \N__36425\,
            I => \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0\
        );

    \I__7550\ : CascadeMux
    port map (
            O => \N__36422\,
            I => \N__36419\
        );

    \I__7549\ : InMux
    port map (
            O => \N__36419\,
            I => \N__36416\
        );

    \I__7548\ : LocalMux
    port map (
            O => \N__36416\,
            I => \N__36413\
        );

    \I__7547\ : Odrv4
    port map (
            O => \N__36413\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\
        );

    \I__7546\ : CascadeMux
    port map (
            O => \N__36410\,
            I => \N__36407\
        );

    \I__7545\ : InMux
    port map (
            O => \N__36407\,
            I => \N__36404\
        );

    \I__7544\ : LocalMux
    port map (
            O => \N__36404\,
            I => \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0\
        );

    \I__7543\ : CascadeMux
    port map (
            O => \N__36401\,
            I => \N__36398\
        );

    \I__7542\ : InMux
    port map (
            O => \N__36398\,
            I => \N__36395\
        );

    \I__7541\ : LocalMux
    port map (
            O => \N__36395\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\
        );

    \I__7540\ : InMux
    port map (
            O => \N__36392\,
            I => \N__36389\
        );

    \I__7539\ : LocalMux
    port map (
            O => \N__36389\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\
        );

    \I__7538\ : CascadeMux
    port map (
            O => \N__36386\,
            I => \N__36383\
        );

    \I__7537\ : InMux
    port map (
            O => \N__36383\,
            I => \N__36380\
        );

    \I__7536\ : LocalMux
    port map (
            O => \N__36380\,
            I => \N__36377\
        );

    \I__7535\ : Odrv4
    port map (
            O => \N__36377\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\
        );

    \I__7534\ : CascadeMux
    port map (
            O => \N__36374\,
            I => \N__36371\
        );

    \I__7533\ : InMux
    port map (
            O => \N__36371\,
            I => \N__36368\
        );

    \I__7532\ : LocalMux
    port map (
            O => \N__36368\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\
        );

    \I__7531\ : InMux
    port map (
            O => \N__36365\,
            I => \N__36362\
        );

    \I__7530\ : LocalMux
    port map (
            O => \N__36362\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\
        );

    \I__7529\ : CascadeMux
    port map (
            O => \N__36359\,
            I => \N__36356\
        );

    \I__7528\ : InMux
    port map (
            O => \N__36356\,
            I => \N__36353\
        );

    \I__7527\ : LocalMux
    port map (
            O => \N__36353\,
            I => \N__36350\
        );

    \I__7526\ : Span4Mux_h
    port map (
            O => \N__36350\,
            I => \N__36347\
        );

    \I__7525\ : Odrv4
    port map (
            O => \N__36347\,
            I => \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\
        );

    \I__7524\ : InMux
    port map (
            O => \N__36344\,
            I => \N__36341\
        );

    \I__7523\ : LocalMux
    port map (
            O => \N__36341\,
            I => \N__36338\
        );

    \I__7522\ : Odrv4
    port map (
            O => \N__36338\,
            I => \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0\
        );

    \I__7521\ : CascadeMux
    port map (
            O => \N__36335\,
            I => \N__36332\
        );

    \I__7520\ : InMux
    port map (
            O => \N__36332\,
            I => \N__36329\
        );

    \I__7519\ : LocalMux
    port map (
            O => \N__36329\,
            I => \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0\
        );

    \I__7518\ : InMux
    port map (
            O => \N__36326\,
            I => \N__36323\
        );

    \I__7517\ : LocalMux
    port map (
            O => \N__36323\,
            I => \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0\
        );

    \I__7516\ : InMux
    port map (
            O => \N__36320\,
            I => \N__36317\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__36317\,
            I => \N__36314\
        );

    \I__7514\ : Odrv4
    port map (
            O => \N__36314\,
            I => \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0\
        );

    \I__7513\ : CascadeMux
    port map (
            O => \N__36311\,
            I => \N__36308\
        );

    \I__7512\ : InMux
    port map (
            O => \N__36308\,
            I => \N__36305\
        );

    \I__7511\ : LocalMux
    port map (
            O => \N__36305\,
            I => \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0\
        );

    \I__7510\ : InMux
    port map (
            O => \N__36302\,
            I => \N__36299\
        );

    \I__7509\ : LocalMux
    port map (
            O => \N__36299\,
            I => \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0\
        );

    \I__7508\ : CascadeMux
    port map (
            O => \N__36296\,
            I => \N__36293\
        );

    \I__7507\ : InMux
    port map (
            O => \N__36293\,
            I => \N__36290\
        );

    \I__7506\ : LocalMux
    port map (
            O => \N__36290\,
            I => \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0\
        );

    \I__7505\ : CascadeMux
    port map (
            O => \N__36287\,
            I => \N__36283\
        );

    \I__7504\ : InMux
    port map (
            O => \N__36286\,
            I => \N__36280\
        );

    \I__7503\ : InMux
    port map (
            O => \N__36283\,
            I => \N__36276\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__36280\,
            I => \N__36273\
        );

    \I__7501\ : InMux
    port map (
            O => \N__36279\,
            I => \N__36270\
        );

    \I__7500\ : LocalMux
    port map (
            O => \N__36276\,
            I => \N__36267\
        );

    \I__7499\ : Span4Mux_v
    port map (
            O => \N__36273\,
            I => \N__36264\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__36270\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__7497\ : Odrv4
    port map (
            O => \N__36267\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__7496\ : Odrv4
    port map (
            O => \N__36264\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__7495\ : InMux
    port map (
            O => \N__36257\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__7494\ : InMux
    port map (
            O => \N__36254\,
            I => \N__36250\
        );

    \I__7493\ : InMux
    port map (
            O => \N__36253\,
            I => \N__36247\
        );

    \I__7492\ : LocalMux
    port map (
            O => \N__36250\,
            I => \N__36244\
        );

    \I__7491\ : LocalMux
    port map (
            O => \N__36247\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__7490\ : Odrv12
    port map (
            O => \N__36244\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__7489\ : CascadeMux
    port map (
            O => \N__36239\,
            I => \N__36236\
        );

    \I__7488\ : InMux
    port map (
            O => \N__36236\,
            I => \N__36231\
        );

    \I__7487\ : InMux
    port map (
            O => \N__36235\,
            I => \N__36228\
        );

    \I__7486\ : InMux
    port map (
            O => \N__36234\,
            I => \N__36225\
        );

    \I__7485\ : LocalMux
    port map (
            O => \N__36231\,
            I => \N__36218\
        );

    \I__7484\ : LocalMux
    port map (
            O => \N__36228\,
            I => \N__36218\
        );

    \I__7483\ : LocalMux
    port map (
            O => \N__36225\,
            I => \N__36218\
        );

    \I__7482\ : Odrv4
    port map (
            O => \N__36218\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__7481\ : InMux
    port map (
            O => \N__36215\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__7480\ : InMux
    port map (
            O => \N__36212\,
            I => \N__36208\
        );

    \I__7479\ : InMux
    port map (
            O => \N__36211\,
            I => \N__36205\
        );

    \I__7478\ : LocalMux
    port map (
            O => \N__36208\,
            I => \N__36202\
        );

    \I__7477\ : LocalMux
    port map (
            O => \N__36205\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__7476\ : Odrv12
    port map (
            O => \N__36202\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__7475\ : CascadeMux
    port map (
            O => \N__36197\,
            I => \N__36194\
        );

    \I__7474\ : InMux
    port map (
            O => \N__36194\,
            I => \N__36189\
        );

    \I__7473\ : InMux
    port map (
            O => \N__36193\,
            I => \N__36186\
        );

    \I__7472\ : InMux
    port map (
            O => \N__36192\,
            I => \N__36183\
        );

    \I__7471\ : LocalMux
    port map (
            O => \N__36189\,
            I => \N__36178\
        );

    \I__7470\ : LocalMux
    port map (
            O => \N__36186\,
            I => \N__36178\
        );

    \I__7469\ : LocalMux
    port map (
            O => \N__36183\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__7468\ : Odrv4
    port map (
            O => \N__36178\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__7467\ : InMux
    port map (
            O => \N__36173\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__7466\ : InMux
    port map (
            O => \N__36170\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__7465\ : CEMux
    port map (
            O => \N__36167\,
            I => \N__36163\
        );

    \I__7464\ : CEMux
    port map (
            O => \N__36166\,
            I => \N__36160\
        );

    \I__7463\ : LocalMux
    port map (
            O => \N__36163\,
            I => \N__36154\
        );

    \I__7462\ : LocalMux
    port map (
            O => \N__36160\,
            I => \N__36151\
        );

    \I__7461\ : CEMux
    port map (
            O => \N__36159\,
            I => \N__36148\
        );

    \I__7460\ : CEMux
    port map (
            O => \N__36158\,
            I => \N__36145\
        );

    \I__7459\ : CEMux
    port map (
            O => \N__36157\,
            I => \N__36142\
        );

    \I__7458\ : Span4Mux_v
    port map (
            O => \N__36154\,
            I => \N__36139\
        );

    \I__7457\ : Span4Mux_v
    port map (
            O => \N__36151\,
            I => \N__36136\
        );

    \I__7456\ : LocalMux
    port map (
            O => \N__36148\,
            I => \N__36133\
        );

    \I__7455\ : LocalMux
    port map (
            O => \N__36145\,
            I => \N__36130\
        );

    \I__7454\ : LocalMux
    port map (
            O => \N__36142\,
            I => \N__36127\
        );

    \I__7453\ : Span4Mux_h
    port map (
            O => \N__36139\,
            I => \N__36124\
        );

    \I__7452\ : Span4Mux_h
    port map (
            O => \N__36136\,
            I => \N__36119\
        );

    \I__7451\ : Span4Mux_h
    port map (
            O => \N__36133\,
            I => \N__36119\
        );

    \I__7450\ : Span4Mux_v
    port map (
            O => \N__36130\,
            I => \N__36116\
        );

    \I__7449\ : Span4Mux_h
    port map (
            O => \N__36127\,
            I => \N__36113\
        );

    \I__7448\ : Span4Mux_v
    port map (
            O => \N__36124\,
            I => \N__36108\
        );

    \I__7447\ : Span4Mux_h
    port map (
            O => \N__36119\,
            I => \N__36108\
        );

    \I__7446\ : Span4Mux_h
    port map (
            O => \N__36116\,
            I => \N__36103\
        );

    \I__7445\ : Span4Mux_h
    port map (
            O => \N__36113\,
            I => \N__36103\
        );

    \I__7444\ : Odrv4
    port map (
            O => \N__36108\,
            I => \delay_measurement_inst.delay_tr_timer.N_204_i\
        );

    \I__7443\ : Odrv4
    port map (
            O => \N__36103\,
            I => \delay_measurement_inst.delay_tr_timer.N_204_i\
        );

    \I__7442\ : InMux
    port map (
            O => \N__36098\,
            I => \N__36095\
        );

    \I__7441\ : LocalMux
    port map (
            O => \N__36095\,
            I => \N__36092\
        );

    \I__7440\ : Span4Mux_h
    port map (
            O => \N__36092\,
            I => \N__36089\
        );

    \I__7439\ : Odrv4
    port map (
            O => \N__36089\,
            I => \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\
        );

    \I__7438\ : CascadeMux
    port map (
            O => \N__36086\,
            I => \N__36083\
        );

    \I__7437\ : InMux
    port map (
            O => \N__36083\,
            I => \N__36080\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__36080\,
            I => \N__36077\
        );

    \I__7435\ : Odrv4
    port map (
            O => \N__36077\,
            I => \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\
        );

    \I__7434\ : InMux
    port map (
            O => \N__36074\,
            I => \N__36071\
        );

    \I__7433\ : LocalMux
    port map (
            O => \N__36071\,
            I => \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\
        );

    \I__7432\ : CascadeMux
    port map (
            O => \N__36068\,
            I => \N__36065\
        );

    \I__7431\ : InMux
    port map (
            O => \N__36065\,
            I => \N__36062\
        );

    \I__7430\ : LocalMux
    port map (
            O => \N__36062\,
            I => \N__36059\
        );

    \I__7429\ : Span4Mux_v
    port map (
            O => \N__36059\,
            I => \N__36056\
        );

    \I__7428\ : Odrv4
    port map (
            O => \N__36056\,
            I => \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0\
        );

    \I__7427\ : InMux
    port map (
            O => \N__36053\,
            I => \N__36050\
        );

    \I__7426\ : LocalMux
    port map (
            O => \N__36050\,
            I => \N__36047\
        );

    \I__7425\ : Sp12to4
    port map (
            O => \N__36047\,
            I => \N__36044\
        );

    \I__7424\ : Odrv12
    port map (
            O => \N__36044\,
            I => \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0\
        );

    \I__7423\ : CascadeMux
    port map (
            O => \N__36041\,
            I => \N__36037\
        );

    \I__7422\ : CascadeMux
    port map (
            O => \N__36040\,
            I => \N__36034\
        );

    \I__7421\ : InMux
    port map (
            O => \N__36037\,
            I => \N__36031\
        );

    \I__7420\ : InMux
    port map (
            O => \N__36034\,
            I => \N__36027\
        );

    \I__7419\ : LocalMux
    port map (
            O => \N__36031\,
            I => \N__36024\
        );

    \I__7418\ : InMux
    port map (
            O => \N__36030\,
            I => \N__36021\
        );

    \I__7417\ : LocalMux
    port map (
            O => \N__36027\,
            I => \N__36018\
        );

    \I__7416\ : Span4Mux_v
    port map (
            O => \N__36024\,
            I => \N__36015\
        );

    \I__7415\ : LocalMux
    port map (
            O => \N__36021\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__7414\ : Odrv4
    port map (
            O => \N__36018\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__7413\ : Odrv4
    port map (
            O => \N__36015\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__7412\ : InMux
    port map (
            O => \N__36008\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__7411\ : CascadeMux
    port map (
            O => \N__36005\,
            I => \N__36002\
        );

    \I__7410\ : InMux
    port map (
            O => \N__36002\,
            I => \N__35997\
        );

    \I__7409\ : InMux
    port map (
            O => \N__36001\,
            I => \N__35994\
        );

    \I__7408\ : InMux
    port map (
            O => \N__36000\,
            I => \N__35991\
        );

    \I__7407\ : LocalMux
    port map (
            O => \N__35997\,
            I => \N__35984\
        );

    \I__7406\ : LocalMux
    port map (
            O => \N__35994\,
            I => \N__35984\
        );

    \I__7405\ : LocalMux
    port map (
            O => \N__35991\,
            I => \N__35984\
        );

    \I__7404\ : Odrv4
    port map (
            O => \N__35984\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__7403\ : InMux
    port map (
            O => \N__35981\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__7402\ : InMux
    port map (
            O => \N__35978\,
            I => \N__35971\
        );

    \I__7401\ : InMux
    port map (
            O => \N__35977\,
            I => \N__35971\
        );

    \I__7400\ : InMux
    port map (
            O => \N__35976\,
            I => \N__35968\
        );

    \I__7399\ : LocalMux
    port map (
            O => \N__35971\,
            I => \N__35965\
        );

    \I__7398\ : LocalMux
    port map (
            O => \N__35968\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__7397\ : Odrv4
    port map (
            O => \N__35965\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__7396\ : InMux
    port map (
            O => \N__35960\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__7395\ : InMux
    port map (
            O => \N__35957\,
            I => \N__35950\
        );

    \I__7394\ : InMux
    port map (
            O => \N__35956\,
            I => \N__35950\
        );

    \I__7393\ : InMux
    port map (
            O => \N__35955\,
            I => \N__35947\
        );

    \I__7392\ : LocalMux
    port map (
            O => \N__35950\,
            I => \N__35944\
        );

    \I__7391\ : LocalMux
    port map (
            O => \N__35947\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__7390\ : Odrv4
    port map (
            O => \N__35944\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__7389\ : InMux
    port map (
            O => \N__35939\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__7388\ : CascadeMux
    port map (
            O => \N__35936\,
            I => \N__35932\
        );

    \I__7387\ : InMux
    port map (
            O => \N__35935\,
            I => \N__35928\
        );

    \I__7386\ : InMux
    port map (
            O => \N__35932\,
            I => \N__35925\
        );

    \I__7385\ : InMux
    port map (
            O => \N__35931\,
            I => \N__35922\
        );

    \I__7384\ : LocalMux
    port map (
            O => \N__35928\,
            I => \N__35917\
        );

    \I__7383\ : LocalMux
    port map (
            O => \N__35925\,
            I => \N__35917\
        );

    \I__7382\ : LocalMux
    port map (
            O => \N__35922\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__7381\ : Odrv12
    port map (
            O => \N__35917\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__7380\ : InMux
    port map (
            O => \N__35912\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__7379\ : CascadeMux
    port map (
            O => \N__35909\,
            I => \N__35905\
        );

    \I__7378\ : CascadeMux
    port map (
            O => \N__35908\,
            I => \N__35902\
        );

    \I__7377\ : InMux
    port map (
            O => \N__35905\,
            I => \N__35896\
        );

    \I__7376\ : InMux
    port map (
            O => \N__35902\,
            I => \N__35896\
        );

    \I__7375\ : InMux
    port map (
            O => \N__35901\,
            I => \N__35893\
        );

    \I__7374\ : LocalMux
    port map (
            O => \N__35896\,
            I => \N__35890\
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__35893\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__7372\ : Odrv12
    port map (
            O => \N__35890\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__7371\ : InMux
    port map (
            O => \N__35885\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__7370\ : CascadeMux
    port map (
            O => \N__35882\,
            I => \N__35878\
        );

    \I__7369\ : CascadeMux
    port map (
            O => \N__35881\,
            I => \N__35875\
        );

    \I__7368\ : InMux
    port map (
            O => \N__35878\,
            I => \N__35869\
        );

    \I__7367\ : InMux
    port map (
            O => \N__35875\,
            I => \N__35869\
        );

    \I__7366\ : InMux
    port map (
            O => \N__35874\,
            I => \N__35866\
        );

    \I__7365\ : LocalMux
    port map (
            O => \N__35869\,
            I => \N__35863\
        );

    \I__7364\ : LocalMux
    port map (
            O => \N__35866\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__7363\ : Odrv4
    port map (
            O => \N__35863\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__7362\ : InMux
    port map (
            O => \N__35858\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__7361\ : CascadeMux
    port map (
            O => \N__35855\,
            I => \N__35852\
        );

    \I__7360\ : InMux
    port map (
            O => \N__35852\,
            I => \N__35848\
        );

    \I__7359\ : InMux
    port map (
            O => \N__35851\,
            I => \N__35845\
        );

    \I__7358\ : LocalMux
    port map (
            O => \N__35848\,
            I => \N__35839\
        );

    \I__7357\ : LocalMux
    port map (
            O => \N__35845\,
            I => \N__35839\
        );

    \I__7356\ : InMux
    port map (
            O => \N__35844\,
            I => \N__35836\
        );

    \I__7355\ : Span4Mux_v
    port map (
            O => \N__35839\,
            I => \N__35833\
        );

    \I__7354\ : LocalMux
    port map (
            O => \N__35836\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__7353\ : Odrv4
    port map (
            O => \N__35833\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__7352\ : InMux
    port map (
            O => \N__35828\,
            I => \bfn_15_13_0_\
        );

    \I__7351\ : CascadeMux
    port map (
            O => \N__35825\,
            I => \N__35820\
        );

    \I__7350\ : InMux
    port map (
            O => \N__35824\,
            I => \N__35817\
        );

    \I__7349\ : InMux
    port map (
            O => \N__35823\,
            I => \N__35814\
        );

    \I__7348\ : InMux
    port map (
            O => \N__35820\,
            I => \N__35811\
        );

    \I__7347\ : LocalMux
    port map (
            O => \N__35817\,
            I => \N__35808\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__35814\,
            I => \N__35801\
        );

    \I__7345\ : LocalMux
    port map (
            O => \N__35811\,
            I => \N__35801\
        );

    \I__7344\ : Span4Mux_v
    port map (
            O => \N__35808\,
            I => \N__35801\
        );

    \I__7343\ : Odrv4
    port map (
            O => \N__35801\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__7342\ : InMux
    port map (
            O => \N__35798\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__7341\ : InMux
    port map (
            O => \N__35795\,
            I => \N__35788\
        );

    \I__7340\ : InMux
    port map (
            O => \N__35794\,
            I => \N__35788\
        );

    \I__7339\ : InMux
    port map (
            O => \N__35793\,
            I => \N__35785\
        );

    \I__7338\ : LocalMux
    port map (
            O => \N__35788\,
            I => \N__35782\
        );

    \I__7337\ : LocalMux
    port map (
            O => \N__35785\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__7336\ : Odrv4
    port map (
            O => \N__35782\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__7335\ : InMux
    port map (
            O => \N__35777\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__7334\ : CascadeMux
    port map (
            O => \N__35774\,
            I => \N__35771\
        );

    \I__7333\ : InMux
    port map (
            O => \N__35771\,
            I => \N__35766\
        );

    \I__7332\ : InMux
    port map (
            O => \N__35770\,
            I => \N__35763\
        );

    \I__7331\ : InMux
    port map (
            O => \N__35769\,
            I => \N__35760\
        );

    \I__7330\ : LocalMux
    port map (
            O => \N__35766\,
            I => \N__35755\
        );

    \I__7329\ : LocalMux
    port map (
            O => \N__35763\,
            I => \N__35755\
        );

    \I__7328\ : LocalMux
    port map (
            O => \N__35760\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__7327\ : Odrv12
    port map (
            O => \N__35755\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__7326\ : InMux
    port map (
            O => \N__35750\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__7325\ : CascadeMux
    port map (
            O => \N__35747\,
            I => \N__35743\
        );

    \I__7324\ : CascadeMux
    port map (
            O => \N__35746\,
            I => \N__35740\
        );

    \I__7323\ : InMux
    port map (
            O => \N__35743\,
            I => \N__35734\
        );

    \I__7322\ : InMux
    port map (
            O => \N__35740\,
            I => \N__35734\
        );

    \I__7321\ : InMux
    port map (
            O => \N__35739\,
            I => \N__35731\
        );

    \I__7320\ : LocalMux
    port map (
            O => \N__35734\,
            I => \N__35728\
        );

    \I__7319\ : LocalMux
    port map (
            O => \N__35731\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__7318\ : Odrv12
    port map (
            O => \N__35728\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__7317\ : InMux
    port map (
            O => \N__35723\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__7316\ : CascadeMux
    port map (
            O => \N__35720\,
            I => \N__35717\
        );

    \I__7315\ : InMux
    port map (
            O => \N__35717\,
            I => \N__35712\
        );

    \I__7314\ : InMux
    port map (
            O => \N__35716\,
            I => \N__35709\
        );

    \I__7313\ : InMux
    port map (
            O => \N__35715\,
            I => \N__35706\
        );

    \I__7312\ : LocalMux
    port map (
            O => \N__35712\,
            I => \N__35701\
        );

    \I__7311\ : LocalMux
    port map (
            O => \N__35709\,
            I => \N__35701\
        );

    \I__7310\ : LocalMux
    port map (
            O => \N__35706\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__7309\ : Odrv12
    port map (
            O => \N__35701\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__7308\ : InMux
    port map (
            O => \N__35696\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__7307\ : CascadeMux
    port map (
            O => \N__35693\,
            I => \N__35690\
        );

    \I__7306\ : InMux
    port map (
            O => \N__35690\,
            I => \N__35685\
        );

    \I__7305\ : InMux
    port map (
            O => \N__35689\,
            I => \N__35682\
        );

    \I__7304\ : InMux
    port map (
            O => \N__35688\,
            I => \N__35679\
        );

    \I__7303\ : LocalMux
    port map (
            O => \N__35685\,
            I => \N__35674\
        );

    \I__7302\ : LocalMux
    port map (
            O => \N__35682\,
            I => \N__35674\
        );

    \I__7301\ : LocalMux
    port map (
            O => \N__35679\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__7300\ : Odrv12
    port map (
            O => \N__35674\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__7299\ : InMux
    port map (
            O => \N__35669\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__7298\ : InMux
    port map (
            O => \N__35666\,
            I => \N__35661\
        );

    \I__7297\ : InMux
    port map (
            O => \N__35665\,
            I => \N__35656\
        );

    \I__7296\ : InMux
    port map (
            O => \N__35664\,
            I => \N__35656\
        );

    \I__7295\ : LocalMux
    port map (
            O => \N__35661\,
            I => \N__35651\
        );

    \I__7294\ : LocalMux
    port map (
            O => \N__35656\,
            I => \N__35651\
        );

    \I__7293\ : Odrv4
    port map (
            O => \N__35651\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__7292\ : InMux
    port map (
            O => \N__35648\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__7291\ : CascadeMux
    port map (
            O => \N__35645\,
            I => \N__35641\
        );

    \I__7290\ : InMux
    port map (
            O => \N__35644\,
            I => \N__35638\
        );

    \I__7289\ : InMux
    port map (
            O => \N__35641\,
            I => \N__35634\
        );

    \I__7288\ : LocalMux
    port map (
            O => \N__35638\,
            I => \N__35631\
        );

    \I__7287\ : InMux
    port map (
            O => \N__35637\,
            I => \N__35628\
        );

    \I__7286\ : LocalMux
    port map (
            O => \N__35634\,
            I => \N__35623\
        );

    \I__7285\ : Span4Mux_v
    port map (
            O => \N__35631\,
            I => \N__35623\
        );

    \I__7284\ : LocalMux
    port map (
            O => \N__35628\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__7283\ : Odrv4
    port map (
            O => \N__35623\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__7282\ : InMux
    port map (
            O => \N__35618\,
            I => \bfn_15_12_0_\
        );

    \I__7281\ : InMux
    port map (
            O => \N__35615\,
            I => \N__35612\
        );

    \I__7280\ : LocalMux
    port map (
            O => \N__35612\,
            I => \N__35608\
        );

    \I__7279\ : InMux
    port map (
            O => \N__35611\,
            I => \N__35605\
        );

    \I__7278\ : Span4Mux_h
    port map (
            O => \N__35608\,
            I => \N__35601\
        );

    \I__7277\ : LocalMux
    port map (
            O => \N__35605\,
            I => \N__35598\
        );

    \I__7276\ : InMux
    port map (
            O => \N__35604\,
            I => \N__35595\
        );

    \I__7275\ : Odrv4
    port map (
            O => \N__35601\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__7274\ : Odrv4
    port map (
            O => \N__35598\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__7273\ : LocalMux
    port map (
            O => \N__35595\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__7272\ : InMux
    port map (
            O => \N__35588\,
            I => \N__35584\
        );

    \I__7271\ : CascadeMux
    port map (
            O => \N__35587\,
            I => \N__35581\
        );

    \I__7270\ : LocalMux
    port map (
            O => \N__35584\,
            I => \N__35578\
        );

    \I__7269\ : InMux
    port map (
            O => \N__35581\,
            I => \N__35574\
        );

    \I__7268\ : Span4Mux_h
    port map (
            O => \N__35578\,
            I => \N__35571\
        );

    \I__7267\ : InMux
    port map (
            O => \N__35577\,
            I => \N__35568\
        );

    \I__7266\ : LocalMux
    port map (
            O => \N__35574\,
            I => \N__35565\
        );

    \I__7265\ : Odrv4
    port map (
            O => \N__35571\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__7264\ : LocalMux
    port map (
            O => \N__35568\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__7263\ : Odrv12
    port map (
            O => \N__35565\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__7262\ : InMux
    port map (
            O => \N__35558\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__7261\ : CascadeMux
    port map (
            O => \N__35555\,
            I => \N__35551\
        );

    \I__7260\ : CascadeMux
    port map (
            O => \N__35554\,
            I => \N__35548\
        );

    \I__7259\ : InMux
    port map (
            O => \N__35551\,
            I => \N__35542\
        );

    \I__7258\ : InMux
    port map (
            O => \N__35548\,
            I => \N__35542\
        );

    \I__7257\ : InMux
    port map (
            O => \N__35547\,
            I => \N__35539\
        );

    \I__7256\ : LocalMux
    port map (
            O => \N__35542\,
            I => \N__35536\
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__35539\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__7254\ : Odrv12
    port map (
            O => \N__35536\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__7253\ : InMux
    port map (
            O => \N__35531\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__7252\ : InMux
    port map (
            O => \N__35528\,
            I => \N__35521\
        );

    \I__7251\ : InMux
    port map (
            O => \N__35527\,
            I => \N__35521\
        );

    \I__7250\ : InMux
    port map (
            O => \N__35526\,
            I => \N__35518\
        );

    \I__7249\ : LocalMux
    port map (
            O => \N__35521\,
            I => \N__35515\
        );

    \I__7248\ : LocalMux
    port map (
            O => \N__35518\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__7247\ : Odrv4
    port map (
            O => \N__35515\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__7246\ : InMux
    port map (
            O => \N__35510\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__7245\ : CascadeMux
    port map (
            O => \N__35507\,
            I => \N__35504\
        );

    \I__7244\ : InMux
    port map (
            O => \N__35504\,
            I => \N__35499\
        );

    \I__7243\ : InMux
    port map (
            O => \N__35503\,
            I => \N__35496\
        );

    \I__7242\ : InMux
    port map (
            O => \N__35502\,
            I => \N__35493\
        );

    \I__7241\ : LocalMux
    port map (
            O => \N__35499\,
            I => \N__35488\
        );

    \I__7240\ : LocalMux
    port map (
            O => \N__35496\,
            I => \N__35488\
        );

    \I__7239\ : LocalMux
    port map (
            O => \N__35493\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__7238\ : Odrv12
    port map (
            O => \N__35488\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__7237\ : InMux
    port map (
            O => \N__35483\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__7236\ : CascadeMux
    port map (
            O => \N__35480\,
            I => \N__35476\
        );

    \I__7235\ : CascadeMux
    port map (
            O => \N__35479\,
            I => \N__35473\
        );

    \I__7234\ : InMux
    port map (
            O => \N__35476\,
            I => \N__35467\
        );

    \I__7233\ : InMux
    port map (
            O => \N__35473\,
            I => \N__35467\
        );

    \I__7232\ : InMux
    port map (
            O => \N__35472\,
            I => \N__35464\
        );

    \I__7231\ : LocalMux
    port map (
            O => \N__35467\,
            I => \N__35461\
        );

    \I__7230\ : LocalMux
    port map (
            O => \N__35464\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__7229\ : Odrv4
    port map (
            O => \N__35461\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__7228\ : InMux
    port map (
            O => \N__35456\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__7227\ : InMux
    port map (
            O => \N__35453\,
            I => \N__35448\
        );

    \I__7226\ : InMux
    port map (
            O => \N__35452\,
            I => \N__35443\
        );

    \I__7225\ : InMux
    port map (
            O => \N__35451\,
            I => \N__35443\
        );

    \I__7224\ : LocalMux
    port map (
            O => \N__35448\,
            I => \N__35438\
        );

    \I__7223\ : LocalMux
    port map (
            O => \N__35443\,
            I => \N__35438\
        );

    \I__7222\ : Odrv4
    port map (
            O => \N__35438\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__7221\ : InMux
    port map (
            O => \N__35435\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__7220\ : CascadeMux
    port map (
            O => \N__35432\,
            I => \N__35429\
        );

    \I__7219\ : InMux
    port map (
            O => \N__35429\,
            I => \N__35424\
        );

    \I__7218\ : InMux
    port map (
            O => \N__35428\,
            I => \N__35421\
        );

    \I__7217\ : InMux
    port map (
            O => \N__35427\,
            I => \N__35418\
        );

    \I__7216\ : LocalMux
    port map (
            O => \N__35424\,
            I => \N__35413\
        );

    \I__7215\ : LocalMux
    port map (
            O => \N__35421\,
            I => \N__35413\
        );

    \I__7214\ : LocalMux
    port map (
            O => \N__35418\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__7213\ : Odrv12
    port map (
            O => \N__35413\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__7212\ : InMux
    port map (
            O => \N__35408\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__7211\ : CascadeMux
    port map (
            O => \N__35405\,
            I => \N__35401\
        );

    \I__7210\ : CascadeMux
    port map (
            O => \N__35404\,
            I => \N__35398\
        );

    \I__7209\ : InMux
    port map (
            O => \N__35401\,
            I => \N__35395\
        );

    \I__7208\ : InMux
    port map (
            O => \N__35398\,
            I => \N__35391\
        );

    \I__7207\ : LocalMux
    port map (
            O => \N__35395\,
            I => \N__35388\
        );

    \I__7206\ : InMux
    port map (
            O => \N__35394\,
            I => \N__35385\
        );

    \I__7205\ : LocalMux
    port map (
            O => \N__35391\,
            I => \N__35382\
        );

    \I__7204\ : Span4Mux_v
    port map (
            O => \N__35388\,
            I => \N__35379\
        );

    \I__7203\ : LocalMux
    port map (
            O => \N__35385\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__7202\ : Odrv4
    port map (
            O => \N__35382\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__7201\ : Odrv4
    port map (
            O => \N__35379\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__7200\ : InMux
    port map (
            O => \N__35372\,
            I => \bfn_15_11_0_\
        );

    \I__7199\ : InMux
    port map (
            O => \N__35369\,
            I => \N__35366\
        );

    \I__7198\ : LocalMux
    port map (
            O => \N__35366\,
            I => \N__35363\
        );

    \I__7197\ : Odrv4
    port map (
            O => \N__35363\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\
        );

    \I__7196\ : CascadeMux
    port map (
            O => \N__35360\,
            I => \N__35357\
        );

    \I__7195\ : InMux
    port map (
            O => \N__35357\,
            I => \N__35354\
        );

    \I__7194\ : LocalMux
    port map (
            O => \N__35354\,
            I => \N__35351\
        );

    \I__7193\ : Span4Mux_v
    port map (
            O => \N__35351\,
            I => \N__35348\
        );

    \I__7192\ : Odrv4
    port map (
            O => \N__35348\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt18\
        );

    \I__7191\ : InMux
    port map (
            O => \N__35345\,
            I => \N__35342\
        );

    \I__7190\ : LocalMux
    port map (
            O => \N__35342\,
            I => \N__35339\
        );

    \I__7189\ : Odrv4
    port map (
            O => \N__35339\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\
        );

    \I__7188\ : CascadeMux
    port map (
            O => \N__35336\,
            I => \N__35333\
        );

    \I__7187\ : InMux
    port map (
            O => \N__35333\,
            I => \N__35329\
        );

    \I__7186\ : InMux
    port map (
            O => \N__35332\,
            I => \N__35326\
        );

    \I__7185\ : LocalMux
    port map (
            O => \N__35329\,
            I => \N__35323\
        );

    \I__7184\ : LocalMux
    port map (
            O => \N__35326\,
            I => \N__35320\
        );

    \I__7183\ : Odrv4
    port map (
            O => \N__35323\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt30\
        );

    \I__7182\ : Odrv4
    port map (
            O => \N__35320\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt30\
        );

    \I__7181\ : InMux
    port map (
            O => \N__35315\,
            I => \N__35312\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__35312\,
            I => \N__35309\
        );

    \I__7179\ : Span4Mux_h
    port map (
            O => \N__35309\,
            I => \N__35306\
        );

    \I__7178\ : Odrv4
    port map (
            O => \N__35306\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO\
        );

    \I__7177\ : InMux
    port map (
            O => \N__35303\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_28\
        );

    \I__7176\ : InMux
    port map (
            O => \N__35300\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_30\
        );

    \I__7175\ : InMux
    port map (
            O => \N__35297\,
            I => \N__35293\
        );

    \I__7174\ : InMux
    port map (
            O => \N__35296\,
            I => \N__35290\
        );

    \I__7173\ : LocalMux
    port map (
            O => \N__35293\,
            I => \N__35287\
        );

    \I__7172\ : LocalMux
    port map (
            O => \N__35290\,
            I => \N__35284\
        );

    \I__7171\ : Span4Mux_h
    port map (
            O => \N__35287\,
            I => \N__35281\
        );

    \I__7170\ : Span4Mux_h
    port map (
            O => \N__35284\,
            I => \N__35278\
        );

    \I__7169\ : Odrv4
    port map (
            O => \N__35281\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__7168\ : Odrv4
    port map (
            O => \N__35278\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__7167\ : InMux
    port map (
            O => \N__35273\,
            I => \N__35269\
        );

    \I__7166\ : InMux
    port map (
            O => \N__35272\,
            I => \N__35266\
        );

    \I__7165\ : LocalMux
    port map (
            O => \N__35269\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__7164\ : LocalMux
    port map (
            O => \N__35266\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__7163\ : InMux
    port map (
            O => \N__35261\,
            I => \N__35258\
        );

    \I__7162\ : LocalMux
    port map (
            O => \N__35258\,
            I => \N__35255\
        );

    \I__7161\ : Odrv4
    port map (
            O => \N__35255\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\
        );

    \I__7160\ : InMux
    port map (
            O => \N__35252\,
            I => \N__35248\
        );

    \I__7159\ : InMux
    port map (
            O => \N__35251\,
            I => \N__35245\
        );

    \I__7158\ : LocalMux
    port map (
            O => \N__35248\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__35245\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__7156\ : CascadeMux
    port map (
            O => \N__35240\,
            I => \N__35237\
        );

    \I__7155\ : InMux
    port map (
            O => \N__35237\,
            I => \N__35234\
        );

    \I__7154\ : LocalMux
    port map (
            O => \N__35234\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\
        );

    \I__7153\ : InMux
    port map (
            O => \N__35231\,
            I => \N__35227\
        );

    \I__7152\ : InMux
    port map (
            O => \N__35230\,
            I => \N__35224\
        );

    \I__7151\ : LocalMux
    port map (
            O => \N__35227\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__7150\ : LocalMux
    port map (
            O => \N__35224\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__7149\ : InMux
    port map (
            O => \N__35219\,
            I => \N__35216\
        );

    \I__7148\ : LocalMux
    port map (
            O => \N__35216\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\
        );

    \I__7147\ : InMux
    port map (
            O => \N__35213\,
            I => \N__35209\
        );

    \I__7146\ : InMux
    port map (
            O => \N__35212\,
            I => \N__35206\
        );

    \I__7145\ : LocalMux
    port map (
            O => \N__35209\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__7144\ : LocalMux
    port map (
            O => \N__35206\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__7143\ : InMux
    port map (
            O => \N__35201\,
            I => \N__35198\
        );

    \I__7142\ : LocalMux
    port map (
            O => \N__35198\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\
        );

    \I__7141\ : InMux
    port map (
            O => \N__35195\,
            I => \N__35192\
        );

    \I__7140\ : LocalMux
    port map (
            O => \N__35192\,
            I => \N__35189\
        );

    \I__7139\ : Span4Mux_h
    port map (
            O => \N__35189\,
            I => \N__35186\
        );

    \I__7138\ : Odrv4
    port map (
            O => \N__35186\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\
        );

    \I__7137\ : InMux
    port map (
            O => \N__35183\,
            I => \N__35179\
        );

    \I__7136\ : InMux
    port map (
            O => \N__35182\,
            I => \N__35176\
        );

    \I__7135\ : LocalMux
    port map (
            O => \N__35179\,
            I => \N__35173\
        );

    \I__7134\ : LocalMux
    port map (
            O => \N__35176\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__7133\ : Odrv4
    port map (
            O => \N__35173\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__7132\ : CascadeMux
    port map (
            O => \N__35168\,
            I => \N__35165\
        );

    \I__7131\ : InMux
    port map (
            O => \N__35165\,
            I => \N__35162\
        );

    \I__7130\ : LocalMux
    port map (
            O => \N__35162\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\
        );

    \I__7129\ : InMux
    port map (
            O => \N__35159\,
            I => \N__35156\
        );

    \I__7128\ : LocalMux
    port map (
            O => \N__35156\,
            I => \N__35153\
        );

    \I__7127\ : Span4Mux_h
    port map (
            O => \N__35153\,
            I => \N__35150\
        );

    \I__7126\ : Span4Mux_h
    port map (
            O => \N__35150\,
            I => \N__35147\
        );

    \I__7125\ : Odrv4
    port map (
            O => \N__35147\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\
        );

    \I__7124\ : InMux
    port map (
            O => \N__35144\,
            I => \N__35140\
        );

    \I__7123\ : InMux
    port map (
            O => \N__35143\,
            I => \N__35137\
        );

    \I__7122\ : LocalMux
    port map (
            O => \N__35140\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__7121\ : LocalMux
    port map (
            O => \N__35137\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__7120\ : CascadeMux
    port map (
            O => \N__35132\,
            I => \N__35129\
        );

    \I__7119\ : InMux
    port map (
            O => \N__35129\,
            I => \N__35126\
        );

    \I__7118\ : LocalMux
    port map (
            O => \N__35126\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\
        );

    \I__7117\ : InMux
    port map (
            O => \N__35123\,
            I => \N__35120\
        );

    \I__7116\ : LocalMux
    port map (
            O => \N__35120\,
            I => \N__35117\
        );

    \I__7115\ : Odrv4
    port map (
            O => \N__35117\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\
        );

    \I__7114\ : InMux
    port map (
            O => \N__35114\,
            I => \N__35110\
        );

    \I__7113\ : InMux
    port map (
            O => \N__35113\,
            I => \N__35107\
        );

    \I__7112\ : LocalMux
    port map (
            O => \N__35110\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__7111\ : LocalMux
    port map (
            O => \N__35107\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__7110\ : CascadeMux
    port map (
            O => \N__35102\,
            I => \N__35099\
        );

    \I__7109\ : InMux
    port map (
            O => \N__35099\,
            I => \N__35096\
        );

    \I__7108\ : LocalMux
    port map (
            O => \N__35096\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\
        );

    \I__7107\ : InMux
    port map (
            O => \N__35093\,
            I => \N__35090\
        );

    \I__7106\ : LocalMux
    port map (
            O => \N__35090\,
            I => \N__35087\
        );

    \I__7105\ : Odrv4
    port map (
            O => \N__35087\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\
        );

    \I__7104\ : CascadeMux
    port map (
            O => \N__35084\,
            I => \N__35081\
        );

    \I__7103\ : InMux
    port map (
            O => \N__35081\,
            I => \N__35078\
        );

    \I__7102\ : LocalMux
    port map (
            O => \N__35078\,
            I => \N__35075\
        );

    \I__7101\ : Odrv12
    port map (
            O => \N__35075\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt16\
        );

    \I__7100\ : InMux
    port map (
            O => \N__35072\,
            I => \N__35068\
        );

    \I__7099\ : InMux
    port map (
            O => \N__35071\,
            I => \N__35065\
        );

    \I__7098\ : LocalMux
    port map (
            O => \N__35068\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__7097\ : LocalMux
    port map (
            O => \N__35065\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__7096\ : InMux
    port map (
            O => \N__35060\,
            I => \N__35057\
        );

    \I__7095\ : LocalMux
    port map (
            O => \N__35057\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\
        );

    \I__7094\ : CascadeMux
    port map (
            O => \N__35054\,
            I => \N__35051\
        );

    \I__7093\ : InMux
    port map (
            O => \N__35051\,
            I => \N__35048\
        );

    \I__7092\ : LocalMux
    port map (
            O => \N__35048\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\
        );

    \I__7091\ : InMux
    port map (
            O => \N__35045\,
            I => \N__35041\
        );

    \I__7090\ : InMux
    port map (
            O => \N__35044\,
            I => \N__35038\
        );

    \I__7089\ : LocalMux
    port map (
            O => \N__35041\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__7088\ : LocalMux
    port map (
            O => \N__35038\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__7087\ : CascadeMux
    port map (
            O => \N__35033\,
            I => \N__35030\
        );

    \I__7086\ : InMux
    port map (
            O => \N__35030\,
            I => \N__35027\
        );

    \I__7085\ : LocalMux
    port map (
            O => \N__35027\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\
        );

    \I__7084\ : InMux
    port map (
            O => \N__35024\,
            I => \N__35021\
        );

    \I__7083\ : LocalMux
    port map (
            O => \N__35021\,
            I => \N__35018\
        );

    \I__7082\ : Odrv4
    port map (
            O => \N__35018\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\
        );

    \I__7081\ : InMux
    port map (
            O => \N__35015\,
            I => \N__35011\
        );

    \I__7080\ : InMux
    port map (
            O => \N__35014\,
            I => \N__35008\
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__35011\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__7078\ : LocalMux
    port map (
            O => \N__35008\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__7077\ : CascadeMux
    port map (
            O => \N__35003\,
            I => \N__35000\
        );

    \I__7076\ : InMux
    port map (
            O => \N__35000\,
            I => \N__34997\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__34997\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\
        );

    \I__7074\ : InMux
    port map (
            O => \N__34994\,
            I => \N__34991\
        );

    \I__7073\ : LocalMux
    port map (
            O => \N__34991\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\
        );

    \I__7072\ : InMux
    port map (
            O => \N__34988\,
            I => \N__34984\
        );

    \I__7071\ : InMux
    port map (
            O => \N__34987\,
            I => \N__34981\
        );

    \I__7070\ : LocalMux
    port map (
            O => \N__34984\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__7069\ : LocalMux
    port map (
            O => \N__34981\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__7068\ : CascadeMux
    port map (
            O => \N__34976\,
            I => \N__34973\
        );

    \I__7067\ : InMux
    port map (
            O => \N__34973\,
            I => \N__34970\
        );

    \I__7066\ : LocalMux
    port map (
            O => \N__34970\,
            I => \N__34967\
        );

    \I__7065\ : Odrv4
    port map (
            O => \N__34967\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\
        );

    \I__7064\ : InMux
    port map (
            O => \N__34964\,
            I => \N__34960\
        );

    \I__7063\ : InMux
    port map (
            O => \N__34963\,
            I => \N__34957\
        );

    \I__7062\ : LocalMux
    port map (
            O => \N__34960\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__7061\ : LocalMux
    port map (
            O => \N__34957\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__7060\ : CascadeMux
    port map (
            O => \N__34952\,
            I => \N__34949\
        );

    \I__7059\ : InMux
    port map (
            O => \N__34949\,
            I => \N__34946\
        );

    \I__7058\ : LocalMux
    port map (
            O => \N__34946\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\
        );

    \I__7057\ : InMux
    port map (
            O => \N__34943\,
            I => \N__34940\
        );

    \I__7056\ : LocalMux
    port map (
            O => \N__34940\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\
        );

    \I__7055\ : InMux
    port map (
            O => \N__34937\,
            I => \N__34933\
        );

    \I__7054\ : InMux
    port map (
            O => \N__34936\,
            I => \N__34930\
        );

    \I__7053\ : LocalMux
    port map (
            O => \N__34933\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__7052\ : LocalMux
    port map (
            O => \N__34930\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__7051\ : CascadeMux
    port map (
            O => \N__34925\,
            I => \N__34922\
        );

    \I__7050\ : InMux
    port map (
            O => \N__34922\,
            I => \N__34919\
        );

    \I__7049\ : LocalMux
    port map (
            O => \N__34919\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\
        );

    \I__7048\ : InMux
    port map (
            O => \N__34916\,
            I => \N__34912\
        );

    \I__7047\ : InMux
    port map (
            O => \N__34915\,
            I => \N__34909\
        );

    \I__7046\ : LocalMux
    port map (
            O => \N__34912\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__7045\ : LocalMux
    port map (
            O => \N__34909\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__7044\ : CascadeMux
    port map (
            O => \N__34904\,
            I => \N__34901\
        );

    \I__7043\ : InMux
    port map (
            O => \N__34901\,
            I => \N__34898\
        );

    \I__7042\ : LocalMux
    port map (
            O => \N__34898\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\
        );

    \I__7041\ : InMux
    port map (
            O => \N__34895\,
            I => \N__34889\
        );

    \I__7040\ : InMux
    port map (
            O => \N__34894\,
            I => \N__34886\
        );

    \I__7039\ : InMux
    port map (
            O => \N__34893\,
            I => \N__34883\
        );

    \I__7038\ : InMux
    port map (
            O => \N__34892\,
            I => \N__34880\
        );

    \I__7037\ : LocalMux
    port map (
            O => \N__34889\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__7036\ : LocalMux
    port map (
            O => \N__34886\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__7035\ : LocalMux
    port map (
            O => \N__34883\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__7034\ : LocalMux
    port map (
            O => \N__34880\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__7033\ : IoInMux
    port map (
            O => \N__34871\,
            I => \N__34868\
        );

    \I__7032\ : LocalMux
    port map (
            O => \N__34868\,
            I => \N__34865\
        );

    \I__7031\ : Span4Mux_s1_v
    port map (
            O => \N__34865\,
            I => \N__34862\
        );

    \I__7030\ : Span4Mux_v
    port map (
            O => \N__34862\,
            I => \N__34857\
        );

    \I__7029\ : InMux
    port map (
            O => \N__34861\,
            I => \N__34854\
        );

    \I__7028\ : InMux
    port map (
            O => \N__34860\,
            I => \N__34851\
        );

    \I__7027\ : Odrv4
    port map (
            O => \N__34857\,
            I => s1_phy_c
        );

    \I__7026\ : LocalMux
    port map (
            O => \N__34854\,
            I => s1_phy_c
        );

    \I__7025\ : LocalMux
    port map (
            O => \N__34851\,
            I => s1_phy_c
        );

    \I__7024\ : CascadeMux
    port map (
            O => \N__34844\,
            I => \N__34839\
        );

    \I__7023\ : InMux
    port map (
            O => \N__34843\,
            I => \N__34835\
        );

    \I__7022\ : InMux
    port map (
            O => \N__34842\,
            I => \N__34832\
        );

    \I__7021\ : InMux
    port map (
            O => \N__34839\,
            I => \N__34829\
        );

    \I__7020\ : InMux
    port map (
            O => \N__34838\,
            I => \N__34826\
        );

    \I__7019\ : LocalMux
    port map (
            O => \N__34835\,
            I => \N__34823\
        );

    \I__7018\ : LocalMux
    port map (
            O => \N__34832\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__7017\ : LocalMux
    port map (
            O => \N__34829\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__7016\ : LocalMux
    port map (
            O => \N__34826\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__7015\ : Odrv4
    port map (
            O => \N__34823\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__7014\ : IoInMux
    port map (
            O => \N__34814\,
            I => \N__34811\
        );

    \I__7013\ : LocalMux
    port map (
            O => \N__34811\,
            I => \N__34808\
        );

    \I__7012\ : Span12Mux_s3_v
    port map (
            O => \N__34808\,
            I => \N__34805\
        );

    \I__7011\ : Odrv12
    port map (
            O => \N__34805\,
            I => s2_phy_c
        );

    \I__7010\ : InMux
    port map (
            O => \N__34802\,
            I => \N__34796\
        );

    \I__7009\ : InMux
    port map (
            O => \N__34801\,
            I => \N__34796\
        );

    \I__7008\ : LocalMux
    port map (
            O => \N__34796\,
            I => \N__34792\
        );

    \I__7007\ : InMux
    port map (
            O => \N__34795\,
            I => \N__34789\
        );

    \I__7006\ : Span4Mux_h
    port map (
            O => \N__34792\,
            I => \N__34786\
        );

    \I__7005\ : LocalMux
    port map (
            O => \N__34789\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__7004\ : Odrv4
    port map (
            O => \N__34786\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__7003\ : CascadeMux
    port map (
            O => \N__34781\,
            I => \N__34777\
        );

    \I__7002\ : CascadeMux
    port map (
            O => \N__34780\,
            I => \N__34774\
        );

    \I__7001\ : InMux
    port map (
            O => \N__34777\,
            I => \N__34771\
        );

    \I__7000\ : InMux
    port map (
            O => \N__34774\,
            I => \N__34768\
        );

    \I__6999\ : LocalMux
    port map (
            O => \N__34771\,
            I => \N__34762\
        );

    \I__6998\ : LocalMux
    port map (
            O => \N__34768\,
            I => \N__34762\
        );

    \I__6997\ : InMux
    port map (
            O => \N__34767\,
            I => \N__34759\
        );

    \I__6996\ : Span4Mux_h
    port map (
            O => \N__34762\,
            I => \N__34756\
        );

    \I__6995\ : LocalMux
    port map (
            O => \N__34759\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__6994\ : Odrv4
    port map (
            O => \N__34756\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__6993\ : InMux
    port map (
            O => \N__34751\,
            I => \N__34745\
        );

    \I__6992\ : InMux
    port map (
            O => \N__34750\,
            I => \N__34745\
        );

    \I__6991\ : LocalMux
    port map (
            O => \N__34745\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\
        );

    \I__6990\ : InMux
    port map (
            O => \N__34742\,
            I => \N__34739\
        );

    \I__6989\ : LocalMux
    port map (
            O => \N__34739\,
            I => \N__34736\
        );

    \I__6988\ : Odrv4
    port map (
            O => \N__34736\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\
        );

    \I__6987\ : CascadeMux
    port map (
            O => \N__34733\,
            I => \N__34730\
        );

    \I__6986\ : InMux
    port map (
            O => \N__34730\,
            I => \N__34725\
        );

    \I__6985\ : InMux
    port map (
            O => \N__34729\,
            I => \N__34722\
        );

    \I__6984\ : CascadeMux
    port map (
            O => \N__34728\,
            I => \N__34719\
        );

    \I__6983\ : LocalMux
    port map (
            O => \N__34725\,
            I => \N__34714\
        );

    \I__6982\ : LocalMux
    port map (
            O => \N__34722\,
            I => \N__34714\
        );

    \I__6981\ : InMux
    port map (
            O => \N__34719\,
            I => \N__34711\
        );

    \I__6980\ : Span4Mux_v
    port map (
            O => \N__34714\,
            I => \N__34708\
        );

    \I__6979\ : LocalMux
    port map (
            O => \N__34711\,
            I => \N__34703\
        );

    \I__6978\ : Span4Mux_h
    port map (
            O => \N__34708\,
            I => \N__34703\
        );

    \I__6977\ : Odrv4
    port map (
            O => \N__34703\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__6976\ : CascadeMux
    port map (
            O => \N__34700\,
            I => \N__34697\
        );

    \I__6975\ : InMux
    port map (
            O => \N__34697\,
            I => \N__34694\
        );

    \I__6974\ : LocalMux
    port map (
            O => \N__34694\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\
        );

    \I__6973\ : CascadeMux
    port map (
            O => \N__34691\,
            I => \N__34685\
        );

    \I__6972\ : InMux
    port map (
            O => \N__34690\,
            I => \N__34682\
        );

    \I__6971\ : InMux
    port map (
            O => \N__34689\,
            I => \N__34677\
        );

    \I__6970\ : InMux
    port map (
            O => \N__34688\,
            I => \N__34677\
        );

    \I__6969\ : InMux
    port map (
            O => \N__34685\,
            I => \N__34674\
        );

    \I__6968\ : LocalMux
    port map (
            O => \N__34682\,
            I => \N__34671\
        );

    \I__6967\ : LocalMux
    port map (
            O => \N__34677\,
            I => \N__34668\
        );

    \I__6966\ : LocalMux
    port map (
            O => \N__34674\,
            I => \N__34663\
        );

    \I__6965\ : Span4Mux_v
    port map (
            O => \N__34671\,
            I => \N__34663\
        );

    \I__6964\ : Sp12to4
    port map (
            O => \N__34668\,
            I => \N__34658\
        );

    \I__6963\ : Span4Mux_v
    port map (
            O => \N__34663\,
            I => \N__34655\
        );

    \I__6962\ : InMux
    port map (
            O => \N__34662\,
            I => \N__34652\
        );

    \I__6961\ : InMux
    port map (
            O => \N__34661\,
            I => \N__34649\
        );

    \I__6960\ : Span12Mux_v
    port map (
            O => \N__34658\,
            I => \N__34642\
        );

    \I__6959\ : Sp12to4
    port map (
            O => \N__34655\,
            I => \N__34642\
        );

    \I__6958\ : LocalMux
    port map (
            O => \N__34652\,
            I => \N__34642\
        );

    \I__6957\ : LocalMux
    port map (
            O => \N__34649\,
            I => phase_controller_inst1_state_4
        );

    \I__6956\ : Odrv12
    port map (
            O => \N__34642\,
            I => phase_controller_inst1_state_4
        );

    \I__6955\ : InMux
    port map (
            O => \N__34637\,
            I => \N__34634\
        );

    \I__6954\ : LocalMux
    port map (
            O => \N__34634\,
            I => \N__34630\
        );

    \I__6953\ : InMux
    port map (
            O => \N__34633\,
            I => \N__34627\
        );

    \I__6952\ : Span4Mux_h
    port map (
            O => \N__34630\,
            I => \N__34622\
        );

    \I__6951\ : LocalMux
    port map (
            O => \N__34627\,
            I => \N__34622\
        );

    \I__6950\ : Odrv4
    port map (
            O => \N__34622\,
            I => \phase_controller_inst1.time_passed_RNIE87F\
        );

    \I__6949\ : CascadeMux
    port map (
            O => \N__34619\,
            I => \N__34616\
        );

    \I__6948\ : InMux
    port map (
            O => \N__34616\,
            I => \N__34611\
        );

    \I__6947\ : InMux
    port map (
            O => \N__34615\,
            I => \N__34608\
        );

    \I__6946\ : InMux
    port map (
            O => \N__34614\,
            I => \N__34605\
        );

    \I__6945\ : LocalMux
    port map (
            O => \N__34611\,
            I => \N__34602\
        );

    \I__6944\ : LocalMux
    port map (
            O => \N__34608\,
            I => \N__34597\
        );

    \I__6943\ : LocalMux
    port map (
            O => \N__34605\,
            I => \N__34597\
        );

    \I__6942\ : Span4Mux_v
    port map (
            O => \N__34602\,
            I => \N__34592\
        );

    \I__6941\ : Span4Mux_v
    port map (
            O => \N__34597\,
            I => \N__34592\
        );

    \I__6940\ : Span4Mux_h
    port map (
            O => \N__34592\,
            I => \N__34589\
        );

    \I__6939\ : Span4Mux_h
    port map (
            O => \N__34589\,
            I => \N__34585\
        );

    \I__6938\ : InMux
    port map (
            O => \N__34588\,
            I => \N__34582\
        );

    \I__6937\ : Span4Mux_v
    port map (
            O => \N__34585\,
            I => \N__34579\
        );

    \I__6936\ : LocalMux
    port map (
            O => \N__34582\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__6935\ : Odrv4
    port map (
            O => \N__34579\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__6934\ : CascadeMux
    port map (
            O => \N__34574\,
            I => \N__34569\
        );

    \I__6933\ : CascadeMux
    port map (
            O => \N__34573\,
            I => \N__34566\
        );

    \I__6932\ : InMux
    port map (
            O => \N__34572\,
            I => \N__34561\
        );

    \I__6931\ : InMux
    port map (
            O => \N__34569\,
            I => \N__34561\
        );

    \I__6930\ : InMux
    port map (
            O => \N__34566\,
            I => \N__34558\
        );

    \I__6929\ : LocalMux
    port map (
            O => \N__34561\,
            I => \N__34555\
        );

    \I__6928\ : LocalMux
    port map (
            O => \N__34558\,
            I => \N__34552\
        );

    \I__6927\ : Span4Mux_v
    port map (
            O => \N__34555\,
            I => \N__34547\
        );

    \I__6926\ : Span4Mux_v
    port map (
            O => \N__34552\,
            I => \N__34547\
        );

    \I__6925\ : Odrv4
    port map (
            O => \N__34547\,
            I => \il_min_comp1_D2\
        );

    \I__6924\ : InMux
    port map (
            O => \N__34544\,
            I => \N__34541\
        );

    \I__6923\ : LocalMux
    port map (
            O => \N__34541\,
            I => \N__34538\
        );

    \I__6922\ : Odrv4
    port map (
            O => \N__34538\,
            I => \phase_controller_inst1.start_timer_tr_RNOZ0Z_0\
        );

    \I__6921\ : InMux
    port map (
            O => \N__34535\,
            I => \N__34530\
        );

    \I__6920\ : InMux
    port map (
            O => \N__34534\,
            I => \N__34526\
        );

    \I__6919\ : InMux
    port map (
            O => \N__34533\,
            I => \N__34523\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__34530\,
            I => \N__34520\
        );

    \I__6917\ : InMux
    port map (
            O => \N__34529\,
            I => \N__34517\
        );

    \I__6916\ : LocalMux
    port map (
            O => \N__34526\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__6915\ : LocalMux
    port map (
            O => \N__34523\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__6914\ : Odrv4
    port map (
            O => \N__34520\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__6913\ : LocalMux
    port map (
            O => \N__34517\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__6912\ : InMux
    port map (
            O => \N__34508\,
            I => \N__34505\
        );

    \I__6911\ : LocalMux
    port map (
            O => \N__34505\,
            I => \N__34502\
        );

    \I__6910\ : Odrv4
    port map (
            O => \N__34502\,
            I => \current_shift_inst.un38_control_input_0_s0_30\
        );

    \I__6909\ : InMux
    port map (
            O => \N__34499\,
            I => \current_shift_inst.un38_control_input_cry_29_s0\
        );

    \I__6908\ : InMux
    port map (
            O => \N__34496\,
            I => \N__34493\
        );

    \I__6907\ : LocalMux
    port map (
            O => \N__34493\,
            I => \N__34490\
        );

    \I__6906\ : Span4Mux_h
    port map (
            O => \N__34490\,
            I => \N__34487\
        );

    \I__6905\ : Odrv4
    port map (
            O => \N__34487\,
            I => \current_shift_inst.un38_control_input_0_s1_31\
        );

    \I__6904\ : InMux
    port map (
            O => \N__34484\,
            I => \current_shift_inst.un38_control_input_cry_30_s0\
        );

    \I__6903\ : InMux
    port map (
            O => \N__34481\,
            I => \N__34478\
        );

    \I__6902\ : LocalMux
    port map (
            O => \N__34478\,
            I => \N__34475\
        );

    \I__6901\ : Span4Mux_h
    port map (
            O => \N__34475\,
            I => \N__34472\
        );

    \I__6900\ : Span4Mux_v
    port map (
            O => \N__34472\,
            I => \N__34469\
        );

    \I__6899\ : Odrv4
    port map (
            O => \N__34469\,
            I => \current_shift_inst.control_input_axb_11\
        );

    \I__6898\ : InMux
    port map (
            O => \N__34466\,
            I => \N__34463\
        );

    \I__6897\ : LocalMux
    port map (
            O => \N__34463\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\
        );

    \I__6896\ : InMux
    port map (
            O => \N__34460\,
            I => \N__34457\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__34457\,
            I => \N__34454\
        );

    \I__6894\ : Odrv12
    port map (
            O => \N__34454\,
            I => \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\
        );

    \I__6893\ : InMux
    port map (
            O => \N__34451\,
            I => \N__34448\
        );

    \I__6892\ : LocalMux
    port map (
            O => \N__34448\,
            I => \N__34445\
        );

    \I__6891\ : Span4Mux_h
    port map (
            O => \N__34445\,
            I => \N__34442\
        );

    \I__6890\ : Odrv4
    port map (
            O => \N__34442\,
            I => \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0\
        );

    \I__6889\ : CascadeMux
    port map (
            O => \N__34439\,
            I => \N__34436\
        );

    \I__6888\ : InMux
    port map (
            O => \N__34436\,
            I => \N__34433\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__34433\,
            I => \N__34430\
        );

    \I__6886\ : Odrv4
    port map (
            O => \N__34430\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\
        );

    \I__6885\ : InMux
    port map (
            O => \N__34427\,
            I => \current_shift_inst.un38_control_input_cry_20_s0\
        );

    \I__6884\ : CascadeMux
    port map (
            O => \N__34424\,
            I => \N__34421\
        );

    \I__6883\ : InMux
    port map (
            O => \N__34421\,
            I => \N__34418\
        );

    \I__6882\ : LocalMux
    port map (
            O => \N__34418\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\
        );

    \I__6881\ : InMux
    port map (
            O => \N__34415\,
            I => \N__34412\
        );

    \I__6880\ : LocalMux
    port map (
            O => \N__34412\,
            I => \N__34409\
        );

    \I__6879\ : Odrv4
    port map (
            O => \N__34409\,
            I => \current_shift_inst.un38_control_input_0_s0_22\
        );

    \I__6878\ : InMux
    port map (
            O => \N__34406\,
            I => \current_shift_inst.un38_control_input_cry_21_s0\
        );

    \I__6877\ : InMux
    port map (
            O => \N__34403\,
            I => \N__34400\
        );

    \I__6876\ : LocalMux
    port map (
            O => \N__34400\,
            I => \N__34397\
        );

    \I__6875\ : Odrv4
    port map (
            O => \N__34397\,
            I => \current_shift_inst.un38_control_input_0_s0_23\
        );

    \I__6874\ : InMux
    port map (
            O => \N__34394\,
            I => \current_shift_inst.un38_control_input_cry_22_s0\
        );

    \I__6873\ : InMux
    port map (
            O => \N__34391\,
            I => \N__34388\
        );

    \I__6872\ : LocalMux
    port map (
            O => \N__34388\,
            I => \current_shift_inst.un38_control_input_0_s0_24\
        );

    \I__6871\ : InMux
    port map (
            O => \N__34385\,
            I => \bfn_14_16_0_\
        );

    \I__6870\ : InMux
    port map (
            O => \N__34382\,
            I => \N__34379\
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__34379\,
            I => \current_shift_inst.un38_control_input_0_s0_25\
        );

    \I__6868\ : InMux
    port map (
            O => \N__34376\,
            I => \current_shift_inst.un38_control_input_cry_24_s0\
        );

    \I__6867\ : InMux
    port map (
            O => \N__34373\,
            I => \N__34370\
        );

    \I__6866\ : LocalMux
    port map (
            O => \N__34370\,
            I => \current_shift_inst.un38_control_input_0_s0_26\
        );

    \I__6865\ : InMux
    port map (
            O => \N__34367\,
            I => \current_shift_inst.un38_control_input_cry_25_s0\
        );

    \I__6864\ : InMux
    port map (
            O => \N__34364\,
            I => \N__34361\
        );

    \I__6863\ : LocalMux
    port map (
            O => \N__34361\,
            I => \current_shift_inst.un38_control_input_0_s0_27\
        );

    \I__6862\ : InMux
    port map (
            O => \N__34358\,
            I => \current_shift_inst.un38_control_input_cry_26_s0\
        );

    \I__6861\ : InMux
    port map (
            O => \N__34355\,
            I => \N__34352\
        );

    \I__6860\ : LocalMux
    port map (
            O => \N__34352\,
            I => \N__34349\
        );

    \I__6859\ : Odrv4
    port map (
            O => \N__34349\,
            I => \current_shift_inst.un38_control_input_0_s0_28\
        );

    \I__6858\ : InMux
    port map (
            O => \N__34346\,
            I => \current_shift_inst.un38_control_input_cry_27_s0\
        );

    \I__6857\ : InMux
    port map (
            O => \N__34343\,
            I => \N__34340\
        );

    \I__6856\ : LocalMux
    port map (
            O => \N__34340\,
            I => \N__34337\
        );

    \I__6855\ : Odrv4
    port map (
            O => \N__34337\,
            I => \current_shift_inst.un38_control_input_0_s0_29\
        );

    \I__6854\ : InMux
    port map (
            O => \N__34334\,
            I => \current_shift_inst.un38_control_input_cry_28_s0\
        );

    \I__6853\ : InMux
    port map (
            O => \N__34331\,
            I => \N__34328\
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__34328\,
            I => \N__34325\
        );

    \I__6851\ : Span4Mux_h
    port map (
            O => \N__34325\,
            I => \N__34322\
        );

    \I__6850\ : Odrv4
    port map (
            O => \N__34322\,
            I => \current_shift_inst.un38_control_input_0_s0_20\
        );

    \I__6849\ : InMux
    port map (
            O => \N__34319\,
            I => \current_shift_inst.un38_control_input_cry_19_s0\
        );

    \I__6848\ : InMux
    port map (
            O => \N__34316\,
            I => \N__34313\
        );

    \I__6847\ : LocalMux
    port map (
            O => \N__34313\,
            I => \N__34310\
        );

    \I__6846\ : Odrv4
    port map (
            O => \N__34310\,
            I => \current_shift_inst.un38_control_input_0_s0_21\
        );

    \I__6845\ : CascadeMux
    port map (
            O => \N__34307\,
            I => \N__34304\
        );

    \I__6844\ : InMux
    port map (
            O => \N__34304\,
            I => \N__34301\
        );

    \I__6843\ : LocalMux
    port map (
            O => \N__34301\,
            I => \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0\
        );

    \I__6842\ : CascadeMux
    port map (
            O => \N__34298\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30_cascade_\
        );

    \I__6841\ : InMux
    port map (
            O => \N__34295\,
            I => \N__34292\
        );

    \I__6840\ : LocalMux
    port map (
            O => \N__34292\,
            I => \N__34288\
        );

    \I__6839\ : InMux
    port map (
            O => \N__34291\,
            I => \N__34285\
        );

    \I__6838\ : Odrv4
    port map (
            O => \N__34288\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__6837\ : LocalMux
    port map (
            O => \N__34285\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__6836\ : CascadeMux
    port map (
            O => \N__34280\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31_cascade_\
        );

    \I__6835\ : InMux
    port map (
            O => \N__34277\,
            I => \N__34274\
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__34274\,
            I => \N__34270\
        );

    \I__6833\ : InMux
    port map (
            O => \N__34273\,
            I => \N__34267\
        );

    \I__6832\ : Odrv4
    port map (
            O => \N__34270\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13\
        );

    \I__6831\ : LocalMux
    port map (
            O => \N__34267\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13\
        );

    \I__6830\ : InMux
    port map (
            O => \N__34262\,
            I => \N__34258\
        );

    \I__6829\ : InMux
    port map (
            O => \N__34261\,
            I => \N__34255\
        );

    \I__6828\ : LocalMux
    port map (
            O => \N__34258\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__6827\ : LocalMux
    port map (
            O => \N__34255\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__6826\ : CascadeMux
    port map (
            O => \N__34250\,
            I => \N__34247\
        );

    \I__6825\ : InMux
    port map (
            O => \N__34247\,
            I => \N__34244\
        );

    \I__6824\ : LocalMux
    port map (
            O => \N__34244\,
            I => \N__34241\
        );

    \I__6823\ : Odrv12
    port map (
            O => \N__34241\,
            I => \current_shift_inst.un38_control_input_cry_0_s0_sf\
        );

    \I__6822\ : CascadeMux
    port map (
            O => \N__34238\,
            I => \N__34235\
        );

    \I__6821\ : InMux
    port map (
            O => \N__34235\,
            I => \N__34232\
        );

    \I__6820\ : LocalMux
    port map (
            O => \N__34232\,
            I => \N__34229\
        );

    \I__6819\ : Span4Mux_h
    port map (
            O => \N__34229\,
            I => \N__34226\
        );

    \I__6818\ : Odrv4
    port map (
            O => \N__34226\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\
        );

    \I__6817\ : InMux
    port map (
            O => \N__34223\,
            I => \bfn_14_11_0_\
        );

    \I__6816\ : InMux
    port map (
            O => \N__34220\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\
        );

    \I__6815\ : InMux
    port map (
            O => \N__34217\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\
        );

    \I__6814\ : InMux
    port map (
            O => \N__34214\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\
        );

    \I__6813\ : InMux
    port map (
            O => \N__34211\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\
        );

    \I__6812\ : InMux
    port map (
            O => \N__34208\,
            I => \N__34198\
        );

    \I__6811\ : InMux
    port map (
            O => \N__34207\,
            I => \N__34198\
        );

    \I__6810\ : InMux
    port map (
            O => \N__34206\,
            I => \N__34198\
        );

    \I__6809\ : InMux
    port map (
            O => \N__34205\,
            I => \N__34195\
        );

    \I__6808\ : LocalMux
    port map (
            O => \N__34198\,
            I => \N__34192\
        );

    \I__6807\ : LocalMux
    port map (
            O => \N__34195\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__6806\ : Odrv4
    port map (
            O => \N__34192\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__6805\ : InMux
    port map (
            O => \N__34187\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\
        );

    \I__6804\ : InMux
    port map (
            O => \N__34184\,
            I => \N__34152\
        );

    \I__6803\ : InMux
    port map (
            O => \N__34183\,
            I => \N__34152\
        );

    \I__6802\ : InMux
    port map (
            O => \N__34182\,
            I => \N__34152\
        );

    \I__6801\ : InMux
    port map (
            O => \N__34181\,
            I => \N__34152\
        );

    \I__6800\ : IoInMux
    port map (
            O => \N__34180\,
            I => \N__34149\
        );

    \I__6799\ : InMux
    port map (
            O => \N__34179\,
            I => \N__34133\
        );

    \I__6798\ : InMux
    port map (
            O => \N__34178\,
            I => \N__34133\
        );

    \I__6797\ : InMux
    port map (
            O => \N__34177\,
            I => \N__34133\
        );

    \I__6796\ : InMux
    port map (
            O => \N__34176\,
            I => \N__34133\
        );

    \I__6795\ : InMux
    port map (
            O => \N__34175\,
            I => \N__34126\
        );

    \I__6794\ : InMux
    port map (
            O => \N__34174\,
            I => \N__34126\
        );

    \I__6793\ : InMux
    port map (
            O => \N__34173\,
            I => \N__34126\
        );

    \I__6792\ : InMux
    port map (
            O => \N__34172\,
            I => \N__34117\
        );

    \I__6791\ : InMux
    port map (
            O => \N__34171\,
            I => \N__34117\
        );

    \I__6790\ : InMux
    port map (
            O => \N__34170\,
            I => \N__34117\
        );

    \I__6789\ : InMux
    port map (
            O => \N__34169\,
            I => \N__34117\
        );

    \I__6788\ : InMux
    port map (
            O => \N__34168\,
            I => \N__34108\
        );

    \I__6787\ : InMux
    port map (
            O => \N__34167\,
            I => \N__34108\
        );

    \I__6786\ : InMux
    port map (
            O => \N__34166\,
            I => \N__34108\
        );

    \I__6785\ : InMux
    port map (
            O => \N__34165\,
            I => \N__34108\
        );

    \I__6784\ : InMux
    port map (
            O => \N__34164\,
            I => \N__34099\
        );

    \I__6783\ : InMux
    port map (
            O => \N__34163\,
            I => \N__34099\
        );

    \I__6782\ : InMux
    port map (
            O => \N__34162\,
            I => \N__34099\
        );

    \I__6781\ : InMux
    port map (
            O => \N__34161\,
            I => \N__34099\
        );

    \I__6780\ : LocalMux
    port map (
            O => \N__34152\,
            I => \N__34096\
        );

    \I__6779\ : LocalMux
    port map (
            O => \N__34149\,
            I => \N__34093\
        );

    \I__6778\ : InMux
    port map (
            O => \N__34148\,
            I => \N__34083\
        );

    \I__6777\ : InMux
    port map (
            O => \N__34147\,
            I => \N__34083\
        );

    \I__6776\ : InMux
    port map (
            O => \N__34146\,
            I => \N__34083\
        );

    \I__6775\ : InMux
    port map (
            O => \N__34145\,
            I => \N__34083\
        );

    \I__6774\ : InMux
    port map (
            O => \N__34144\,
            I => \N__34076\
        );

    \I__6773\ : InMux
    port map (
            O => \N__34143\,
            I => \N__34076\
        );

    \I__6772\ : InMux
    port map (
            O => \N__34142\,
            I => \N__34076\
        );

    \I__6771\ : LocalMux
    port map (
            O => \N__34133\,
            I => \N__34073\
        );

    \I__6770\ : LocalMux
    port map (
            O => \N__34126\,
            I => \N__34064\
        );

    \I__6769\ : LocalMux
    port map (
            O => \N__34117\,
            I => \N__34064\
        );

    \I__6768\ : LocalMux
    port map (
            O => \N__34108\,
            I => \N__34064\
        );

    \I__6767\ : LocalMux
    port map (
            O => \N__34099\,
            I => \N__34064\
        );

    \I__6766\ : Span4Mux_h
    port map (
            O => \N__34096\,
            I => \N__34061\
        );

    \I__6765\ : Span4Mux_s0_v
    port map (
            O => \N__34093\,
            I => \N__34058\
        );

    \I__6764\ : InMux
    port map (
            O => \N__34092\,
            I => \N__34055\
        );

    \I__6763\ : LocalMux
    port map (
            O => \N__34083\,
            I => \N__34046\
        );

    \I__6762\ : LocalMux
    port map (
            O => \N__34076\,
            I => \N__34046\
        );

    \I__6761\ : Span4Mux_v
    port map (
            O => \N__34073\,
            I => \N__34046\
        );

    \I__6760\ : Span4Mux_v
    port map (
            O => \N__34064\,
            I => \N__34046\
        );

    \I__6759\ : Span4Mux_v
    port map (
            O => \N__34061\,
            I => \N__34041\
        );

    \I__6758\ : Span4Mux_v
    port map (
            O => \N__34058\,
            I => \N__34041\
        );

    \I__6757\ : LocalMux
    port map (
            O => \N__34055\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__6756\ : Odrv4
    port map (
            O => \N__34046\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__6755\ : Odrv4
    port map (
            O => \N__34041\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__6754\ : InMux
    port map (
            O => \N__34034\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\
        );

    \I__6753\ : CascadeMux
    port map (
            O => \N__34031\,
            I => \N__34027\
        );

    \I__6752\ : CascadeMux
    port map (
            O => \N__34030\,
            I => \N__34024\
        );

    \I__6751\ : InMux
    port map (
            O => \N__34027\,
            I => \N__34016\
        );

    \I__6750\ : InMux
    port map (
            O => \N__34024\,
            I => \N__34016\
        );

    \I__6749\ : InMux
    port map (
            O => \N__34023\,
            I => \N__34016\
        );

    \I__6748\ : LocalMux
    port map (
            O => \N__34016\,
            I => \N__34012\
        );

    \I__6747\ : InMux
    port map (
            O => \N__34015\,
            I => \N__34009\
        );

    \I__6746\ : Span4Mux_v
    port map (
            O => \N__34012\,
            I => \N__34006\
        );

    \I__6745\ : LocalMux
    port map (
            O => \N__34009\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__6744\ : Odrv4
    port map (
            O => \N__34006\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__6743\ : InMux
    port map (
            O => \N__34001\,
            I => \N__33998\
        );

    \I__6742\ : LocalMux
    port map (
            O => \N__33998\,
            I => \N__33994\
        );

    \I__6741\ : InMux
    port map (
            O => \N__33997\,
            I => \N__33991\
        );

    \I__6740\ : Odrv4
    port map (
            O => \N__33994\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30\
        );

    \I__6739\ : LocalMux
    port map (
            O => \N__33991\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30\
        );

    \I__6738\ : InMux
    port map (
            O => \N__33986\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\
        );

    \I__6737\ : InMux
    port map (
            O => \N__33983\,
            I => \bfn_14_10_0_\
        );

    \I__6736\ : InMux
    port map (
            O => \N__33980\,
            I => \N__33973\
        );

    \I__6735\ : InMux
    port map (
            O => \N__33979\,
            I => \N__33973\
        );

    \I__6734\ : InMux
    port map (
            O => \N__33978\,
            I => \N__33970\
        );

    \I__6733\ : LocalMux
    port map (
            O => \N__33973\,
            I => \N__33967\
        );

    \I__6732\ : LocalMux
    port map (
            O => \N__33970\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__6731\ : Odrv4
    port map (
            O => \N__33967\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__6730\ : InMux
    port map (
            O => \N__33962\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\
        );

    \I__6729\ : CascadeMux
    port map (
            O => \N__33959\,
            I => \N__33956\
        );

    \I__6728\ : InMux
    port map (
            O => \N__33956\,
            I => \N__33949\
        );

    \I__6727\ : InMux
    port map (
            O => \N__33955\,
            I => \N__33949\
        );

    \I__6726\ : InMux
    port map (
            O => \N__33954\,
            I => \N__33946\
        );

    \I__6725\ : LocalMux
    port map (
            O => \N__33949\,
            I => \N__33943\
        );

    \I__6724\ : LocalMux
    port map (
            O => \N__33946\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__6723\ : Odrv4
    port map (
            O => \N__33943\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__6722\ : InMux
    port map (
            O => \N__33938\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\
        );

    \I__6721\ : InMux
    port map (
            O => \N__33935\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\
        );

    \I__6720\ : InMux
    port map (
            O => \N__33932\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__6719\ : InMux
    port map (
            O => \N__33929\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\
        );

    \I__6718\ : InMux
    port map (
            O => \N__33926\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\
        );

    \I__6717\ : InMux
    port map (
            O => \N__33923\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\
        );

    \I__6716\ : InMux
    port map (
            O => \N__33920\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\
        );

    \I__6715\ : InMux
    port map (
            O => \N__33917\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\
        );

    \I__6714\ : InMux
    port map (
            O => \N__33914\,
            I => \bfn_14_9_0_\
        );

    \I__6713\ : InMux
    port map (
            O => \N__33911\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\
        );

    \I__6712\ : InMux
    port map (
            O => \N__33908\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\
        );

    \I__6711\ : InMux
    port map (
            O => \N__33905\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\
        );

    \I__6710\ : InMux
    port map (
            O => \N__33902\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\
        );

    \I__6709\ : InMux
    port map (
            O => \N__33899\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\
        );

    \I__6708\ : InMux
    port map (
            O => \N__33896\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\
        );

    \I__6707\ : CascadeMux
    port map (
            O => \N__33893\,
            I => \N__33890\
        );

    \I__6706\ : InMux
    port map (
            O => \N__33890\,
            I => \N__33884\
        );

    \I__6705\ : InMux
    port map (
            O => \N__33889\,
            I => \N__33884\
        );

    \I__6704\ : LocalMux
    port map (
            O => \N__33884\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\
        );

    \I__6703\ : InMux
    port map (
            O => \N__33881\,
            I => \N__33878\
        );

    \I__6702\ : LocalMux
    port map (
            O => \N__33878\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\
        );

    \I__6701\ : InMux
    port map (
            O => \N__33875\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\
        );

    \I__6700\ : CascadeMux
    port map (
            O => \N__33872\,
            I => \N__33869\
        );

    \I__6699\ : InMux
    port map (
            O => \N__33869\,
            I => \N__33866\
        );

    \I__6698\ : LocalMux
    port map (
            O => \N__33866\,
            I => \N__33863\
        );

    \I__6697\ : Odrv4
    port map (
            O => \N__33863\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34Z0Z_28\
        );

    \I__6696\ : InMux
    port map (
            O => \N__33860\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\
        );

    \I__6695\ : InMux
    port map (
            O => \N__33857\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\
        );

    \I__6694\ : InMux
    port map (
            O => \N__33854\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\
        );

    \I__6693\ : InMux
    port map (
            O => \N__33851\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\
        );

    \I__6692\ : InMux
    port map (
            O => \N__33848\,
            I => \N__33842\
        );

    \I__6691\ : InMux
    port map (
            O => \N__33847\,
            I => \N__33842\
        );

    \I__6690\ : LocalMux
    port map (
            O => \N__33842\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\
        );

    \I__6689\ : InMux
    port map (
            O => \N__33839\,
            I => \N__33836\
        );

    \I__6688\ : LocalMux
    port map (
            O => \N__33836\,
            I => \current_shift_inst.un38_control_input_0_s1_29\
        );

    \I__6687\ : InMux
    port map (
            O => \N__33833\,
            I => \N__33830\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__33830\,
            I => \N__33827\
        );

    \I__6685\ : Span4Mux_h
    port map (
            O => \N__33827\,
            I => \N__33824\
        );

    \I__6684\ : Odrv4
    port map (
            O => \N__33824\,
            I => \current_shift_inst.control_input_axb_9\
        );

    \I__6683\ : InMux
    port map (
            O => \N__33821\,
            I => \N__33818\
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__33818\,
            I => \current_shift_inst.un38_control_input_0_s1_30\
        );

    \I__6681\ : InMux
    port map (
            O => \N__33815\,
            I => \N__33812\
        );

    \I__6680\ : LocalMux
    port map (
            O => \N__33812\,
            I => \N__33809\
        );

    \I__6679\ : Span4Mux_v
    port map (
            O => \N__33809\,
            I => \N__33806\
        );

    \I__6678\ : Odrv4
    port map (
            O => \N__33806\,
            I => \current_shift_inst.control_input_axb_10\
        );

    \I__6677\ : CascadeMux
    port map (
            O => \N__33803\,
            I => \N__33800\
        );

    \I__6676\ : InMux
    port map (
            O => \N__33800\,
            I => \N__33797\
        );

    \I__6675\ : LocalMux
    port map (
            O => \N__33797\,
            I => \N__33794\
        );

    \I__6674\ : Odrv4
    port map (
            O => \N__33794\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\
        );

    \I__6673\ : InMux
    port map (
            O => \N__33791\,
            I => \N__33788\
        );

    \I__6672\ : LocalMux
    port map (
            O => \N__33788\,
            I => \N__33784\
        );

    \I__6671\ : InMux
    port map (
            O => \N__33787\,
            I => \N__33781\
        );

    \I__6670\ : Span4Mux_v
    port map (
            O => \N__33784\,
            I => \N__33778\
        );

    \I__6669\ : LocalMux
    port map (
            O => \N__33781\,
            I => \N__33775\
        );

    \I__6668\ : Span4Mux_v
    port map (
            O => \N__33778\,
            I => \N__33772\
        );

    \I__6667\ : Span4Mux_v
    port map (
            O => \N__33775\,
            I => \N__33769\
        );

    \I__6666\ : Odrv4
    port map (
            O => \N__33772\,
            I => state_ns_i_a2_1
        );

    \I__6665\ : Odrv4
    port map (
            O => \N__33769\,
            I => state_ns_i_a2_1
        );

    \I__6664\ : InMux
    port map (
            O => \N__33764\,
            I => \N__33757\
        );

    \I__6663\ : InMux
    port map (
            O => \N__33763\,
            I => \N__33757\
        );

    \I__6662\ : InMux
    port map (
            O => \N__33762\,
            I => \N__33754\
        );

    \I__6661\ : LocalMux
    port map (
            O => \N__33757\,
            I => \N__33751\
        );

    \I__6660\ : LocalMux
    port map (
            O => \N__33754\,
            I => \N__33748\
        );

    \I__6659\ : Span4Mux_v
    port map (
            O => \N__33751\,
            I => \N__33745\
        );

    \I__6658\ : Span4Mux_h
    port map (
            O => \N__33748\,
            I => \N__33742\
        );

    \I__6657\ : Sp12to4
    port map (
            O => \N__33745\,
            I => \N__33738\
        );

    \I__6656\ : Span4Mux_h
    port map (
            O => \N__33742\,
            I => \N__33735\
        );

    \I__6655\ : InMux
    port map (
            O => \N__33741\,
            I => \N__33732\
        );

    \I__6654\ : Span12Mux_h
    port map (
            O => \N__33738\,
            I => \N__33729\
        );

    \I__6653\ : Odrv4
    port map (
            O => \N__33735\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__6652\ : LocalMux
    port map (
            O => \N__33732\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__6651\ : Odrv12
    port map (
            O => \N__33729\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__6650\ : InMux
    port map (
            O => \N__33722\,
            I => \N__33719\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__33719\,
            I => \phase_controller_inst1.start_timer_hc_0_sqmuxa\
        );

    \I__6648\ : CascadeMux
    port map (
            O => \N__33716\,
            I => \N__33712\
        );

    \I__6647\ : InMux
    port map (
            O => \N__33715\,
            I => \N__33709\
        );

    \I__6646\ : InMux
    port map (
            O => \N__33712\,
            I => \N__33705\
        );

    \I__6645\ : LocalMux
    port map (
            O => \N__33709\,
            I => \N__33702\
        );

    \I__6644\ : InMux
    port map (
            O => \N__33708\,
            I => \N__33699\
        );

    \I__6643\ : LocalMux
    port map (
            O => \N__33705\,
            I => \N__33692\
        );

    \I__6642\ : Span4Mux_v
    port map (
            O => \N__33702\,
            I => \N__33692\
        );

    \I__6641\ : LocalMux
    port map (
            O => \N__33699\,
            I => \N__33692\
        );

    \I__6640\ : Span4Mux_v
    port map (
            O => \N__33692\,
            I => \N__33689\
        );

    \I__6639\ : Odrv4
    port map (
            O => \N__33689\,
            I => \il_max_comp1_D2\
        );

    \I__6638\ : IoInMux
    port map (
            O => \N__33686\,
            I => \N__33683\
        );

    \I__6637\ : LocalMux
    port map (
            O => \N__33683\,
            I => \N__33680\
        );

    \I__6636\ : Odrv12
    port map (
            O => \N__33680\,
            I => \current_shift_inst.timer_s1.N_162_i\
        );

    \I__6635\ : InMux
    port map (
            O => \N__33677\,
            I => \N__33674\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__33674\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\
        );

    \I__6633\ : InMux
    port map (
            O => \N__33671\,
            I => \N__33668\
        );

    \I__6632\ : LocalMux
    port map (
            O => \N__33668\,
            I => \current_shift_inst.un38_control_input_0_s1_22\
        );

    \I__6631\ : InMux
    port map (
            O => \N__33665\,
            I => \N__33662\
        );

    \I__6630\ : LocalMux
    port map (
            O => \N__33662\,
            I => \N__33659\
        );

    \I__6629\ : Span4Mux_v
    port map (
            O => \N__33659\,
            I => \N__33656\
        );

    \I__6628\ : Odrv4
    port map (
            O => \N__33656\,
            I => \current_shift_inst.control_input_axb_2\
        );

    \I__6627\ : InMux
    port map (
            O => \N__33653\,
            I => \N__33650\
        );

    \I__6626\ : LocalMux
    port map (
            O => \N__33650\,
            I => \current_shift_inst.un38_control_input_0_s1_23\
        );

    \I__6625\ : InMux
    port map (
            O => \N__33647\,
            I => \N__33644\
        );

    \I__6624\ : LocalMux
    port map (
            O => \N__33644\,
            I => \N__33641\
        );

    \I__6623\ : Span4Mux_v
    port map (
            O => \N__33641\,
            I => \N__33638\
        );

    \I__6622\ : Odrv4
    port map (
            O => \N__33638\,
            I => \current_shift_inst.control_input_axb_3\
        );

    \I__6621\ : InMux
    port map (
            O => \N__33635\,
            I => \N__33632\
        );

    \I__6620\ : LocalMux
    port map (
            O => \N__33632\,
            I => \current_shift_inst.un38_control_input_0_s1_24\
        );

    \I__6619\ : InMux
    port map (
            O => \N__33629\,
            I => \N__33626\
        );

    \I__6618\ : LocalMux
    port map (
            O => \N__33626\,
            I => \N__33623\
        );

    \I__6617\ : Span4Mux_h
    port map (
            O => \N__33623\,
            I => \N__33620\
        );

    \I__6616\ : Odrv4
    port map (
            O => \N__33620\,
            I => \current_shift_inst.control_input_axb_4\
        );

    \I__6615\ : InMux
    port map (
            O => \N__33617\,
            I => \N__33614\
        );

    \I__6614\ : LocalMux
    port map (
            O => \N__33614\,
            I => \current_shift_inst.un38_control_input_0_s1_25\
        );

    \I__6613\ : InMux
    port map (
            O => \N__33611\,
            I => \N__33608\
        );

    \I__6612\ : LocalMux
    port map (
            O => \N__33608\,
            I => \N__33605\
        );

    \I__6611\ : Span4Mux_h
    port map (
            O => \N__33605\,
            I => \N__33602\
        );

    \I__6610\ : Odrv4
    port map (
            O => \N__33602\,
            I => \current_shift_inst.control_input_axb_5\
        );

    \I__6609\ : InMux
    port map (
            O => \N__33599\,
            I => \N__33596\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__33596\,
            I => \current_shift_inst.un38_control_input_0_s1_26\
        );

    \I__6607\ : InMux
    port map (
            O => \N__33593\,
            I => \N__33590\
        );

    \I__6606\ : LocalMux
    port map (
            O => \N__33590\,
            I => \N__33587\
        );

    \I__6605\ : Span4Mux_h
    port map (
            O => \N__33587\,
            I => \N__33584\
        );

    \I__6604\ : Odrv4
    port map (
            O => \N__33584\,
            I => \current_shift_inst.control_input_axb_6\
        );

    \I__6603\ : InMux
    port map (
            O => \N__33581\,
            I => \N__33578\
        );

    \I__6602\ : LocalMux
    port map (
            O => \N__33578\,
            I => \current_shift_inst.un38_control_input_0_s1_27\
        );

    \I__6601\ : InMux
    port map (
            O => \N__33575\,
            I => \N__33572\
        );

    \I__6600\ : LocalMux
    port map (
            O => \N__33572\,
            I => \N__33569\
        );

    \I__6599\ : Span4Mux_h
    port map (
            O => \N__33569\,
            I => \N__33566\
        );

    \I__6598\ : Odrv4
    port map (
            O => \N__33566\,
            I => \current_shift_inst.control_input_axb_7\
        );

    \I__6597\ : InMux
    port map (
            O => \N__33563\,
            I => \N__33560\
        );

    \I__6596\ : LocalMux
    port map (
            O => \N__33560\,
            I => \current_shift_inst.un38_control_input_0_s1_28\
        );

    \I__6595\ : InMux
    port map (
            O => \N__33557\,
            I => \N__33554\
        );

    \I__6594\ : LocalMux
    port map (
            O => \N__33554\,
            I => \N__33551\
        );

    \I__6593\ : Span4Mux_h
    port map (
            O => \N__33551\,
            I => \N__33548\
        );

    \I__6592\ : Odrv4
    port map (
            O => \N__33548\,
            I => \current_shift_inst.control_input_axb_8\
        );

    \I__6591\ : InMux
    port map (
            O => \N__33545\,
            I => \N__33542\
        );

    \I__6590\ : LocalMux
    port map (
            O => \N__33542\,
            I => \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0\
        );

    \I__6589\ : CascadeMux
    port map (
            O => \N__33539\,
            I => \N__33536\
        );

    \I__6588\ : InMux
    port map (
            O => \N__33536\,
            I => \N__33533\
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__33533\,
            I => \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0\
        );

    \I__6586\ : CascadeMux
    port map (
            O => \N__33530\,
            I => \N__33527\
        );

    \I__6585\ : InMux
    port map (
            O => \N__33527\,
            I => \N__33524\
        );

    \I__6584\ : LocalMux
    port map (
            O => \N__33524\,
            I => \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0\
        );

    \I__6583\ : InMux
    port map (
            O => \N__33521\,
            I => \N__33518\
        );

    \I__6582\ : LocalMux
    port map (
            O => \N__33518\,
            I => \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0\
        );

    \I__6581\ : CascadeMux
    port map (
            O => \N__33515\,
            I => \N__33512\
        );

    \I__6580\ : InMux
    port map (
            O => \N__33512\,
            I => \N__33509\
        );

    \I__6579\ : LocalMux
    port map (
            O => \N__33509\,
            I => \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0\
        );

    \I__6578\ : CascadeMux
    port map (
            O => \N__33506\,
            I => \N__33503\
        );

    \I__6577\ : InMux
    port map (
            O => \N__33503\,
            I => \N__33500\
        );

    \I__6576\ : LocalMux
    port map (
            O => \N__33500\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\
        );

    \I__6575\ : InMux
    port map (
            O => \N__33497\,
            I => \N__33494\
        );

    \I__6574\ : LocalMux
    port map (
            O => \N__33494\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\
        );

    \I__6573\ : InMux
    port map (
            O => \N__33491\,
            I => \N__33488\
        );

    \I__6572\ : LocalMux
    port map (
            O => \N__33488\,
            I => \current_shift_inst.un38_control_input_0_s1_21\
        );

    \I__6571\ : InMux
    port map (
            O => \N__33485\,
            I => \N__33482\
        );

    \I__6570\ : LocalMux
    port map (
            O => \N__33482\,
            I => \N__33479\
        );

    \I__6569\ : Span4Mux_h
    port map (
            O => \N__33479\,
            I => \N__33476\
        );

    \I__6568\ : Odrv4
    port map (
            O => \N__33476\,
            I => \current_shift_inst.control_input_axb_1\
        );

    \I__6567\ : InMux
    port map (
            O => \N__33473\,
            I => \N__33470\
        );

    \I__6566\ : LocalMux
    port map (
            O => \N__33470\,
            I => \current_shift_inst.elapsed_time_ns_s1_fast_31\
        );

    \I__6565\ : CascadeMux
    port map (
            O => \N__33467\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\
        );

    \I__6564\ : CascadeMux
    port map (
            O => \N__33464\,
            I => \N__33460\
        );

    \I__6563\ : InMux
    port map (
            O => \N__33463\,
            I => \N__33457\
        );

    \I__6562\ : InMux
    port map (
            O => \N__33460\,
            I => \N__33454\
        );

    \I__6561\ : LocalMux
    port map (
            O => \N__33457\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__6560\ : LocalMux
    port map (
            O => \N__33454\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__6559\ : InMux
    port map (
            O => \N__33449\,
            I => \N__33446\
        );

    \I__6558\ : LocalMux
    port map (
            O => \N__33446\,
            I => \N__33440\
        );

    \I__6557\ : InMux
    port map (
            O => \N__33445\,
            I => \N__33437\
        );

    \I__6556\ : InMux
    port map (
            O => \N__33444\,
            I => \N__33432\
        );

    \I__6555\ : InMux
    port map (
            O => \N__33443\,
            I => \N__33432\
        );

    \I__6554\ : Span4Mux_h
    port map (
            O => \N__33440\,
            I => \N__33429\
        );

    \I__6553\ : LocalMux
    port map (
            O => \N__33437\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__6552\ : LocalMux
    port map (
            O => \N__33432\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__6551\ : Odrv4
    port map (
            O => \N__33429\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__6550\ : InMux
    port map (
            O => \N__33422\,
            I => \N__33384\
        );

    \I__6549\ : InMux
    port map (
            O => \N__33421\,
            I => \N__33384\
        );

    \I__6548\ : InMux
    port map (
            O => \N__33420\,
            I => \N__33384\
        );

    \I__6547\ : InMux
    port map (
            O => \N__33419\,
            I => \N__33384\
        );

    \I__6546\ : InMux
    port map (
            O => \N__33418\,
            I => \N__33375\
        );

    \I__6545\ : InMux
    port map (
            O => \N__33417\,
            I => \N__33375\
        );

    \I__6544\ : InMux
    port map (
            O => \N__33416\,
            I => \N__33375\
        );

    \I__6543\ : InMux
    port map (
            O => \N__33415\,
            I => \N__33375\
        );

    \I__6542\ : InMux
    port map (
            O => \N__33414\,
            I => \N__33370\
        );

    \I__6541\ : InMux
    port map (
            O => \N__33413\,
            I => \N__33370\
        );

    \I__6540\ : InMux
    port map (
            O => \N__33412\,
            I => \N__33361\
        );

    \I__6539\ : InMux
    port map (
            O => \N__33411\,
            I => \N__33361\
        );

    \I__6538\ : InMux
    port map (
            O => \N__33410\,
            I => \N__33361\
        );

    \I__6537\ : InMux
    port map (
            O => \N__33409\,
            I => \N__33361\
        );

    \I__6536\ : InMux
    port map (
            O => \N__33408\,
            I => \N__33352\
        );

    \I__6535\ : InMux
    port map (
            O => \N__33407\,
            I => \N__33352\
        );

    \I__6534\ : InMux
    port map (
            O => \N__33406\,
            I => \N__33352\
        );

    \I__6533\ : InMux
    port map (
            O => \N__33405\,
            I => \N__33352\
        );

    \I__6532\ : InMux
    port map (
            O => \N__33404\,
            I => \N__33343\
        );

    \I__6531\ : InMux
    port map (
            O => \N__33403\,
            I => \N__33343\
        );

    \I__6530\ : InMux
    port map (
            O => \N__33402\,
            I => \N__33343\
        );

    \I__6529\ : InMux
    port map (
            O => \N__33401\,
            I => \N__33343\
        );

    \I__6528\ : InMux
    port map (
            O => \N__33400\,
            I => \N__33334\
        );

    \I__6527\ : InMux
    port map (
            O => \N__33399\,
            I => \N__33334\
        );

    \I__6526\ : InMux
    port map (
            O => \N__33398\,
            I => \N__33334\
        );

    \I__6525\ : InMux
    port map (
            O => \N__33397\,
            I => \N__33334\
        );

    \I__6524\ : InMux
    port map (
            O => \N__33396\,
            I => \N__33325\
        );

    \I__6523\ : InMux
    port map (
            O => \N__33395\,
            I => \N__33325\
        );

    \I__6522\ : InMux
    port map (
            O => \N__33394\,
            I => \N__33325\
        );

    \I__6521\ : InMux
    port map (
            O => \N__33393\,
            I => \N__33325\
        );

    \I__6520\ : LocalMux
    port map (
            O => \N__33384\,
            I => \N__33322\
        );

    \I__6519\ : LocalMux
    port map (
            O => \N__33375\,
            I => \N__33319\
        );

    \I__6518\ : LocalMux
    port map (
            O => \N__33370\,
            I => \N__33314\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__33361\,
            I => \N__33314\
        );

    \I__6516\ : LocalMux
    port map (
            O => \N__33352\,
            I => \N__33305\
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__33343\,
            I => \N__33305\
        );

    \I__6514\ : LocalMux
    port map (
            O => \N__33334\,
            I => \N__33305\
        );

    \I__6513\ : LocalMux
    port map (
            O => \N__33325\,
            I => \N__33305\
        );

    \I__6512\ : Odrv4
    port map (
            O => \N__33322\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__6511\ : Odrv4
    port map (
            O => \N__33319\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__6510\ : Odrv4
    port map (
            O => \N__33314\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__6509\ : Odrv12
    port map (
            O => \N__33305\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__6508\ : InMux
    port map (
            O => \N__33296\,
            I => \N__33293\
        );

    \I__6507\ : LocalMux
    port map (
            O => \N__33293\,
            I => \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0\
        );

    \I__6506\ : CascadeMux
    port map (
            O => \N__33290\,
            I => \N__33287\
        );

    \I__6505\ : InMux
    port map (
            O => \N__33287\,
            I => \N__33284\
        );

    \I__6504\ : LocalMux
    port map (
            O => \N__33284\,
            I => \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0\
        );

    \I__6503\ : InMux
    port map (
            O => \N__33281\,
            I => \N__33278\
        );

    \I__6502\ : LocalMux
    port map (
            O => \N__33278\,
            I => \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0\
        );

    \I__6501\ : InMux
    port map (
            O => \N__33275\,
            I => \N__33272\
        );

    \I__6500\ : LocalMux
    port map (
            O => \N__33272\,
            I => \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0\
        );

    \I__6499\ : CascadeMux
    port map (
            O => \N__33269\,
            I => \N__33266\
        );

    \I__6498\ : InMux
    port map (
            O => \N__33266\,
            I => \N__33263\
        );

    \I__6497\ : LocalMux
    port map (
            O => \N__33263\,
            I => \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0\
        );

    \I__6496\ : InMux
    port map (
            O => \N__33260\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_24\
        );

    \I__6495\ : InMux
    port map (
            O => \N__33257\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_25\
        );

    \I__6494\ : InMux
    port map (
            O => \N__33254\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_26\
        );

    \I__6493\ : InMux
    port map (
            O => \N__33251\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_27\
        );

    \I__6492\ : InMux
    port map (
            O => \N__33248\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_28\
        );

    \I__6491\ : CEMux
    port map (
            O => \N__33245\,
            I => \N__33241\
        );

    \I__6490\ : CEMux
    port map (
            O => \N__33244\,
            I => \N__33238\
        );

    \I__6489\ : LocalMux
    port map (
            O => \N__33241\,
            I => \N__33233\
        );

    \I__6488\ : LocalMux
    port map (
            O => \N__33238\,
            I => \N__33230\
        );

    \I__6487\ : CEMux
    port map (
            O => \N__33237\,
            I => \N__33227\
        );

    \I__6486\ : CEMux
    port map (
            O => \N__33236\,
            I => \N__33224\
        );

    \I__6485\ : Span4Mux_v
    port map (
            O => \N__33233\,
            I => \N__33217\
        );

    \I__6484\ : Span4Mux_h
    port map (
            O => \N__33230\,
            I => \N__33217\
        );

    \I__6483\ : LocalMux
    port map (
            O => \N__33227\,
            I => \N__33217\
        );

    \I__6482\ : LocalMux
    port map (
            O => \N__33224\,
            I => \N__33214\
        );

    \I__6481\ : Span4Mux_v
    port map (
            O => \N__33217\,
            I => \N__33211\
        );

    \I__6480\ : Span4Mux_h
    port map (
            O => \N__33214\,
            I => \N__33208\
        );

    \I__6479\ : Odrv4
    port map (
            O => \N__33211\,
            I => \delay_measurement_inst.delay_tr_timer.N_205_i\
        );

    \I__6478\ : Odrv4
    port map (
            O => \N__33208\,
            I => \delay_measurement_inst.delay_tr_timer.N_205_i\
        );

    \I__6477\ : CascadeMux
    port map (
            O => \N__33203\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\
        );

    \I__6476\ : CascadeMux
    port map (
            O => \N__33200\,
            I => \N__33196\
        );

    \I__6475\ : InMux
    port map (
            O => \N__33199\,
            I => \N__33191\
        );

    \I__6474\ : InMux
    port map (
            O => \N__33196\,
            I => \N__33184\
        );

    \I__6473\ : InMux
    port map (
            O => \N__33195\,
            I => \N__33184\
        );

    \I__6472\ : InMux
    port map (
            O => \N__33194\,
            I => \N__33184\
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__33191\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__6470\ : LocalMux
    port map (
            O => \N__33184\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__6469\ : InMux
    port map (
            O => \N__33179\,
            I => \N__33176\
        );

    \I__6468\ : LocalMux
    port map (
            O => \N__33176\,
            I => \current_shift_inst.un4_control_input1_1\
        );

    \I__6467\ : InMux
    port map (
            O => \N__33173\,
            I => \bfn_13_12_0_\
        );

    \I__6466\ : InMux
    port map (
            O => \N__33170\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_16\
        );

    \I__6465\ : InMux
    port map (
            O => \N__33167\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_17\
        );

    \I__6464\ : InMux
    port map (
            O => \N__33164\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_18\
        );

    \I__6463\ : InMux
    port map (
            O => \N__33161\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_19\
        );

    \I__6462\ : InMux
    port map (
            O => \N__33158\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_20\
        );

    \I__6461\ : InMux
    port map (
            O => \N__33155\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_21\
        );

    \I__6460\ : InMux
    port map (
            O => \N__33152\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_22\
        );

    \I__6459\ : InMux
    port map (
            O => \N__33149\,
            I => \bfn_13_13_0_\
        );

    \I__6458\ : InMux
    port map (
            O => \N__33146\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_6\
        );

    \I__6457\ : InMux
    port map (
            O => \N__33143\,
            I => \bfn_13_11_0_\
        );

    \I__6456\ : InMux
    port map (
            O => \N__33140\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_8\
        );

    \I__6455\ : InMux
    port map (
            O => \N__33137\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_9\
        );

    \I__6454\ : InMux
    port map (
            O => \N__33134\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_10\
        );

    \I__6453\ : InMux
    port map (
            O => \N__33131\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_11\
        );

    \I__6452\ : InMux
    port map (
            O => \N__33128\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_12\
        );

    \I__6451\ : InMux
    port map (
            O => \N__33125\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_13\
        );

    \I__6450\ : InMux
    port map (
            O => \N__33122\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_14\
        );

    \I__6449\ : CascadeMux
    port map (
            O => \N__33119\,
            I => \N__33115\
        );

    \I__6448\ : InMux
    port map (
            O => \N__33118\,
            I => \N__33107\
        );

    \I__6447\ : InMux
    port map (
            O => \N__33115\,
            I => \N__33107\
        );

    \I__6446\ : InMux
    port map (
            O => \N__33114\,
            I => \N__33107\
        );

    \I__6445\ : LocalMux
    port map (
            O => \N__33107\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_31\
        );

    \I__6444\ : InMux
    port map (
            O => \N__33104\,
            I => \bfn_13_10_0_\
        );

    \I__6443\ : InMux
    port map (
            O => \N__33101\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_0\
        );

    \I__6442\ : InMux
    port map (
            O => \N__33098\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_1\
        );

    \I__6441\ : InMux
    port map (
            O => \N__33095\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_2\
        );

    \I__6440\ : InMux
    port map (
            O => \N__33092\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_3\
        );

    \I__6439\ : InMux
    port map (
            O => \N__33089\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_4\
        );

    \I__6438\ : InMux
    port map (
            O => \N__33086\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_5\
        );

    \I__6437\ : CascadeMux
    port map (
            O => \N__33083\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\
        );

    \I__6436\ : InMux
    port map (
            O => \N__33080\,
            I => \N__33073\
        );

    \I__6435\ : InMux
    port map (
            O => \N__33079\,
            I => \N__33068\
        );

    \I__6434\ : InMux
    port map (
            O => \N__33078\,
            I => \N__33068\
        );

    \I__6433\ : InMux
    port map (
            O => \N__33077\,
            I => \N__33065\
        );

    \I__6432\ : InMux
    port map (
            O => \N__33076\,
            I => \N__33062\
        );

    \I__6431\ : LocalMux
    port map (
            O => \N__33073\,
            I => \N__33057\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__33068\,
            I => \N__33057\
        );

    \I__6429\ : LocalMux
    port map (
            O => \N__33065\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__6428\ : LocalMux
    port map (
            O => \N__33062\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__6427\ : Odrv4
    port map (
            O => \N__33057\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__6426\ : InMux
    port map (
            O => \N__33050\,
            I => \N__33046\
        );

    \I__6425\ : InMux
    port map (
            O => \N__33049\,
            I => \N__33043\
        );

    \I__6424\ : LocalMux
    port map (
            O => \N__33046\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\
        );

    \I__6423\ : LocalMux
    port map (
            O => \N__33043\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\
        );

    \I__6422\ : CascadeMux
    port map (
            O => \N__33038\,
            I => \N__33035\
        );

    \I__6421\ : InMux
    port map (
            O => \N__33035\,
            I => \N__33032\
        );

    \I__6420\ : LocalMux
    port map (
            O => \N__33032\,
            I => \N__33029\
        );

    \I__6419\ : Odrv4
    port map (
            O => \N__33029\,
            I => \phase_controller_inst2.stoper_tr.un4_running_df30\
        );

    \I__6418\ : InMux
    port map (
            O => \N__33026\,
            I => \N__33017\
        );

    \I__6417\ : InMux
    port map (
            O => \N__33025\,
            I => \N__33017\
        );

    \I__6416\ : InMux
    port map (
            O => \N__33024\,
            I => \N__33017\
        );

    \I__6415\ : LocalMux
    port map (
            O => \N__33017\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_30\
        );

    \I__6414\ : CascadeMux
    port map (
            O => \N__33014\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13_cascade_\
        );

    \I__6413\ : InMux
    port map (
            O => \N__33011\,
            I => \N__33007\
        );

    \I__6412\ : CascadeMux
    port map (
            O => \N__33010\,
            I => \N__33004\
        );

    \I__6411\ : LocalMux
    port map (
            O => \N__33007\,
            I => \N__32999\
        );

    \I__6410\ : InMux
    port map (
            O => \N__33004\,
            I => \N__32996\
        );

    \I__6409\ : InMux
    port map (
            O => \N__33003\,
            I => \N__32991\
        );

    \I__6408\ : InMux
    port map (
            O => \N__33002\,
            I => \N__32991\
        );

    \I__6407\ : Span12Mux_v
    port map (
            O => \N__32999\,
            I => \N__32988\
        );

    \I__6406\ : LocalMux
    port map (
            O => \N__32996\,
            I => \N__32985\
        );

    \I__6405\ : LocalMux
    port map (
            O => \N__32991\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__6404\ : Odrv12
    port map (
            O => \N__32988\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__6403\ : Odrv4
    port map (
            O => \N__32985\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__6402\ : IoInMux
    port map (
            O => \N__32978\,
            I => \N__32975\
        );

    \I__6401\ : LocalMux
    port map (
            O => \N__32975\,
            I => \N__32972\
        );

    \I__6400\ : IoSpan4Mux
    port map (
            O => \N__32972\,
            I => \N__32969\
        );

    \I__6399\ : Sp12to4
    port map (
            O => \N__32969\,
            I => \N__32966\
        );

    \I__6398\ : Odrv12
    port map (
            O => \N__32966\,
            I => s4_phy_c
        );

    \I__6397\ : InMux
    port map (
            O => \N__32963\,
            I => \N__32960\
        );

    \I__6396\ : LocalMux
    port map (
            O => \N__32960\,
            I => \N__32956\
        );

    \I__6395\ : InMux
    port map (
            O => \N__32959\,
            I => \N__32953\
        );

    \I__6394\ : Span4Mux_h
    port map (
            O => \N__32956\,
            I => \N__32948\
        );

    \I__6393\ : LocalMux
    port map (
            O => \N__32953\,
            I => \N__32948\
        );

    \I__6392\ : Span4Mux_h
    port map (
            O => \N__32948\,
            I => \N__32943\
        );

    \I__6391\ : InMux
    port map (
            O => \N__32947\,
            I => \N__32940\
        );

    \I__6390\ : InMux
    port map (
            O => \N__32946\,
            I => \N__32937\
        );

    \I__6389\ : Span4Mux_v
    port map (
            O => \N__32943\,
            I => \N__32934\
        );

    \I__6388\ : LocalMux
    port map (
            O => \N__32940\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__6387\ : LocalMux
    port map (
            O => \N__32937\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__6386\ : Odrv4
    port map (
            O => \N__32934\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__6385\ : ClkMux
    port map (
            O => \N__32927\,
            I => \N__32921\
        );

    \I__6384\ : ClkMux
    port map (
            O => \N__32926\,
            I => \N__32921\
        );

    \I__6383\ : GlobalMux
    port map (
            O => \N__32921\,
            I => \N__32918\
        );

    \I__6382\ : gio2CtrlBuf
    port map (
            O => \N__32918\,
            I => delay_hc_input_c_g
        );

    \I__6381\ : IoInMux
    port map (
            O => \N__32915\,
            I => \N__32912\
        );

    \I__6380\ : LocalMux
    port map (
            O => \N__32912\,
            I => \N__32909\
        );

    \I__6379\ : Span4Mux_s0_v
    port map (
            O => \N__32909\,
            I => \N__32906\
        );

    \I__6378\ : Odrv4
    port map (
            O => \N__32906\,
            I => \pll_inst.red_c_i\
        );

    \I__6377\ : InMux
    port map (
            O => \N__32903\,
            I => \N__32899\
        );

    \I__6376\ : InMux
    port map (
            O => \N__32902\,
            I => \N__32896\
        );

    \I__6375\ : LocalMux
    port map (
            O => \N__32899\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__6374\ : LocalMux
    port map (
            O => \N__32896\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__6373\ : InMux
    port map (
            O => \N__32891\,
            I => \N__32887\
        );

    \I__6372\ : InMux
    port map (
            O => \N__32890\,
            I => \N__32884\
        );

    \I__6371\ : LocalMux
    port map (
            O => \N__32887\,
            I => \phase_controller_inst2.state_RNI9M3OZ0Z_0\
        );

    \I__6370\ : LocalMux
    port map (
            O => \N__32884\,
            I => \phase_controller_inst2.state_RNI9M3OZ0Z_0\
        );

    \I__6369\ : InMux
    port map (
            O => \N__32879\,
            I => \N__32875\
        );

    \I__6368\ : CascadeMux
    port map (
            O => \N__32878\,
            I => \N__32872\
        );

    \I__6367\ : LocalMux
    port map (
            O => \N__32875\,
            I => \N__32867\
        );

    \I__6366\ : InMux
    port map (
            O => \N__32872\,
            I => \N__32864\
        );

    \I__6365\ : InMux
    port map (
            O => \N__32871\,
            I => \N__32859\
        );

    \I__6364\ : InMux
    port map (
            O => \N__32870\,
            I => \N__32859\
        );

    \I__6363\ : Odrv4
    port map (
            O => \N__32867\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__6362\ : LocalMux
    port map (
            O => \N__32864\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__6361\ : LocalMux
    port map (
            O => \N__32859\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__6360\ : CascadeMux
    port map (
            O => \N__32852\,
            I => \N__32848\
        );

    \I__6359\ : InMux
    port map (
            O => \N__32851\,
            I => \N__32844\
        );

    \I__6358\ : InMux
    port map (
            O => \N__32848\,
            I => \N__32841\
        );

    \I__6357\ : InMux
    port map (
            O => \N__32847\,
            I => \N__32838\
        );

    \I__6356\ : LocalMux
    port map (
            O => \N__32844\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__6355\ : LocalMux
    port map (
            O => \N__32841\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__6354\ : LocalMux
    port map (
            O => \N__32838\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__6353\ : CascadeMux
    port map (
            O => \N__32831\,
            I => \N__32827\
        );

    \I__6352\ : InMux
    port map (
            O => \N__32830\,
            I => \N__32824\
        );

    \I__6351\ : InMux
    port map (
            O => \N__32827\,
            I => \N__32821\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__32824\,
            I => \N__32818\
        );

    \I__6349\ : LocalMux
    port map (
            O => \N__32821\,
            I => \phase_controller_inst2.stoper_tr.runningZ0\
        );

    \I__6348\ : Odrv4
    port map (
            O => \N__32818\,
            I => \phase_controller_inst2.stoper_tr.runningZ0\
        );

    \I__6347\ : CascadeMux
    port map (
            O => \N__32813\,
            I => \N__32808\
        );

    \I__6346\ : InMux
    port map (
            O => \N__32812\,
            I => \N__32803\
        );

    \I__6345\ : InMux
    port map (
            O => \N__32811\,
            I => \N__32803\
        );

    \I__6344\ : InMux
    port map (
            O => \N__32808\,
            I => \N__32798\
        );

    \I__6343\ : LocalMux
    port map (
            O => \N__32803\,
            I => \N__32795\
        );

    \I__6342\ : InMux
    port map (
            O => \N__32802\,
            I => \N__32790\
        );

    \I__6341\ : InMux
    port map (
            O => \N__32801\,
            I => \N__32790\
        );

    \I__6340\ : LocalMux
    port map (
            O => \N__32798\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__6339\ : Odrv4
    port map (
            O => \N__32795\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__6338\ : LocalMux
    port map (
            O => \N__32790\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__6337\ : InMux
    port map (
            O => \N__32783\,
            I => \N__32780\
        );

    \I__6336\ : LocalMux
    port map (
            O => \N__32780\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\
        );

    \I__6335\ : InMux
    port map (
            O => \N__32777\,
            I => \current_shift_inst.un38_control_input_cry_24_s1\
        );

    \I__6334\ : InMux
    port map (
            O => \N__32774\,
            I => \current_shift_inst.un38_control_input_cry_25_s1\
        );

    \I__6333\ : InMux
    port map (
            O => \N__32771\,
            I => \current_shift_inst.un38_control_input_cry_26_s1\
        );

    \I__6332\ : InMux
    port map (
            O => \N__32768\,
            I => \current_shift_inst.un38_control_input_cry_27_s1\
        );

    \I__6331\ : InMux
    port map (
            O => \N__32765\,
            I => \current_shift_inst.un38_control_input_cry_28_s1\
        );

    \I__6330\ : InMux
    port map (
            O => \N__32762\,
            I => \current_shift_inst.un38_control_input_cry_29_s1\
        );

    \I__6329\ : InMux
    port map (
            O => \N__32759\,
            I => \current_shift_inst.un38_control_input_cry_30_s1\
        );

    \I__6328\ : InMux
    port map (
            O => \N__32756\,
            I => \N__32753\
        );

    \I__6327\ : LocalMux
    port map (
            O => \N__32753\,
            I => \N__32750\
        );

    \I__6326\ : Span4Mux_v
    port map (
            O => \N__32750\,
            I => \N__32747\
        );

    \I__6325\ : Span4Mux_h
    port map (
            O => \N__32747\,
            I => \N__32744\
        );

    \I__6324\ : Sp12to4
    port map (
            O => \N__32744\,
            I => \N__32741\
        );

    \I__6323\ : Span12Mux_v
    port map (
            O => \N__32741\,
            I => \N__32738\
        );

    \I__6322\ : Odrv12
    port map (
            O => \N__32738\,
            I => il_min_comp1_c
        );

    \I__6321\ : InMux
    port map (
            O => \N__32735\,
            I => \N__32732\
        );

    \I__6320\ : LocalMux
    port map (
            O => \N__32732\,
            I => \il_min_comp1_D1\
        );

    \I__6319\ : InMux
    port map (
            O => \N__32729\,
            I => \N__32726\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__32726\,
            I => \N__32723\
        );

    \I__6317\ : Odrv4
    port map (
            O => \N__32723\,
            I => \current_shift_inst.un38_control_input_0_s1_20\
        );

    \I__6316\ : InMux
    port map (
            O => \N__32720\,
            I => \current_shift_inst.un38_control_input_cry_19_s1\
        );

    \I__6315\ : InMux
    port map (
            O => \N__32717\,
            I => \current_shift_inst.un38_control_input_cry_20_s1\
        );

    \I__6314\ : CascadeMux
    port map (
            O => \N__32714\,
            I => \N__32711\
        );

    \I__6313\ : InMux
    port map (
            O => \N__32711\,
            I => \N__32708\
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__32708\,
            I => \N__32705\
        );

    \I__6311\ : Odrv4
    port map (
            O => \N__32705\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\
        );

    \I__6310\ : InMux
    port map (
            O => \N__32702\,
            I => \current_shift_inst.un38_control_input_cry_21_s1\
        );

    \I__6309\ : InMux
    port map (
            O => \N__32699\,
            I => \current_shift_inst.un38_control_input_cry_22_s1\
        );

    \I__6308\ : InMux
    port map (
            O => \N__32696\,
            I => \bfn_12_18_0_\
        );

    \I__6307\ : CascadeMux
    port map (
            O => \N__32693\,
            I => \N__32690\
        );

    \I__6306\ : InMux
    port map (
            O => \N__32690\,
            I => \N__32687\
        );

    \I__6305\ : LocalMux
    port map (
            O => \N__32687\,
            I => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\
        );

    \I__6304\ : InMux
    port map (
            O => \N__32684\,
            I => \N__32681\
        );

    \I__6303\ : LocalMux
    port map (
            O => \N__32681\,
            I => \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\
        );

    \I__6302\ : InMux
    port map (
            O => \N__32678\,
            I => \N__32675\
        );

    \I__6301\ : LocalMux
    port map (
            O => \N__32675\,
            I => \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0\
        );

    \I__6300\ : CEMux
    port map (
            O => \N__32672\,
            I => \N__32649\
        );

    \I__6299\ : CEMux
    port map (
            O => \N__32671\,
            I => \N__32644\
        );

    \I__6298\ : InMux
    port map (
            O => \N__32670\,
            I => \N__32635\
        );

    \I__6297\ : InMux
    port map (
            O => \N__32669\,
            I => \N__32635\
        );

    \I__6296\ : InMux
    port map (
            O => \N__32668\,
            I => \N__32635\
        );

    \I__6295\ : InMux
    port map (
            O => \N__32667\,
            I => \N__32635\
        );

    \I__6294\ : InMux
    port map (
            O => \N__32666\,
            I => \N__32626\
        );

    \I__6293\ : InMux
    port map (
            O => \N__32665\,
            I => \N__32626\
        );

    \I__6292\ : InMux
    port map (
            O => \N__32664\,
            I => \N__32626\
        );

    \I__6291\ : InMux
    port map (
            O => \N__32663\,
            I => \N__32626\
        );

    \I__6290\ : InMux
    port map (
            O => \N__32662\,
            I => \N__32617\
        );

    \I__6289\ : InMux
    port map (
            O => \N__32661\,
            I => \N__32617\
        );

    \I__6288\ : InMux
    port map (
            O => \N__32660\,
            I => \N__32617\
        );

    \I__6287\ : InMux
    port map (
            O => \N__32659\,
            I => \N__32617\
        );

    \I__6286\ : CEMux
    port map (
            O => \N__32658\,
            I => \N__32613\
        );

    \I__6285\ : CEMux
    port map (
            O => \N__32657\,
            I => \N__32602\
        );

    \I__6284\ : CEMux
    port map (
            O => \N__32656\,
            I => \N__32595\
        );

    \I__6283\ : CEMux
    port map (
            O => \N__32655\,
            I => \N__32591\
        );

    \I__6282\ : CEMux
    port map (
            O => \N__32654\,
            I => \N__32587\
        );

    \I__6281\ : CEMux
    port map (
            O => \N__32653\,
            I => \N__32584\
        );

    \I__6280\ : CEMux
    port map (
            O => \N__32652\,
            I => \N__32581\
        );

    \I__6279\ : LocalMux
    port map (
            O => \N__32649\,
            I => \N__32578\
        );

    \I__6278\ : CEMux
    port map (
            O => \N__32648\,
            I => \N__32575\
        );

    \I__6277\ : CEMux
    port map (
            O => \N__32647\,
            I => \N__32568\
        );

    \I__6276\ : LocalMux
    port map (
            O => \N__32644\,
            I => \N__32559\
        );

    \I__6275\ : LocalMux
    port map (
            O => \N__32635\,
            I => \N__32559\
        );

    \I__6274\ : LocalMux
    port map (
            O => \N__32626\,
            I => \N__32559\
        );

    \I__6273\ : LocalMux
    port map (
            O => \N__32617\,
            I => \N__32559\
        );

    \I__6272\ : CEMux
    port map (
            O => \N__32616\,
            I => \N__32556\
        );

    \I__6271\ : LocalMux
    port map (
            O => \N__32613\,
            I => \N__32549\
        );

    \I__6270\ : InMux
    port map (
            O => \N__32612\,
            I => \N__32540\
        );

    \I__6269\ : InMux
    port map (
            O => \N__32611\,
            I => \N__32540\
        );

    \I__6268\ : InMux
    port map (
            O => \N__32610\,
            I => \N__32540\
        );

    \I__6267\ : InMux
    port map (
            O => \N__32609\,
            I => \N__32540\
        );

    \I__6266\ : InMux
    port map (
            O => \N__32608\,
            I => \N__32531\
        );

    \I__6265\ : InMux
    port map (
            O => \N__32607\,
            I => \N__32531\
        );

    \I__6264\ : InMux
    port map (
            O => \N__32606\,
            I => \N__32531\
        );

    \I__6263\ : InMux
    port map (
            O => \N__32605\,
            I => \N__32531\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__32602\,
            I => \N__32528\
        );

    \I__6261\ : CEMux
    port map (
            O => \N__32601\,
            I => \N__32525\
        );

    \I__6260\ : InMux
    port map (
            O => \N__32600\,
            I => \N__32518\
        );

    \I__6259\ : InMux
    port map (
            O => \N__32599\,
            I => \N__32518\
        );

    \I__6258\ : InMux
    port map (
            O => \N__32598\,
            I => \N__32518\
        );

    \I__6257\ : LocalMux
    port map (
            O => \N__32595\,
            I => \N__32515\
        );

    \I__6256\ : CEMux
    port map (
            O => \N__32594\,
            I => \N__32512\
        );

    \I__6255\ : LocalMux
    port map (
            O => \N__32591\,
            I => \N__32509\
        );

    \I__6254\ : CEMux
    port map (
            O => \N__32590\,
            I => \N__32506\
        );

    \I__6253\ : LocalMux
    port map (
            O => \N__32587\,
            I => \N__32503\
        );

    \I__6252\ : LocalMux
    port map (
            O => \N__32584\,
            I => \N__32498\
        );

    \I__6251\ : LocalMux
    port map (
            O => \N__32581\,
            I => \N__32498\
        );

    \I__6250\ : Span4Mux_s3_v
    port map (
            O => \N__32578\,
            I => \N__32492\
        );

    \I__6249\ : LocalMux
    port map (
            O => \N__32575\,
            I => \N__32492\
        );

    \I__6248\ : CEMux
    port map (
            O => \N__32574\,
            I => \N__32489\
        );

    \I__6247\ : InMux
    port map (
            O => \N__32573\,
            I => \N__32482\
        );

    \I__6246\ : InMux
    port map (
            O => \N__32572\,
            I => \N__32482\
        );

    \I__6245\ : InMux
    port map (
            O => \N__32571\,
            I => \N__32482\
        );

    \I__6244\ : LocalMux
    port map (
            O => \N__32568\,
            I => \N__32475\
        );

    \I__6243\ : Span4Mux_v
    port map (
            O => \N__32559\,
            I => \N__32475\
        );

    \I__6242\ : LocalMux
    port map (
            O => \N__32556\,
            I => \N__32475\
        );

    \I__6241\ : InMux
    port map (
            O => \N__32555\,
            I => \N__32466\
        );

    \I__6240\ : InMux
    port map (
            O => \N__32554\,
            I => \N__32466\
        );

    \I__6239\ : InMux
    port map (
            O => \N__32553\,
            I => \N__32466\
        );

    \I__6238\ : InMux
    port map (
            O => \N__32552\,
            I => \N__32466\
        );

    \I__6237\ : Span4Mux_h
    port map (
            O => \N__32549\,
            I => \N__32453\
        );

    \I__6236\ : LocalMux
    port map (
            O => \N__32540\,
            I => \N__32453\
        );

    \I__6235\ : LocalMux
    port map (
            O => \N__32531\,
            I => \N__32453\
        );

    \I__6234\ : Span4Mux_s3_v
    port map (
            O => \N__32528\,
            I => \N__32453\
        );

    \I__6233\ : LocalMux
    port map (
            O => \N__32525\,
            I => \N__32453\
        );

    \I__6232\ : LocalMux
    port map (
            O => \N__32518\,
            I => \N__32453\
        );

    \I__6231\ : Span4Mux_v
    port map (
            O => \N__32515\,
            I => \N__32448\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__32512\,
            I => \N__32448\
        );

    \I__6229\ : Span4Mux_v
    port map (
            O => \N__32509\,
            I => \N__32443\
        );

    \I__6228\ : LocalMux
    port map (
            O => \N__32506\,
            I => \N__32443\
        );

    \I__6227\ : Span4Mux_v
    port map (
            O => \N__32503\,
            I => \N__32438\
        );

    \I__6226\ : Span4Mux_v
    port map (
            O => \N__32498\,
            I => \N__32438\
        );

    \I__6225\ : InMux
    port map (
            O => \N__32497\,
            I => \N__32435\
        );

    \I__6224\ : Span4Mux_v
    port map (
            O => \N__32492\,
            I => \N__32432\
        );

    \I__6223\ : LocalMux
    port map (
            O => \N__32489\,
            I => \N__32419\
        );

    \I__6222\ : LocalMux
    port map (
            O => \N__32482\,
            I => \N__32419\
        );

    \I__6221\ : Span4Mux_v
    port map (
            O => \N__32475\,
            I => \N__32419\
        );

    \I__6220\ : LocalMux
    port map (
            O => \N__32466\,
            I => \N__32419\
        );

    \I__6219\ : Span4Mux_v
    port map (
            O => \N__32453\,
            I => \N__32419\
        );

    \I__6218\ : Span4Mux_h
    port map (
            O => \N__32448\,
            I => \N__32419\
        );

    \I__6217\ : Sp12to4
    port map (
            O => \N__32443\,
            I => \N__32412\
        );

    \I__6216\ : Sp12to4
    port map (
            O => \N__32438\,
            I => \N__32412\
        );

    \I__6215\ : LocalMux
    port map (
            O => \N__32435\,
            I => \N__32412\
        );

    \I__6214\ : Span4Mux_h
    port map (
            O => \N__32432\,
            I => \N__32409\
        );

    \I__6213\ : Span4Mux_h
    port map (
            O => \N__32419\,
            I => \N__32406\
        );

    \I__6212\ : Odrv12
    port map (
            O => \N__32412\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__6211\ : Odrv4
    port map (
            O => \N__32409\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__6210\ : Odrv4
    port map (
            O => \N__32406\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__6209\ : InMux
    port map (
            O => \N__32399\,
            I => \N__32396\
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__32396\,
            I => \N__32392\
        );

    \I__6207\ : InMux
    port map (
            O => \N__32395\,
            I => \N__32389\
        );

    \I__6206\ : Odrv12
    port map (
            O => \N__32392\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\
        );

    \I__6205\ : LocalMux
    port map (
            O => \N__32389\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\
        );

    \I__6204\ : CascadeMux
    port map (
            O => \N__32384\,
            I => \N__32381\
        );

    \I__6203\ : InMux
    port map (
            O => \N__32381\,
            I => \N__32378\
        );

    \I__6202\ : LocalMux
    port map (
            O => \N__32378\,
            I => \N__32374\
        );

    \I__6201\ : CascadeMux
    port map (
            O => \N__32377\,
            I => \N__32369\
        );

    \I__6200\ : Span4Mux_h
    port map (
            O => \N__32374\,
            I => \N__32365\
        );

    \I__6199\ : InMux
    port map (
            O => \N__32373\,
            I => \N__32360\
        );

    \I__6198\ : InMux
    port map (
            O => \N__32372\,
            I => \N__32360\
        );

    \I__6197\ : InMux
    port map (
            O => \N__32369\,
            I => \N__32357\
        );

    \I__6196\ : InMux
    port map (
            O => \N__32368\,
            I => \N__32354\
        );

    \I__6195\ : Span4Mux_h
    port map (
            O => \N__32365\,
            I => \N__32349\
        );

    \I__6194\ : LocalMux
    port map (
            O => \N__32360\,
            I => \N__32349\
        );

    \I__6193\ : LocalMux
    port map (
            O => \N__32357\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__6192\ : LocalMux
    port map (
            O => \N__32354\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__6191\ : Odrv4
    port map (
            O => \N__32349\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__6190\ : CascadeMux
    port map (
            O => \N__32342\,
            I => \N__32339\
        );

    \I__6189\ : InMux
    port map (
            O => \N__32339\,
            I => \N__32336\
        );

    \I__6188\ : LocalMux
    port map (
            O => \N__32336\,
            I => \N__32332\
        );

    \I__6187\ : InMux
    port map (
            O => \N__32335\,
            I => \N__32329\
        );

    \I__6186\ : Span4Mux_v
    port map (
            O => \N__32332\,
            I => \N__32323\
        );

    \I__6185\ : LocalMux
    port map (
            O => \N__32329\,
            I => \N__32323\
        );

    \I__6184\ : InMux
    port map (
            O => \N__32328\,
            I => \N__32320\
        );

    \I__6183\ : Span4Mux_v
    port map (
            O => \N__32323\,
            I => \N__32317\
        );

    \I__6182\ : LocalMux
    port map (
            O => \N__32320\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__6181\ : Odrv4
    port map (
            O => \N__32317\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__6180\ : CascadeMux
    port map (
            O => \N__32312\,
            I => \N__32309\
        );

    \I__6179\ : InMux
    port map (
            O => \N__32309\,
            I => \N__32305\
        );

    \I__6178\ : InMux
    port map (
            O => \N__32308\,
            I => \N__32302\
        );

    \I__6177\ : LocalMux
    port map (
            O => \N__32305\,
            I => \phase_controller_inst2.stoper_hc.runningZ0\
        );

    \I__6176\ : LocalMux
    port map (
            O => \N__32302\,
            I => \phase_controller_inst2.stoper_hc.runningZ0\
        );

    \I__6175\ : InMux
    port map (
            O => \N__32297\,
            I => \N__32287\
        );

    \I__6174\ : InMux
    port map (
            O => \N__32296\,
            I => \N__32287\
        );

    \I__6173\ : InMux
    port map (
            O => \N__32295\,
            I => \N__32287\
        );

    \I__6172\ : CascadeMux
    port map (
            O => \N__32294\,
            I => \N__32283\
        );

    \I__6171\ : LocalMux
    port map (
            O => \N__32287\,
            I => \N__32280\
        );

    \I__6170\ : InMux
    port map (
            O => \N__32286\,
            I => \N__32275\
        );

    \I__6169\ : InMux
    port map (
            O => \N__32283\,
            I => \N__32275\
        );

    \I__6168\ : Span4Mux_h
    port map (
            O => \N__32280\,
            I => \N__32272\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__32275\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__6166\ : Odrv4
    port map (
            O => \N__32272\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__6165\ : InMux
    port map (
            O => \N__32267\,
            I => \N__32263\
        );

    \I__6164\ : InMux
    port map (
            O => \N__32266\,
            I => \N__32258\
        );

    \I__6163\ : LocalMux
    port map (
            O => \N__32263\,
            I => \N__32255\
        );

    \I__6162\ : InMux
    port map (
            O => \N__32262\,
            I => \N__32252\
        );

    \I__6161\ : CascadeMux
    port map (
            O => \N__32261\,
            I => \N__32249\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__32258\,
            I => \N__32242\
        );

    \I__6159\ : Span4Mux_v
    port map (
            O => \N__32255\,
            I => \N__32242\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__32252\,
            I => \N__32242\
        );

    \I__6157\ : InMux
    port map (
            O => \N__32249\,
            I => \N__32239\
        );

    \I__6156\ : Span4Mux_v
    port map (
            O => \N__32242\,
            I => \N__32236\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__32239\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__6154\ : Odrv4
    port map (
            O => \N__32236\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__6153\ : InMux
    port map (
            O => \N__32231\,
            I => \N__32225\
        );

    \I__6152\ : InMux
    port map (
            O => \N__32230\,
            I => \N__32222\
        );

    \I__6151\ : InMux
    port map (
            O => \N__32229\,
            I => \N__32216\
        );

    \I__6150\ : InMux
    port map (
            O => \N__32228\,
            I => \N__32216\
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__32225\,
            I => \N__32213\
        );

    \I__6148\ : LocalMux
    port map (
            O => \N__32222\,
            I => \N__32210\
        );

    \I__6147\ : InMux
    port map (
            O => \N__32221\,
            I => \N__32207\
        );

    \I__6146\ : LocalMux
    port map (
            O => \N__32216\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__6145\ : Odrv12
    port map (
            O => \N__32213\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__6144\ : Odrv4
    port map (
            O => \N__32210\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__6143\ : LocalMux
    port map (
            O => \N__32207\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__6142\ : IoInMux
    port map (
            O => \N__32198\,
            I => \N__32195\
        );

    \I__6141\ : LocalMux
    port map (
            O => \N__32195\,
            I => \N__32192\
        );

    \I__6140\ : Span4Mux_s1_v
    port map (
            O => \N__32192\,
            I => \N__32169\
        );

    \I__6139\ : InMux
    port map (
            O => \N__32191\,
            I => \N__32156\
        );

    \I__6138\ : InMux
    port map (
            O => \N__32190\,
            I => \N__32156\
        );

    \I__6137\ : InMux
    port map (
            O => \N__32189\,
            I => \N__32156\
        );

    \I__6136\ : InMux
    port map (
            O => \N__32188\,
            I => \N__32156\
        );

    \I__6135\ : InMux
    port map (
            O => \N__32187\,
            I => \N__32147\
        );

    \I__6134\ : InMux
    port map (
            O => \N__32186\,
            I => \N__32147\
        );

    \I__6133\ : InMux
    port map (
            O => \N__32185\,
            I => \N__32147\
        );

    \I__6132\ : InMux
    port map (
            O => \N__32184\,
            I => \N__32147\
        );

    \I__6131\ : InMux
    port map (
            O => \N__32183\,
            I => \N__32140\
        );

    \I__6130\ : InMux
    port map (
            O => \N__32182\,
            I => \N__32140\
        );

    \I__6129\ : InMux
    port map (
            O => \N__32181\,
            I => \N__32140\
        );

    \I__6128\ : InMux
    port map (
            O => \N__32180\,
            I => \N__32131\
        );

    \I__6127\ : InMux
    port map (
            O => \N__32179\,
            I => \N__32131\
        );

    \I__6126\ : InMux
    port map (
            O => \N__32178\,
            I => \N__32131\
        );

    \I__6125\ : InMux
    port map (
            O => \N__32177\,
            I => \N__32131\
        );

    \I__6124\ : InMux
    port map (
            O => \N__32176\,
            I => \N__32122\
        );

    \I__6123\ : InMux
    port map (
            O => \N__32175\,
            I => \N__32122\
        );

    \I__6122\ : InMux
    port map (
            O => \N__32174\,
            I => \N__32122\
        );

    \I__6121\ : InMux
    port map (
            O => \N__32173\,
            I => \N__32122\
        );

    \I__6120\ : InMux
    port map (
            O => \N__32172\,
            I => \N__32119\
        );

    \I__6119\ : Sp12to4
    port map (
            O => \N__32169\,
            I => \N__32116\
        );

    \I__6118\ : InMux
    port map (
            O => \N__32168\,
            I => \N__32100\
        );

    \I__6117\ : InMux
    port map (
            O => \N__32167\,
            I => \N__32100\
        );

    \I__6116\ : InMux
    port map (
            O => \N__32166\,
            I => \N__32100\
        );

    \I__6115\ : InMux
    port map (
            O => \N__32165\,
            I => \N__32100\
        );

    \I__6114\ : LocalMux
    port map (
            O => \N__32156\,
            I => \N__32097\
        );

    \I__6113\ : LocalMux
    port map (
            O => \N__32147\,
            I => \N__32086\
        );

    \I__6112\ : LocalMux
    port map (
            O => \N__32140\,
            I => \N__32086\
        );

    \I__6111\ : LocalMux
    port map (
            O => \N__32131\,
            I => \N__32086\
        );

    \I__6110\ : LocalMux
    port map (
            O => \N__32122\,
            I => \N__32086\
        );

    \I__6109\ : LocalMux
    port map (
            O => \N__32119\,
            I => \N__32086\
        );

    \I__6108\ : Span12Mux_h
    port map (
            O => \N__32116\,
            I => \N__32083\
        );

    \I__6107\ : InMux
    port map (
            O => \N__32115\,
            I => \N__32076\
        );

    \I__6106\ : InMux
    port map (
            O => \N__32114\,
            I => \N__32076\
        );

    \I__6105\ : InMux
    port map (
            O => \N__32113\,
            I => \N__32076\
        );

    \I__6104\ : InMux
    port map (
            O => \N__32112\,
            I => \N__32067\
        );

    \I__6103\ : InMux
    port map (
            O => \N__32111\,
            I => \N__32067\
        );

    \I__6102\ : InMux
    port map (
            O => \N__32110\,
            I => \N__32067\
        );

    \I__6101\ : InMux
    port map (
            O => \N__32109\,
            I => \N__32067\
        );

    \I__6100\ : LocalMux
    port map (
            O => \N__32100\,
            I => \N__32064\
        );

    \I__6099\ : Span4Mux_v
    port map (
            O => \N__32097\,
            I => \N__32059\
        );

    \I__6098\ : Span4Mux_v
    port map (
            O => \N__32086\,
            I => \N__32059\
        );

    \I__6097\ : Span12Mux_v
    port map (
            O => \N__32083\,
            I => \N__32056\
        );

    \I__6096\ : LocalMux
    port map (
            O => \N__32076\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__6095\ : LocalMux
    port map (
            O => \N__32067\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__6094\ : Odrv4
    port map (
            O => \N__32064\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__6093\ : Odrv4
    port map (
            O => \N__32059\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__6092\ : Odrv12
    port map (
            O => \N__32056\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__6091\ : InMux
    port map (
            O => \N__32045\,
            I => \N__32042\
        );

    \I__6090\ : LocalMux
    port map (
            O => \N__32042\,
            I => \N__32036\
        );

    \I__6089\ : InMux
    port map (
            O => \N__32041\,
            I => \N__32033\
        );

    \I__6088\ : InMux
    port map (
            O => \N__32040\,
            I => \N__32030\
        );

    \I__6087\ : InMux
    port map (
            O => \N__32039\,
            I => \N__32027\
        );

    \I__6086\ : Span4Mux_v
    port map (
            O => \N__32036\,
            I => \N__32022\
        );

    \I__6085\ : LocalMux
    port map (
            O => \N__32033\,
            I => \N__32022\
        );

    \I__6084\ : LocalMux
    port map (
            O => \N__32030\,
            I => \N__32017\
        );

    \I__6083\ : LocalMux
    port map (
            O => \N__32027\,
            I => \N__32017\
        );

    \I__6082\ : Span4Mux_v
    port map (
            O => \N__32022\,
            I => \N__32012\
        );

    \I__6081\ : Span4Mux_v
    port map (
            O => \N__32017\,
            I => \N__32012\
        );

    \I__6080\ : Odrv4
    port map (
            O => \N__32012\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__6079\ : InMux
    port map (
            O => \N__32009\,
            I => \N__32000\
        );

    \I__6078\ : InMux
    port map (
            O => \N__32008\,
            I => \N__31997\
        );

    \I__6077\ : InMux
    port map (
            O => \N__32007\,
            I => \N__31960\
        );

    \I__6076\ : InMux
    port map (
            O => \N__32006\,
            I => \N__31953\
        );

    \I__6075\ : InMux
    port map (
            O => \N__32005\,
            I => \N__31950\
        );

    \I__6074\ : InMux
    port map (
            O => \N__32004\,
            I => \N__31947\
        );

    \I__6073\ : InMux
    port map (
            O => \N__32003\,
            I => \N__31944\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__32000\,
            I => \N__31932\
        );

    \I__6071\ : LocalMux
    port map (
            O => \N__31997\,
            I => \N__31932\
        );

    \I__6070\ : InMux
    port map (
            O => \N__31996\,
            I => \N__31925\
        );

    \I__6069\ : InMux
    port map (
            O => \N__31995\,
            I => \N__31925\
        );

    \I__6068\ : InMux
    port map (
            O => \N__31994\,
            I => \N__31925\
        );

    \I__6067\ : InMux
    port map (
            O => \N__31993\,
            I => \N__31922\
        );

    \I__6066\ : InMux
    port map (
            O => \N__31992\,
            I => \N__31913\
        );

    \I__6065\ : InMux
    port map (
            O => \N__31991\,
            I => \N__31913\
        );

    \I__6064\ : InMux
    port map (
            O => \N__31990\,
            I => \N__31913\
        );

    \I__6063\ : InMux
    port map (
            O => \N__31989\,
            I => \N__31913\
        );

    \I__6062\ : CascadeMux
    port map (
            O => \N__31988\,
            I => \N__31895\
        );

    \I__6061\ : InMux
    port map (
            O => \N__31987\,
            I => \N__31885\
        );

    \I__6060\ : InMux
    port map (
            O => \N__31986\,
            I => \N__31885\
        );

    \I__6059\ : InMux
    port map (
            O => \N__31985\,
            I => \N__31885\
        );

    \I__6058\ : InMux
    port map (
            O => \N__31984\,
            I => \N__31885\
        );

    \I__6057\ : InMux
    port map (
            O => \N__31983\,
            I => \N__31882\
        );

    \I__6056\ : InMux
    port map (
            O => \N__31982\,
            I => \N__31865\
        );

    \I__6055\ : InMux
    port map (
            O => \N__31981\,
            I => \N__31865\
        );

    \I__6054\ : InMux
    port map (
            O => \N__31980\,
            I => \N__31865\
        );

    \I__6053\ : InMux
    port map (
            O => \N__31979\,
            I => \N__31865\
        );

    \I__6052\ : InMux
    port map (
            O => \N__31978\,
            I => \N__31865\
        );

    \I__6051\ : InMux
    port map (
            O => \N__31977\,
            I => \N__31865\
        );

    \I__6050\ : InMux
    port map (
            O => \N__31976\,
            I => \N__31865\
        );

    \I__6049\ : InMux
    port map (
            O => \N__31975\,
            I => \N__31865\
        );

    \I__6048\ : InMux
    port map (
            O => \N__31974\,
            I => \N__31854\
        );

    \I__6047\ : InMux
    port map (
            O => \N__31973\,
            I => \N__31854\
        );

    \I__6046\ : InMux
    port map (
            O => \N__31972\,
            I => \N__31854\
        );

    \I__6045\ : InMux
    port map (
            O => \N__31971\,
            I => \N__31854\
        );

    \I__6044\ : InMux
    port map (
            O => \N__31970\,
            I => \N__31854\
        );

    \I__6043\ : InMux
    port map (
            O => \N__31969\,
            I => \N__31849\
        );

    \I__6042\ : InMux
    port map (
            O => \N__31968\,
            I => \N__31849\
        );

    \I__6041\ : InMux
    port map (
            O => \N__31967\,
            I => \N__31838\
        );

    \I__6040\ : InMux
    port map (
            O => \N__31966\,
            I => \N__31838\
        );

    \I__6039\ : InMux
    port map (
            O => \N__31965\,
            I => \N__31838\
        );

    \I__6038\ : InMux
    port map (
            O => \N__31964\,
            I => \N__31838\
        );

    \I__6037\ : InMux
    port map (
            O => \N__31963\,
            I => \N__31838\
        );

    \I__6036\ : LocalMux
    port map (
            O => \N__31960\,
            I => \N__31835\
        );

    \I__6035\ : InMux
    port map (
            O => \N__31959\,
            I => \N__31830\
        );

    \I__6034\ : InMux
    port map (
            O => \N__31958\,
            I => \N__31823\
        );

    \I__6033\ : InMux
    port map (
            O => \N__31957\,
            I => \N__31823\
        );

    \I__6032\ : InMux
    port map (
            O => \N__31956\,
            I => \N__31823\
        );

    \I__6031\ : LocalMux
    port map (
            O => \N__31953\,
            I => \N__31816\
        );

    \I__6030\ : LocalMux
    port map (
            O => \N__31950\,
            I => \N__31816\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__31947\,
            I => \N__31816\
        );

    \I__6028\ : LocalMux
    port map (
            O => \N__31944\,
            I => \N__31809\
        );

    \I__6027\ : InMux
    port map (
            O => \N__31943\,
            I => \N__31806\
        );

    \I__6026\ : InMux
    port map (
            O => \N__31942\,
            I => \N__31801\
        );

    \I__6025\ : InMux
    port map (
            O => \N__31941\,
            I => \N__31801\
        );

    \I__6024\ : InMux
    port map (
            O => \N__31940\,
            I => \N__31796\
        );

    \I__6023\ : InMux
    port map (
            O => \N__31939\,
            I => \N__31796\
        );

    \I__6022\ : InMux
    port map (
            O => \N__31938\,
            I => \N__31793\
        );

    \I__6021\ : InMux
    port map (
            O => \N__31937\,
            I => \N__31790\
        );

    \I__6020\ : Span4Mux_h
    port map (
            O => \N__31932\,
            I => \N__31781\
        );

    \I__6019\ : LocalMux
    port map (
            O => \N__31925\,
            I => \N__31781\
        );

    \I__6018\ : LocalMux
    port map (
            O => \N__31922\,
            I => \N__31781\
        );

    \I__6017\ : LocalMux
    port map (
            O => \N__31913\,
            I => \N__31781\
        );

    \I__6016\ : InMux
    port map (
            O => \N__31912\,
            I => \N__31766\
        );

    \I__6015\ : InMux
    port map (
            O => \N__31911\,
            I => \N__31761\
        );

    \I__6014\ : InMux
    port map (
            O => \N__31910\,
            I => \N__31750\
        );

    \I__6013\ : InMux
    port map (
            O => \N__31909\,
            I => \N__31750\
        );

    \I__6012\ : InMux
    port map (
            O => \N__31908\,
            I => \N__31750\
        );

    \I__6011\ : InMux
    port map (
            O => \N__31907\,
            I => \N__31750\
        );

    \I__6010\ : InMux
    port map (
            O => \N__31906\,
            I => \N__31750\
        );

    \I__6009\ : InMux
    port map (
            O => \N__31905\,
            I => \N__31743\
        );

    \I__6008\ : InMux
    port map (
            O => \N__31904\,
            I => \N__31740\
        );

    \I__6007\ : InMux
    port map (
            O => \N__31903\,
            I => \N__31731\
        );

    \I__6006\ : InMux
    port map (
            O => \N__31902\,
            I => \N__31731\
        );

    \I__6005\ : InMux
    port map (
            O => \N__31901\,
            I => \N__31731\
        );

    \I__6004\ : InMux
    port map (
            O => \N__31900\,
            I => \N__31731\
        );

    \I__6003\ : InMux
    port map (
            O => \N__31899\,
            I => \N__31722\
        );

    \I__6002\ : InMux
    port map (
            O => \N__31898\,
            I => \N__31722\
        );

    \I__6001\ : InMux
    port map (
            O => \N__31895\,
            I => \N__31722\
        );

    \I__6000\ : InMux
    port map (
            O => \N__31894\,
            I => \N__31722\
        );

    \I__5999\ : LocalMux
    port map (
            O => \N__31885\,
            I => \N__31719\
        );

    \I__5998\ : LocalMux
    port map (
            O => \N__31882\,
            I => \N__31706\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__31865\,
            I => \N__31706\
        );

    \I__5996\ : LocalMux
    port map (
            O => \N__31854\,
            I => \N__31706\
        );

    \I__5995\ : LocalMux
    port map (
            O => \N__31849\,
            I => \N__31706\
        );

    \I__5994\ : LocalMux
    port map (
            O => \N__31838\,
            I => \N__31706\
        );

    \I__5993\ : Span4Mux_s3_v
    port map (
            O => \N__31835\,
            I => \N__31706\
        );

    \I__5992\ : InMux
    port map (
            O => \N__31834\,
            I => \N__31701\
        );

    \I__5991\ : InMux
    port map (
            O => \N__31833\,
            I => \N__31701\
        );

    \I__5990\ : LocalMux
    port map (
            O => \N__31830\,
            I => \N__31698\
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__31823\,
            I => \N__31693\
        );

    \I__5988\ : Span4Mux_v
    port map (
            O => \N__31816\,
            I => \N__31693\
        );

    \I__5987\ : InMux
    port map (
            O => \N__31815\,
            I => \N__31684\
        );

    \I__5986\ : InMux
    port map (
            O => \N__31814\,
            I => \N__31684\
        );

    \I__5985\ : InMux
    port map (
            O => \N__31813\,
            I => \N__31684\
        );

    \I__5984\ : InMux
    port map (
            O => \N__31812\,
            I => \N__31684\
        );

    \I__5983\ : Span4Mux_h
    port map (
            O => \N__31809\,
            I => \N__31679\
        );

    \I__5982\ : LocalMux
    port map (
            O => \N__31806\,
            I => \N__31679\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__31801\,
            I => \N__31674\
        );

    \I__5980\ : LocalMux
    port map (
            O => \N__31796\,
            I => \N__31674\
        );

    \I__5979\ : LocalMux
    port map (
            O => \N__31793\,
            I => \N__31671\
        );

    \I__5978\ : LocalMux
    port map (
            O => \N__31790\,
            I => \N__31668\
        );

    \I__5977\ : Span4Mux_v
    port map (
            O => \N__31781\,
            I => \N__31665\
        );

    \I__5976\ : InMux
    port map (
            O => \N__31780\,
            I => \N__31656\
        );

    \I__5975\ : InMux
    port map (
            O => \N__31779\,
            I => \N__31656\
        );

    \I__5974\ : InMux
    port map (
            O => \N__31778\,
            I => \N__31656\
        );

    \I__5973\ : InMux
    port map (
            O => \N__31777\,
            I => \N__31656\
        );

    \I__5972\ : InMux
    port map (
            O => \N__31776\,
            I => \N__31645\
        );

    \I__5971\ : InMux
    port map (
            O => \N__31775\,
            I => \N__31645\
        );

    \I__5970\ : InMux
    port map (
            O => \N__31774\,
            I => \N__31645\
        );

    \I__5969\ : InMux
    port map (
            O => \N__31773\,
            I => \N__31645\
        );

    \I__5968\ : InMux
    port map (
            O => \N__31772\,
            I => \N__31645\
        );

    \I__5967\ : InMux
    port map (
            O => \N__31771\,
            I => \N__31638\
        );

    \I__5966\ : InMux
    port map (
            O => \N__31770\,
            I => \N__31638\
        );

    \I__5965\ : InMux
    port map (
            O => \N__31769\,
            I => \N__31638\
        );

    \I__5964\ : LocalMux
    port map (
            O => \N__31766\,
            I => \N__31635\
        );

    \I__5963\ : InMux
    port map (
            O => \N__31765\,
            I => \N__31630\
        );

    \I__5962\ : InMux
    port map (
            O => \N__31764\,
            I => \N__31630\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__31761\,
            I => \N__31625\
        );

    \I__5960\ : LocalMux
    port map (
            O => \N__31750\,
            I => \N__31625\
        );

    \I__5959\ : InMux
    port map (
            O => \N__31749\,
            I => \N__31616\
        );

    \I__5958\ : InMux
    port map (
            O => \N__31748\,
            I => \N__31616\
        );

    \I__5957\ : InMux
    port map (
            O => \N__31747\,
            I => \N__31616\
        );

    \I__5956\ : InMux
    port map (
            O => \N__31746\,
            I => \N__31616\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__31743\,
            I => \N__31603\
        );

    \I__5954\ : LocalMux
    port map (
            O => \N__31740\,
            I => \N__31603\
        );

    \I__5953\ : LocalMux
    port map (
            O => \N__31731\,
            I => \N__31603\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__31722\,
            I => \N__31603\
        );

    \I__5951\ : Span4Mux_h
    port map (
            O => \N__31719\,
            I => \N__31603\
        );

    \I__5950\ : Span4Mux_v
    port map (
            O => \N__31706\,
            I => \N__31603\
        );

    \I__5949\ : LocalMux
    port map (
            O => \N__31701\,
            I => \N__31584\
        );

    \I__5948\ : Span4Mux_v
    port map (
            O => \N__31698\,
            I => \N__31584\
        );

    \I__5947\ : Span4Mux_v
    port map (
            O => \N__31693\,
            I => \N__31584\
        );

    \I__5946\ : LocalMux
    port map (
            O => \N__31684\,
            I => \N__31584\
        );

    \I__5945\ : Span4Mux_v
    port map (
            O => \N__31679\,
            I => \N__31584\
        );

    \I__5944\ : Span4Mux_v
    port map (
            O => \N__31674\,
            I => \N__31584\
        );

    \I__5943\ : Span4Mux_h
    port map (
            O => \N__31671\,
            I => \N__31584\
        );

    \I__5942\ : Span4Mux_v
    port map (
            O => \N__31668\,
            I => \N__31584\
        );

    \I__5941\ : Span4Mux_v
    port map (
            O => \N__31665\,
            I => \N__31584\
        );

    \I__5940\ : LocalMux
    port map (
            O => \N__31656\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__31645\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__5938\ : LocalMux
    port map (
            O => \N__31638\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__5937\ : Odrv4
    port map (
            O => \N__31635\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__5936\ : LocalMux
    port map (
            O => \N__31630\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__5935\ : Odrv12
    port map (
            O => \N__31625\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__5934\ : LocalMux
    port map (
            O => \N__31616\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__5933\ : Odrv4
    port map (
            O => \N__31603\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__5932\ : Odrv4
    port map (
            O => \N__31584\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__5931\ : InMux
    port map (
            O => \N__31565\,
            I => \N__31562\
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__31562\,
            I => \N__31557\
        );

    \I__5929\ : InMux
    port map (
            O => \N__31561\,
            I => \N__31554\
        );

    \I__5928\ : InMux
    port map (
            O => \N__31560\,
            I => \N__31551\
        );

    \I__5927\ : Span4Mux_h
    port map (
            O => \N__31557\,
            I => \N__31548\
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__31554\,
            I => \N__31545\
        );

    \I__5925\ : LocalMux
    port map (
            O => \N__31551\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20\
        );

    \I__5924\ : Odrv4
    port map (
            O => \N__31548\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20\
        );

    \I__5923\ : Odrv12
    port map (
            O => \N__31545\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20\
        );

    \I__5922\ : CascadeMux
    port map (
            O => \N__31538\,
            I => \current_shift_inst.un4_control_input1_1_cascade_\
        );

    \I__5921\ : CascadeMux
    port map (
            O => \N__31535\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7_cascade_\
        );

    \I__5920\ : InMux
    port map (
            O => \N__31532\,
            I => \N__31529\
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__31529\,
            I => \N__31526\
        );

    \I__5918\ : Span4Mux_h
    port map (
            O => \N__31526\,
            I => \N__31523\
        );

    \I__5917\ : Odrv4
    port map (
            O => \N__31523\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\
        );

    \I__5916\ : InMux
    port map (
            O => \N__31520\,
            I => \N__31517\
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__31517\,
            I => \N__31514\
        );

    \I__5914\ : Odrv12
    port map (
            O => \N__31514\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt20\
        );

    \I__5913\ : CascadeMux
    port map (
            O => \N__31511\,
            I => \N__31506\
        );

    \I__5912\ : InMux
    port map (
            O => \N__31510\,
            I => \N__31503\
        );

    \I__5911\ : InMux
    port map (
            O => \N__31509\,
            I => \N__31498\
        );

    \I__5910\ : InMux
    port map (
            O => \N__31506\,
            I => \N__31498\
        );

    \I__5909\ : LocalMux
    port map (
            O => \N__31503\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__31498\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__5907\ : CascadeMux
    port map (
            O => \N__31493\,
            I => \N__31488\
        );

    \I__5906\ : InMux
    port map (
            O => \N__31492\,
            I => \N__31485\
        );

    \I__5905\ : InMux
    port map (
            O => \N__31491\,
            I => \N__31480\
        );

    \I__5904\ : InMux
    port map (
            O => \N__31488\,
            I => \N__31480\
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__31485\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__5902\ : LocalMux
    port map (
            O => \N__31480\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__5901\ : CascadeMux
    port map (
            O => \N__31475\,
            I => \N__31472\
        );

    \I__5900\ : InMux
    port map (
            O => \N__31472\,
            I => \N__31469\
        );

    \I__5899\ : LocalMux
    port map (
            O => \N__31469\,
            I => \N__31466\
        );

    \I__5898\ : Odrv4
    port map (
            O => \N__31466\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20\
        );

    \I__5897\ : InMux
    port map (
            O => \N__31463\,
            I => \N__31457\
        );

    \I__5896\ : InMux
    port map (
            O => \N__31462\,
            I => \N__31457\
        );

    \I__5895\ : LocalMux
    port map (
            O => \N__31457\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_20\
        );

    \I__5894\ : InMux
    port map (
            O => \N__31454\,
            I => \N__31450\
        );

    \I__5893\ : InMux
    port map (
            O => \N__31453\,
            I => \N__31447\
        );

    \I__5892\ : LocalMux
    port map (
            O => \N__31450\,
            I => \N__31443\
        );

    \I__5891\ : LocalMux
    port map (
            O => \N__31447\,
            I => \N__31440\
        );

    \I__5890\ : InMux
    port map (
            O => \N__31446\,
            I => \N__31437\
        );

    \I__5889\ : Span12Mux_h
    port map (
            O => \N__31443\,
            I => \N__31434\
        );

    \I__5888\ : Span4Mux_h
    port map (
            O => \N__31440\,
            I => \N__31431\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__31437\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21\
        );

    \I__5886\ : Odrv12
    port map (
            O => \N__31434\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21\
        );

    \I__5885\ : Odrv4
    port map (
            O => \N__31431\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21\
        );

    \I__5884\ : InMux
    port map (
            O => \N__31424\,
            I => \N__31421\
        );

    \I__5883\ : LocalMux
    port map (
            O => \N__31421\,
            I => \N__31417\
        );

    \I__5882\ : InMux
    port map (
            O => \N__31420\,
            I => \N__31414\
        );

    \I__5881\ : Span4Mux_v
    port map (
            O => \N__31417\,
            I => \N__31410\
        );

    \I__5880\ : LocalMux
    port map (
            O => \N__31414\,
            I => \N__31406\
        );

    \I__5879\ : InMux
    port map (
            O => \N__31413\,
            I => \N__31403\
        );

    \I__5878\ : Span4Mux_v
    port map (
            O => \N__31410\,
            I => \N__31400\
        );

    \I__5877\ : InMux
    port map (
            O => \N__31409\,
            I => \N__31397\
        );

    \I__5876\ : Span4Mux_h
    port map (
            O => \N__31406\,
            I => \N__31392\
        );

    \I__5875\ : LocalMux
    port map (
            O => \N__31403\,
            I => \N__31392\
        );

    \I__5874\ : Span4Mux_h
    port map (
            O => \N__31400\,
            I => \N__31387\
        );

    \I__5873\ : LocalMux
    port map (
            O => \N__31397\,
            I => \N__31387\
        );

    \I__5872\ : Odrv4
    port map (
            O => \N__31392\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__5871\ : Odrv4
    port map (
            O => \N__31387\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__5870\ : InMux
    port map (
            O => \N__31382\,
            I => \N__31376\
        );

    \I__5869\ : InMux
    port map (
            O => \N__31381\,
            I => \N__31376\
        );

    \I__5868\ : LocalMux
    port map (
            O => \N__31376\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_21\
        );

    \I__5867\ : InMux
    port map (
            O => \N__31373\,
            I => \N__31368\
        );

    \I__5866\ : InMux
    port map (
            O => \N__31372\,
            I => \N__31363\
        );

    \I__5865\ : InMux
    port map (
            O => \N__31371\,
            I => \N__31363\
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__31368\,
            I => \N__31359\
        );

    \I__5863\ : LocalMux
    port map (
            O => \N__31363\,
            I => \N__31356\
        );

    \I__5862\ : InMux
    port map (
            O => \N__31362\,
            I => \N__31353\
        );

    \I__5861\ : Span4Mux_v
    port map (
            O => \N__31359\,
            I => \N__31350\
        );

    \I__5860\ : Span4Mux_h
    port map (
            O => \N__31356\,
            I => \N__31345\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__31353\,
            I => \N__31345\
        );

    \I__5858\ : Odrv4
    port map (
            O => \N__31350\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__5857\ : Odrv4
    port map (
            O => \N__31345\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__5856\ : InMux
    port map (
            O => \N__31340\,
            I => \N__31336\
        );

    \I__5855\ : InMux
    port map (
            O => \N__31339\,
            I => \N__31333\
        );

    \I__5854\ : LocalMux
    port map (
            O => \N__31336\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7\
        );

    \I__5853\ : LocalMux
    port map (
            O => \N__31333\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7\
        );

    \I__5852\ : InMux
    port map (
            O => \N__31328\,
            I => \N__31325\
        );

    \I__5851\ : LocalMux
    port map (
            O => \N__31325\,
            I => \N__31322\
        );

    \I__5850\ : Span4Mux_v
    port map (
            O => \N__31322\,
            I => \N__31319\
        );

    \I__5849\ : Odrv4
    port map (
            O => \N__31319\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\
        );

    \I__5848\ : CEMux
    port map (
            O => \N__31316\,
            I => \N__31286\
        );

    \I__5847\ : CEMux
    port map (
            O => \N__31315\,
            I => \N__31286\
        );

    \I__5846\ : CEMux
    port map (
            O => \N__31314\,
            I => \N__31286\
        );

    \I__5845\ : CEMux
    port map (
            O => \N__31313\,
            I => \N__31286\
        );

    \I__5844\ : CEMux
    port map (
            O => \N__31312\,
            I => \N__31286\
        );

    \I__5843\ : CEMux
    port map (
            O => \N__31311\,
            I => \N__31286\
        );

    \I__5842\ : CEMux
    port map (
            O => \N__31310\,
            I => \N__31286\
        );

    \I__5841\ : CEMux
    port map (
            O => \N__31309\,
            I => \N__31286\
        );

    \I__5840\ : CEMux
    port map (
            O => \N__31308\,
            I => \N__31286\
        );

    \I__5839\ : CEMux
    port map (
            O => \N__31307\,
            I => \N__31286\
        );

    \I__5838\ : GlobalMux
    port map (
            O => \N__31286\,
            I => \N__31283\
        );

    \I__5837\ : gio2CtrlBuf
    port map (
            O => \N__31283\,
            I => \phase_controller_inst2.stoper_hc.un1_start_g\
        );

    \I__5836\ : CascadeMux
    port map (
            O => \N__31280\,
            I => \N__31277\
        );

    \I__5835\ : InMux
    port map (
            O => \N__31277\,
            I => \N__31271\
        );

    \I__5834\ : InMux
    port map (
            O => \N__31276\,
            I => \N__31266\
        );

    \I__5833\ : InMux
    port map (
            O => \N__31275\,
            I => \N__31266\
        );

    \I__5832\ : InMux
    port map (
            O => \N__31274\,
            I => \N__31263\
        );

    \I__5831\ : LocalMux
    port map (
            O => \N__31271\,
            I => \N__31258\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__31266\,
            I => \N__31258\
        );

    \I__5829\ : LocalMux
    port map (
            O => \N__31263\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__5828\ : Odrv12
    port map (
            O => \N__31258\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__5827\ : InMux
    port map (
            O => \N__31253\,
            I => \N__31247\
        );

    \I__5826\ : InMux
    port map (
            O => \N__31252\,
            I => \N__31247\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__31247\,
            I => \N__31244\
        );

    \I__5824\ : Span4Mux_h
    port map (
            O => \N__31244\,
            I => \N__31241\
        );

    \I__5823\ : Odrv4
    port map (
            O => \N__31241\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__5822\ : InMux
    port map (
            O => \N__31238\,
            I => \N__31233\
        );

    \I__5821\ : InMux
    port map (
            O => \N__31237\,
            I => \N__31228\
        );

    \I__5820\ : InMux
    port map (
            O => \N__31236\,
            I => \N__31228\
        );

    \I__5819\ : LocalMux
    port map (
            O => \N__31233\,
            I => \N__31225\
        );

    \I__5818\ : LocalMux
    port map (
            O => \N__31228\,
            I => \N__31222\
        );

    \I__5817\ : Span4Mux_h
    port map (
            O => \N__31225\,
            I => \N__31219\
        );

    \I__5816\ : Span12Mux_h
    port map (
            O => \N__31222\,
            I => \N__31216\
        );

    \I__5815\ : IoSpan4Mux
    port map (
            O => \N__31219\,
            I => \N__31213\
        );

    \I__5814\ : Odrv12
    port map (
            O => \N__31216\,
            I => il_min_comp2_c
        );

    \I__5813\ : Odrv4
    port map (
            O => \N__31213\,
            I => il_min_comp2_c
        );

    \I__5812\ : InMux
    port map (
            O => \N__31208\,
            I => \N__31205\
        );

    \I__5811\ : LocalMux
    port map (
            O => \N__31205\,
            I => \N__31200\
        );

    \I__5810\ : InMux
    port map (
            O => \N__31204\,
            I => \N__31197\
        );

    \I__5809\ : InMux
    port map (
            O => \N__31203\,
            I => \N__31194\
        );

    \I__5808\ : Span4Mux_v
    port map (
            O => \N__31200\,
            I => \N__31187\
        );

    \I__5807\ : LocalMux
    port map (
            O => \N__31197\,
            I => \N__31187\
        );

    \I__5806\ : LocalMux
    port map (
            O => \N__31194\,
            I => \N__31187\
        );

    \I__5805\ : Span4Mux_h
    port map (
            O => \N__31187\,
            I => \N__31184\
        );

    \I__5804\ : Span4Mux_h
    port map (
            O => \N__31184\,
            I => \N__31181\
        );

    \I__5803\ : Odrv4
    port map (
            O => \N__31181\,
            I => il_max_comp2_c
        );

    \I__5802\ : InMux
    port map (
            O => \N__31178\,
            I => \N__31175\
        );

    \I__5801\ : LocalMux
    port map (
            O => \N__31175\,
            I => \N__31170\
        );

    \I__5800\ : CascadeMux
    port map (
            O => \N__31174\,
            I => \N__31166\
        );

    \I__5799\ : InMux
    port map (
            O => \N__31173\,
            I => \N__31163\
        );

    \I__5798\ : Span12Mux_s11_h
    port map (
            O => \N__31170\,
            I => \N__31160\
        );

    \I__5797\ : InMux
    port map (
            O => \N__31169\,
            I => \N__31157\
        );

    \I__5796\ : InMux
    port map (
            O => \N__31166\,
            I => \N__31154\
        );

    \I__5795\ : LocalMux
    port map (
            O => \N__31163\,
            I => \N__31151\
        );

    \I__5794\ : Span12Mux_v
    port map (
            O => \N__31160\,
            I => \N__31148\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__31157\,
            I => \N__31145\
        );

    \I__5792\ : LocalMux
    port map (
            O => \N__31154\,
            I => \N__31138\
        );

    \I__5791\ : Span12Mux_s5_v
    port map (
            O => \N__31151\,
            I => \N__31138\
        );

    \I__5790\ : Span12Mux_v
    port map (
            O => \N__31148\,
            I => \N__31138\
        );

    \I__5789\ : Odrv4
    port map (
            O => \N__31145\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__5788\ : Odrv12
    port map (
            O => \N__31138\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__5787\ : InMux
    port map (
            O => \N__31133\,
            I => \N__31129\
        );

    \I__5786\ : InMux
    port map (
            O => \N__31132\,
            I => \N__31125\
        );

    \I__5785\ : LocalMux
    port map (
            O => \N__31129\,
            I => \N__31122\
        );

    \I__5784\ : CascadeMux
    port map (
            O => \N__31128\,
            I => \N__31118\
        );

    \I__5783\ : LocalMux
    port map (
            O => \N__31125\,
            I => \N__31113\
        );

    \I__5782\ : Span4Mux_h
    port map (
            O => \N__31122\,
            I => \N__31113\
        );

    \I__5781\ : InMux
    port map (
            O => \N__31121\,
            I => \N__31110\
        );

    \I__5780\ : InMux
    port map (
            O => \N__31118\,
            I => \N__31107\
        );

    \I__5779\ : Span4Mux_v
    port map (
            O => \N__31113\,
            I => \N__31100\
        );

    \I__5778\ : LocalMux
    port map (
            O => \N__31110\,
            I => \N__31100\
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__31107\,
            I => \N__31100\
        );

    \I__5776\ : Odrv4
    port map (
            O => \N__31100\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__5775\ : InMux
    port map (
            O => \N__31097\,
            I => \N__31093\
        );

    \I__5774\ : InMux
    port map (
            O => \N__31096\,
            I => \N__31090\
        );

    \I__5773\ : LocalMux
    port map (
            O => \N__31093\,
            I => \N__31087\
        );

    \I__5772\ : LocalMux
    port map (
            O => \N__31090\,
            I => \N__31083\
        );

    \I__5771\ : Span4Mux_h
    port map (
            O => \N__31087\,
            I => \N__31080\
        );

    \I__5770\ : InMux
    port map (
            O => \N__31086\,
            I => \N__31077\
        );

    \I__5769\ : Span4Mux_v
    port map (
            O => \N__31083\,
            I => \N__31074\
        );

    \I__5768\ : Sp12to4
    port map (
            O => \N__31080\,
            I => \N__31071\
        );

    \I__5767\ : LocalMux
    port map (
            O => \N__31077\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28\
        );

    \I__5766\ : Odrv4
    port map (
            O => \N__31074\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28\
        );

    \I__5765\ : Odrv12
    port map (
            O => \N__31071\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28\
        );

    \I__5764\ : CascadeMux
    port map (
            O => \N__31064\,
            I => \N__31061\
        );

    \I__5763\ : InMux
    port map (
            O => \N__31061\,
            I => \N__31058\
        );

    \I__5762\ : LocalMux
    port map (
            O => \N__31058\,
            I => \N__31055\
        );

    \I__5761\ : Span4Mux_v
    port map (
            O => \N__31055\,
            I => \N__31052\
        );

    \I__5760\ : Span4Mux_h
    port map (
            O => \N__31052\,
            I => \N__31049\
        );

    \I__5759\ : Odrv4
    port map (
            O => \N__31049\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt28\
        );

    \I__5758\ : InMux
    port map (
            O => \N__31046\,
            I => \N__31043\
        );

    \I__5757\ : LocalMux
    port map (
            O => \N__31043\,
            I => \N__31040\
        );

    \I__5756\ : Span4Mux_h
    port map (
            O => \N__31040\,
            I => \N__31036\
        );

    \I__5755\ : InMux
    port map (
            O => \N__31039\,
            I => \N__31033\
        );

    \I__5754\ : Odrv4
    port map (
            O => \N__31036\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__31033\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29\
        );

    \I__5752\ : CascadeMux
    port map (
            O => \N__31028\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29_cascade_\
        );

    \I__5751\ : InMux
    port map (
            O => \N__31025\,
            I => \N__31018\
        );

    \I__5750\ : InMux
    port map (
            O => \N__31024\,
            I => \N__31018\
        );

    \I__5749\ : InMux
    port map (
            O => \N__31023\,
            I => \N__31015\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__31018\,
            I => \N__31012\
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__31015\,
            I => \N__31006\
        );

    \I__5746\ : Span4Mux_h
    port map (
            O => \N__31012\,
            I => \N__31006\
        );

    \I__5745\ : CascadeMux
    port map (
            O => \N__31011\,
            I => \N__31003\
        );

    \I__5744\ : Span4Mux_v
    port map (
            O => \N__31006\,
            I => \N__31000\
        );

    \I__5743\ : InMux
    port map (
            O => \N__31003\,
            I => \N__30997\
        );

    \I__5742\ : Odrv4
    port map (
            O => \N__31000\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__30997\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__5740\ : InMux
    port map (
            O => \N__30992\,
            I => \N__30986\
        );

    \I__5739\ : InMux
    port map (
            O => \N__30991\,
            I => \N__30986\
        );

    \I__5738\ : LocalMux
    port map (
            O => \N__30986\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_28\
        );

    \I__5737\ : InMux
    port map (
            O => \N__30983\,
            I => \N__30976\
        );

    \I__5736\ : InMux
    port map (
            O => \N__30982\,
            I => \N__30976\
        );

    \I__5735\ : InMux
    port map (
            O => \N__30981\,
            I => \N__30973\
        );

    \I__5734\ : LocalMux
    port map (
            O => \N__30976\,
            I => \N__30970\
        );

    \I__5733\ : LocalMux
    port map (
            O => \N__30973\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__5732\ : Odrv12
    port map (
            O => \N__30970\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__5731\ : CascadeMux
    port map (
            O => \N__30965\,
            I => \N__30961\
        );

    \I__5730\ : CascadeMux
    port map (
            O => \N__30964\,
            I => \N__30958\
        );

    \I__5729\ : InMux
    port map (
            O => \N__30961\,
            I => \N__30952\
        );

    \I__5728\ : InMux
    port map (
            O => \N__30958\,
            I => \N__30952\
        );

    \I__5727\ : InMux
    port map (
            O => \N__30957\,
            I => \N__30949\
        );

    \I__5726\ : LocalMux
    port map (
            O => \N__30952\,
            I => \N__30946\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__30949\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__5724\ : Odrv12
    port map (
            O => \N__30946\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__5723\ : InMux
    port map (
            O => \N__30941\,
            I => \N__30935\
        );

    \I__5722\ : InMux
    port map (
            O => \N__30940\,
            I => \N__30935\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__30935\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_29\
        );

    \I__5720\ : InMux
    port map (
            O => \N__30932\,
            I => \N__30929\
        );

    \I__5719\ : LocalMux
    port map (
            O => \N__30929\,
            I => \N__30926\
        );

    \I__5718\ : Span4Mux_h
    port map (
            O => \N__30926\,
            I => \N__30923\
        );

    \I__5717\ : Odrv4
    port map (
            O => \N__30923\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28\
        );

    \I__5716\ : InMux
    port map (
            O => \N__30920\,
            I => \N__30916\
        );

    \I__5715\ : InMux
    port map (
            O => \N__30919\,
            I => \N__30912\
        );

    \I__5714\ : LocalMux
    port map (
            O => \N__30916\,
            I => \N__30909\
        );

    \I__5713\ : InMux
    port map (
            O => \N__30915\,
            I => \N__30906\
        );

    \I__5712\ : LocalMux
    port map (
            O => \N__30912\,
            I => \N__30903\
        );

    \I__5711\ : Span4Mux_v
    port map (
            O => \N__30909\,
            I => \N__30900\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__30906\,
            I => \N__30895\
        );

    \I__5709\ : Span4Mux_h
    port map (
            O => \N__30903\,
            I => \N__30895\
        );

    \I__5708\ : Span4Mux_h
    port map (
            O => \N__30900\,
            I => \N__30890\
        );

    \I__5707\ : Span4Mux_v
    port map (
            O => \N__30895\,
            I => \N__30890\
        );

    \I__5706\ : Odrv4
    port map (
            O => \N__30890\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__5705\ : InMux
    port map (
            O => \N__30887\,
            I => \N__30884\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__30884\,
            I => \N__30881\
        );

    \I__5703\ : Glb2LocalMux
    port map (
            O => \N__30881\,
            I => \N__30878\
        );

    \I__5702\ : GlobalMux
    port map (
            O => \N__30878\,
            I => clk_12mhz
        );

    \I__5701\ : IoInMux
    port map (
            O => \N__30875\,
            I => \N__30872\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__30872\,
            I => \GB_BUFFER_clk_12mhz_THRU_CO\
        );

    \I__5699\ : InMux
    port map (
            O => \N__30869\,
            I => \N__30866\
        );

    \I__5698\ : LocalMux
    port map (
            O => \N__30866\,
            I => \phase_controller_inst2.start_timer_tr_RNO_0_0\
        );

    \I__5697\ : InMux
    port map (
            O => \N__30863\,
            I => \N__30858\
        );

    \I__5696\ : InMux
    port map (
            O => \N__30862\,
            I => \N__30853\
        );

    \I__5695\ : InMux
    port map (
            O => \N__30861\,
            I => \N__30853\
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__30858\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__5693\ : LocalMux
    port map (
            O => \N__30853\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__5692\ : InMux
    port map (
            O => \N__30848\,
            I => \N__30845\
        );

    \I__5691\ : LocalMux
    port map (
            O => \N__30845\,
            I => \phase_controller_inst2.start_timer_hc_0_sqmuxa\
        );

    \I__5690\ : InMux
    port map (
            O => \N__30842\,
            I => \N__30839\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__30839\,
            I => \N__30835\
        );

    \I__5688\ : InMux
    port map (
            O => \N__30838\,
            I => \N__30832\
        );

    \I__5687\ : Odrv4
    port map (
            O => \N__30835\,
            I => \phase_controller_inst2.state_RNIG7JFZ0Z_2\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__30832\,
            I => \phase_controller_inst2.state_RNIG7JFZ0Z_2\
        );

    \I__5685\ : InMux
    port map (
            O => \N__30827\,
            I => \N__30821\
        );

    \I__5684\ : InMux
    port map (
            O => \N__30826\,
            I => \N__30821\
        );

    \I__5683\ : LocalMux
    port map (
            O => \N__30821\,
            I => \N__30818\
        );

    \I__5682\ : Span4Mux_s3_v
    port map (
            O => \N__30818\,
            I => \N__30815\
        );

    \I__5681\ : Span4Mux_h
    port map (
            O => \N__30815\,
            I => \N__30812\
        );

    \I__5680\ : Sp12to4
    port map (
            O => \N__30812\,
            I => \N__30807\
        );

    \I__5679\ : InMux
    port map (
            O => \N__30811\,
            I => \N__30804\
        );

    \I__5678\ : InMux
    port map (
            O => \N__30810\,
            I => \N__30801\
        );

    \I__5677\ : Span12Mux_v
    port map (
            O => \N__30807\,
            I => \N__30798\
        );

    \I__5676\ : LocalMux
    port map (
            O => \N__30804\,
            I => \N__30793\
        );

    \I__5675\ : LocalMux
    port map (
            O => \N__30801\,
            I => \N__30793\
        );

    \I__5674\ : Span12Mux_v
    port map (
            O => \N__30798\,
            I => \N__30790\
        );

    \I__5673\ : Span12Mux_h
    port map (
            O => \N__30793\,
            I => \N__30787\
        );

    \I__5672\ : Span12Mux_h
    port map (
            O => \N__30790\,
            I => \N__30782\
        );

    \I__5671\ : Span12Mux_v
    port map (
            O => \N__30787\,
            I => \N__30782\
        );

    \I__5670\ : Odrv12
    port map (
            O => \N__30782\,
            I => start_stop_c
        );

    \I__5669\ : InMux
    port map (
            O => \N__30779\,
            I => \N__30776\
        );

    \I__5668\ : LocalMux
    port map (
            O => \N__30776\,
            I => \N__30772\
        );

    \I__5667\ : InMux
    port map (
            O => \N__30775\,
            I => \N__30769\
        );

    \I__5666\ : Span4Mux_h
    port map (
            O => \N__30772\,
            I => \N__30762\
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__30769\,
            I => \N__30762\
        );

    \I__5664\ : InMux
    port map (
            O => \N__30768\,
            I => \N__30759\
        );

    \I__5663\ : InMux
    port map (
            O => \N__30767\,
            I => \N__30756\
        );

    \I__5662\ : Odrv4
    port map (
            O => \N__30762\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__30759\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__5660\ : LocalMux
    port map (
            O => \N__30756\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__5659\ : InMux
    port map (
            O => \N__30749\,
            I => \N__30746\
        );

    \I__5658\ : LocalMux
    port map (
            O => \N__30746\,
            I => \N__30741\
        );

    \I__5657\ : InMux
    port map (
            O => \N__30745\,
            I => \N__30738\
        );

    \I__5656\ : InMux
    port map (
            O => \N__30744\,
            I => \N__30735\
        );

    \I__5655\ : Span4Mux_h
    port map (
            O => \N__30741\,
            I => \N__30730\
        );

    \I__5654\ : LocalMux
    port map (
            O => \N__30738\,
            I => \N__30730\
        );

    \I__5653\ : LocalMux
    port map (
            O => \N__30735\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26\
        );

    \I__5652\ : Odrv4
    port map (
            O => \N__30730\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26\
        );

    \I__5651\ : CascadeMux
    port map (
            O => \N__30725\,
            I => \N__30721\
        );

    \I__5650\ : InMux
    port map (
            O => \N__30724\,
            I => \N__30716\
        );

    \I__5649\ : InMux
    port map (
            O => \N__30721\,
            I => \N__30713\
        );

    \I__5648\ : InMux
    port map (
            O => \N__30720\,
            I => \N__30710\
        );

    \I__5647\ : InMux
    port map (
            O => \N__30719\,
            I => \N__30707\
        );

    \I__5646\ : LocalMux
    port map (
            O => \N__30716\,
            I => \N__30702\
        );

    \I__5645\ : LocalMux
    port map (
            O => \N__30713\,
            I => \N__30702\
        );

    \I__5644\ : LocalMux
    port map (
            O => \N__30710\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__30707\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__5642\ : Odrv4
    port map (
            O => \N__30702\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__5641\ : InMux
    port map (
            O => \N__30695\,
            I => \N__30690\
        );

    \I__5640\ : InMux
    port map (
            O => \N__30694\,
            I => \N__30685\
        );

    \I__5639\ : InMux
    port map (
            O => \N__30693\,
            I => \N__30685\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__30690\,
            I => \N__30680\
        );

    \I__5637\ : LocalMux
    port map (
            O => \N__30685\,
            I => \N__30680\
        );

    \I__5636\ : Odrv4
    port map (
            O => \N__30680\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__5635\ : ClkMux
    port map (
            O => \N__30677\,
            I => \N__30671\
        );

    \I__5634\ : ClkMux
    port map (
            O => \N__30676\,
            I => \N__30671\
        );

    \I__5633\ : GlobalMux
    port map (
            O => \N__30671\,
            I => \N__30668\
        );

    \I__5632\ : gio2CtrlBuf
    port map (
            O => \N__30668\,
            I => delay_tr_input_c_g
        );

    \I__5631\ : InMux
    port map (
            O => \N__30665\,
            I => \N__30660\
        );

    \I__5630\ : InMux
    port map (
            O => \N__30664\,
            I => \N__30657\
        );

    \I__5629\ : InMux
    port map (
            O => \N__30663\,
            I => \N__30654\
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__30660\,
            I => \N__30651\
        );

    \I__5627\ : LocalMux
    port map (
            O => \N__30657\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__5626\ : LocalMux
    port map (
            O => \N__30654\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__5625\ : Odrv4
    port map (
            O => \N__30651\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__5624\ : InMux
    port map (
            O => \N__30644\,
            I => \N__30639\
        );

    \I__5623\ : InMux
    port map (
            O => \N__30643\,
            I => \N__30636\
        );

    \I__5622\ : InMux
    port map (
            O => \N__30642\,
            I => \N__30633\
        );

    \I__5621\ : LocalMux
    port map (
            O => \N__30639\,
            I => \N__30630\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__30636\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__5619\ : LocalMux
    port map (
            O => \N__30633\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__5618\ : Odrv4
    port map (
            O => \N__30630\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__5617\ : InMux
    port map (
            O => \N__30623\,
            I => \N__30619\
        );

    \I__5616\ : InMux
    port map (
            O => \N__30622\,
            I => \N__30615\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__30619\,
            I => \N__30612\
        );

    \I__5614\ : InMux
    port map (
            O => \N__30618\,
            I => \N__30609\
        );

    \I__5613\ : LocalMux
    port map (
            O => \N__30615\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__5612\ : Odrv4
    port map (
            O => \N__30612\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__30609\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__5610\ : InMux
    port map (
            O => \N__30602\,
            I => \N__30599\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__30599\,
            I => \pwm_generator_inst.un1_counterlto9_2\
        );

    \I__5608\ : CascadeMux
    port map (
            O => \N__30596\,
            I => \N__30592\
        );

    \I__5607\ : InMux
    port map (
            O => \N__30595\,
            I => \N__30588\
        );

    \I__5606\ : InMux
    port map (
            O => \N__30592\,
            I => \N__30585\
        );

    \I__5605\ : InMux
    port map (
            O => \N__30591\,
            I => \N__30582\
        );

    \I__5604\ : LocalMux
    port map (
            O => \N__30588\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__5603\ : LocalMux
    port map (
            O => \N__30585\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__30582\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__5601\ : InMux
    port map (
            O => \N__30575\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\
        );

    \I__5600\ : InMux
    port map (
            O => \N__30572\,
            I => \N__30567\
        );

    \I__5599\ : InMux
    port map (
            O => \N__30571\,
            I => \N__30564\
        );

    \I__5598\ : InMux
    port map (
            O => \N__30570\,
            I => \N__30561\
        );

    \I__5597\ : LocalMux
    port map (
            O => \N__30567\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__5596\ : LocalMux
    port map (
            O => \N__30564\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__5595\ : LocalMux
    port map (
            O => \N__30561\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__5594\ : InMux
    port map (
            O => \N__30554\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\
        );

    \I__5593\ : InMux
    port map (
            O => \N__30551\,
            I => \N__30541\
        );

    \I__5592\ : InMux
    port map (
            O => \N__30550\,
            I => \N__30541\
        );

    \I__5591\ : InMux
    port map (
            O => \N__30549\,
            I => \N__30541\
        );

    \I__5590\ : InMux
    port map (
            O => \N__30548\,
            I => \N__30538\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__30541\,
            I => \N__30535\
        );

    \I__5588\ : LocalMux
    port map (
            O => \N__30538\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__5587\ : Odrv12
    port map (
            O => \N__30535\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__5586\ : InMux
    port map (
            O => \N__30530\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\
        );

    \I__5585\ : InMux
    port map (
            O => \N__30527\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\
        );

    \I__5584\ : InMux
    port map (
            O => \N__30524\,
            I => \N__30521\
        );

    \I__5583\ : LocalMux
    port map (
            O => \N__30521\,
            I => \N__30515\
        );

    \I__5582\ : InMux
    port map (
            O => \N__30520\,
            I => \N__30510\
        );

    \I__5581\ : InMux
    port map (
            O => \N__30519\,
            I => \N__30510\
        );

    \I__5580\ : InMux
    port map (
            O => \N__30518\,
            I => \N__30507\
        );

    \I__5579\ : Sp12to4
    port map (
            O => \N__30515\,
            I => \N__30502\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__30510\,
            I => \N__30502\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__30507\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__5576\ : Odrv12
    port map (
            O => \N__30502\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__5575\ : InMux
    port map (
            O => \N__30497\,
            I => \N__30494\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__30494\,
            I => \N__30490\
        );

    \I__5573\ : InMux
    port map (
            O => \N__30493\,
            I => \N__30487\
        );

    \I__5572\ : Odrv4
    port map (
            O => \N__30490\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\
        );

    \I__5571\ : LocalMux
    port map (
            O => \N__30487\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\
        );

    \I__5570\ : InMux
    port map (
            O => \N__30482\,
            I => \N__30479\
        );

    \I__5569\ : LocalMux
    port map (
            O => \N__30479\,
            I => \N__30476\
        );

    \I__5568\ : Span4Mux_v
    port map (
            O => \N__30476\,
            I => \N__30473\
        );

    \I__5567\ : Odrv4
    port map (
            O => \N__30473\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\
        );

    \I__5566\ : InMux
    port map (
            O => \N__30470\,
            I => \N__30467\
        );

    \I__5565\ : LocalMux
    port map (
            O => \N__30467\,
            I => \N__30461\
        );

    \I__5564\ : InMux
    port map (
            O => \N__30466\,
            I => \N__30458\
        );

    \I__5563\ : InMux
    port map (
            O => \N__30465\,
            I => \N__30455\
        );

    \I__5562\ : InMux
    port map (
            O => \N__30464\,
            I => \N__30452\
        );

    \I__5561\ : Odrv4
    port map (
            O => \N__30461\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__5560\ : LocalMux
    port map (
            O => \N__30458\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__5559\ : LocalMux
    port map (
            O => \N__30455\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__5558\ : LocalMux
    port map (
            O => \N__30452\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__5557\ : InMux
    port map (
            O => \N__30443\,
            I => \N__30440\
        );

    \I__5556\ : LocalMux
    port map (
            O => \N__30440\,
            I => \N__30436\
        );

    \I__5555\ : InMux
    port map (
            O => \N__30439\,
            I => \N__30432\
        );

    \I__5554\ : Span4Mux_h
    port map (
            O => \N__30436\,
            I => \N__30429\
        );

    \I__5553\ : InMux
    port map (
            O => \N__30435\,
            I => \N__30426\
        );

    \I__5552\ : LocalMux
    port map (
            O => \N__30432\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13\
        );

    \I__5551\ : Odrv4
    port map (
            O => \N__30429\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13\
        );

    \I__5550\ : LocalMux
    port map (
            O => \N__30426\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13\
        );

    \I__5549\ : CascadeMux
    port map (
            O => \N__30419\,
            I => \N__30416\
        );

    \I__5548\ : InMux
    port map (
            O => \N__30416\,
            I => \N__30410\
        );

    \I__5547\ : InMux
    port map (
            O => \N__30415\,
            I => \N__30410\
        );

    \I__5546\ : LocalMux
    port map (
            O => \N__30410\,
            I => \N__30406\
        );

    \I__5545\ : InMux
    port map (
            O => \N__30409\,
            I => \N__30403\
        );

    \I__5544\ : Span4Mux_h
    port map (
            O => \N__30406\,
            I => \N__30400\
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__30403\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__5542\ : Odrv4
    port map (
            O => \N__30400\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__5541\ : InMux
    port map (
            O => \N__30395\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\
        );

    \I__5540\ : InMux
    port map (
            O => \N__30392\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\
        );

    \I__5539\ : InMux
    port map (
            O => \N__30389\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__5538\ : CascadeMux
    port map (
            O => \N__30386\,
            I => \N__30383\
        );

    \I__5537\ : InMux
    port map (
            O => \N__30383\,
            I => \N__30377\
        );

    \I__5536\ : InMux
    port map (
            O => \N__30382\,
            I => \N__30377\
        );

    \I__5535\ : LocalMux
    port map (
            O => \N__30377\,
            I => \N__30373\
        );

    \I__5534\ : InMux
    port map (
            O => \N__30376\,
            I => \N__30370\
        );

    \I__5533\ : Span4Mux_h
    port map (
            O => \N__30373\,
            I => \N__30367\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__30370\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__5531\ : Odrv4
    port map (
            O => \N__30367\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__5530\ : InMux
    port map (
            O => \N__30362\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\
        );

    \I__5529\ : InMux
    port map (
            O => \N__30359\,
            I => \N__30353\
        );

    \I__5528\ : InMux
    port map (
            O => \N__30358\,
            I => \N__30353\
        );

    \I__5527\ : LocalMux
    port map (
            O => \N__30353\,
            I => \N__30349\
        );

    \I__5526\ : InMux
    port map (
            O => \N__30352\,
            I => \N__30346\
        );

    \I__5525\ : Span4Mux_h
    port map (
            O => \N__30349\,
            I => \N__30343\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__30346\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__5523\ : Odrv4
    port map (
            O => \N__30343\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__5522\ : InMux
    port map (
            O => \N__30338\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\
        );

    \I__5521\ : InMux
    port map (
            O => \N__30335\,
            I => \N__30330\
        );

    \I__5520\ : InMux
    port map (
            O => \N__30334\,
            I => \N__30325\
        );

    \I__5519\ : InMux
    port map (
            O => \N__30333\,
            I => \N__30325\
        );

    \I__5518\ : LocalMux
    port map (
            O => \N__30330\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__5517\ : LocalMux
    port map (
            O => \N__30325\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__5516\ : InMux
    port map (
            O => \N__30320\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\
        );

    \I__5515\ : CascadeMux
    port map (
            O => \N__30317\,
            I => \N__30312\
        );

    \I__5514\ : InMux
    port map (
            O => \N__30316\,
            I => \N__30309\
        );

    \I__5513\ : InMux
    port map (
            O => \N__30315\,
            I => \N__30304\
        );

    \I__5512\ : InMux
    port map (
            O => \N__30312\,
            I => \N__30304\
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__30309\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__30304\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__5509\ : InMux
    port map (
            O => \N__30299\,
            I => \bfn_11_11_0_\
        );

    \I__5508\ : InMux
    port map (
            O => \N__30296\,
            I => \N__30291\
        );

    \I__5507\ : InMux
    port map (
            O => \N__30295\,
            I => \N__30288\
        );

    \I__5506\ : InMux
    port map (
            O => \N__30294\,
            I => \N__30285\
        );

    \I__5505\ : LocalMux
    port map (
            O => \N__30291\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__30288\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__30285\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__5502\ : InMux
    port map (
            O => \N__30278\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\
        );

    \I__5501\ : CascadeMux
    port map (
            O => \N__30275\,
            I => \N__30271\
        );

    \I__5500\ : CascadeMux
    port map (
            O => \N__30274\,
            I => \N__30267\
        );

    \I__5499\ : InMux
    port map (
            O => \N__30271\,
            I => \N__30264\
        );

    \I__5498\ : InMux
    port map (
            O => \N__30270\,
            I => \N__30261\
        );

    \I__5497\ : InMux
    port map (
            O => \N__30267\,
            I => \N__30258\
        );

    \I__5496\ : LocalMux
    port map (
            O => \N__30264\,
            I => \N__30255\
        );

    \I__5495\ : LocalMux
    port map (
            O => \N__30261\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__5494\ : LocalMux
    port map (
            O => \N__30258\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__5493\ : Odrv4
    port map (
            O => \N__30255\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__5492\ : InMux
    port map (
            O => \N__30248\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\
        );

    \I__5491\ : InMux
    port map (
            O => \N__30245\,
            I => \N__30241\
        );

    \I__5490\ : InMux
    port map (
            O => \N__30244\,
            I => \N__30238\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__30241\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__5488\ : LocalMux
    port map (
            O => \N__30238\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__5487\ : InMux
    port map (
            O => \N__30233\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\
        );

    \I__5486\ : InMux
    port map (
            O => \N__30230\,
            I => \N__30226\
        );

    \I__5485\ : InMux
    port map (
            O => \N__30229\,
            I => \N__30223\
        );

    \I__5484\ : LocalMux
    port map (
            O => \N__30226\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__30223\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__5482\ : InMux
    port map (
            O => \N__30218\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\
        );

    \I__5481\ : InMux
    port map (
            O => \N__30215\,
            I => \N__30211\
        );

    \I__5480\ : InMux
    port map (
            O => \N__30214\,
            I => \N__30208\
        );

    \I__5479\ : LocalMux
    port map (
            O => \N__30211\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__30208\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__5477\ : InMux
    port map (
            O => \N__30203\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\
        );

    \I__5476\ : InMux
    port map (
            O => \N__30200\,
            I => \N__30196\
        );

    \I__5475\ : InMux
    port map (
            O => \N__30199\,
            I => \N__30193\
        );

    \I__5474\ : LocalMux
    port map (
            O => \N__30196\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__30193\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__5472\ : InMux
    port map (
            O => \N__30188\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\
        );

    \I__5471\ : InMux
    port map (
            O => \N__30185\,
            I => \N__30181\
        );

    \I__5470\ : InMux
    port map (
            O => \N__30184\,
            I => \N__30178\
        );

    \I__5469\ : LocalMux
    port map (
            O => \N__30181\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__30178\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__5467\ : InMux
    port map (
            O => \N__30173\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\
        );

    \I__5466\ : CascadeMux
    port map (
            O => \N__30170\,
            I => \N__30166\
        );

    \I__5465\ : InMux
    port map (
            O => \N__30169\,
            I => \N__30161\
        );

    \I__5464\ : InMux
    port map (
            O => \N__30166\,
            I => \N__30161\
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__30161\,
            I => \N__30157\
        );

    \I__5462\ : InMux
    port map (
            O => \N__30160\,
            I => \N__30154\
        );

    \I__5461\ : Span4Mux_h
    port map (
            O => \N__30157\,
            I => \N__30151\
        );

    \I__5460\ : LocalMux
    port map (
            O => \N__30154\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__5459\ : Odrv4
    port map (
            O => \N__30151\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__5458\ : InMux
    port map (
            O => \N__30146\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\
        );

    \I__5457\ : CascadeMux
    port map (
            O => \N__30143\,
            I => \N__30140\
        );

    \I__5456\ : InMux
    port map (
            O => \N__30140\,
            I => \N__30135\
        );

    \I__5455\ : InMux
    port map (
            O => \N__30139\,
            I => \N__30132\
        );

    \I__5454\ : InMux
    port map (
            O => \N__30138\,
            I => \N__30129\
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__30135\,
            I => \N__30124\
        );

    \I__5452\ : LocalMux
    port map (
            O => \N__30132\,
            I => \N__30124\
        );

    \I__5451\ : LocalMux
    port map (
            O => \N__30129\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__5450\ : Odrv12
    port map (
            O => \N__30124\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__5449\ : InMux
    port map (
            O => \N__30119\,
            I => \bfn_11_10_0_\
        );

    \I__5448\ : InMux
    port map (
            O => \N__30116\,
            I => \N__30110\
        );

    \I__5447\ : InMux
    port map (
            O => \N__30115\,
            I => \N__30110\
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__30110\,
            I => \N__30106\
        );

    \I__5445\ : InMux
    port map (
            O => \N__30109\,
            I => \N__30103\
        );

    \I__5444\ : Span4Mux_h
    port map (
            O => \N__30106\,
            I => \N__30100\
        );

    \I__5443\ : LocalMux
    port map (
            O => \N__30103\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__5442\ : Odrv4
    port map (
            O => \N__30100\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__5441\ : InMux
    port map (
            O => \N__30095\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\
        );

    \I__5440\ : CascadeMux
    port map (
            O => \N__30092\,
            I => \N__30089\
        );

    \I__5439\ : InMux
    port map (
            O => \N__30089\,
            I => \N__30086\
        );

    \I__5438\ : LocalMux
    port map (
            O => \N__30086\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3Z0Z_28\
        );

    \I__5437\ : InMux
    port map (
            O => \N__30083\,
            I => \N__30079\
        );

    \I__5436\ : InMux
    port map (
            O => \N__30082\,
            I => \N__30076\
        );

    \I__5435\ : LocalMux
    port map (
            O => \N__30079\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__30076\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__5433\ : InMux
    port map (
            O => \N__30071\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\
        );

    \I__5432\ : InMux
    port map (
            O => \N__30068\,
            I => \N__30064\
        );

    \I__5431\ : InMux
    port map (
            O => \N__30067\,
            I => \N__30061\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__30064\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__5429\ : LocalMux
    port map (
            O => \N__30061\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__5428\ : InMux
    port map (
            O => \N__30056\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\
        );

    \I__5427\ : InMux
    port map (
            O => \N__30053\,
            I => \N__30049\
        );

    \I__5426\ : InMux
    port map (
            O => \N__30052\,
            I => \N__30046\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__30049\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__30046\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__5423\ : InMux
    port map (
            O => \N__30041\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\
        );

    \I__5422\ : InMux
    port map (
            O => \N__30038\,
            I => \N__30034\
        );

    \I__5421\ : InMux
    port map (
            O => \N__30037\,
            I => \N__30031\
        );

    \I__5420\ : LocalMux
    port map (
            O => \N__30034\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__5419\ : LocalMux
    port map (
            O => \N__30031\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__5418\ : InMux
    port map (
            O => \N__30026\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\
        );

    \I__5417\ : InMux
    port map (
            O => \N__30023\,
            I => \N__30019\
        );

    \I__5416\ : InMux
    port map (
            O => \N__30022\,
            I => \N__30016\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__30019\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__5414\ : LocalMux
    port map (
            O => \N__30016\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__5413\ : InMux
    port map (
            O => \N__30011\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\
        );

    \I__5412\ : InMux
    port map (
            O => \N__30008\,
            I => \N__30004\
        );

    \I__5411\ : InMux
    port map (
            O => \N__30007\,
            I => \N__30001\
        );

    \I__5410\ : LocalMux
    port map (
            O => \N__30004\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__5409\ : LocalMux
    port map (
            O => \N__30001\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__5408\ : InMux
    port map (
            O => \N__29996\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\
        );

    \I__5407\ : InMux
    port map (
            O => \N__29993\,
            I => \N__29989\
        );

    \I__5406\ : InMux
    port map (
            O => \N__29992\,
            I => \N__29986\
        );

    \I__5405\ : LocalMux
    port map (
            O => \N__29989\,
            I => \N__29983\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__29986\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__5403\ : Odrv4
    port map (
            O => \N__29983\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__5402\ : InMux
    port map (
            O => \N__29978\,
            I => \bfn_11_9_0_\
        );

    \I__5401\ : InMux
    port map (
            O => \N__29975\,
            I => \N__29971\
        );

    \I__5400\ : InMux
    port map (
            O => \N__29974\,
            I => \N__29968\
        );

    \I__5399\ : LocalMux
    port map (
            O => \N__29971\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__5398\ : LocalMux
    port map (
            O => \N__29968\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__5397\ : InMux
    port map (
            O => \N__29963\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\
        );

    \I__5396\ : CascadeMux
    port map (
            O => \N__29960\,
            I => \phase_controller_inst2.stoper_hc.un4_running_df30_cascade_\
        );

    \I__5395\ : InMux
    port map (
            O => \N__29957\,
            I => \N__29954\
        );

    \I__5394\ : LocalMux
    port map (
            O => \N__29954\,
            I => \N__29951\
        );

    \I__5393\ : Odrv4
    port map (
            O => \N__29951\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO\
        );

    \I__5392\ : CascadeMux
    port map (
            O => \N__29948\,
            I => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\
        );

    \I__5391\ : CascadeMux
    port map (
            O => \N__29945\,
            I => \N__29942\
        );

    \I__5390\ : InMux
    port map (
            O => \N__29942\,
            I => \N__29939\
        );

    \I__5389\ : LocalMux
    port map (
            O => \N__29939\,
            I => \N__29936\
        );

    \I__5388\ : Span4Mux_v
    port map (
            O => \N__29936\,
            I => \N__29932\
        );

    \I__5387\ : InMux
    port map (
            O => \N__29935\,
            I => \N__29929\
        );

    \I__5386\ : Odrv4
    port map (
            O => \N__29932\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt30\
        );

    \I__5385\ : LocalMux
    port map (
            O => \N__29929\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt30\
        );

    \I__5384\ : CascadeMux
    port map (
            O => \N__29924\,
            I => \N__29921\
        );

    \I__5383\ : InMux
    port map (
            O => \N__29921\,
            I => \N__29916\
        );

    \I__5382\ : InMux
    port map (
            O => \N__29920\,
            I => \N__29911\
        );

    \I__5381\ : InMux
    port map (
            O => \N__29919\,
            I => \N__29911\
        );

    \I__5380\ : LocalMux
    port map (
            O => \N__29916\,
            I => \N__29908\
        );

    \I__5379\ : LocalMux
    port map (
            O => \N__29911\,
            I => \N__29905\
        );

    \I__5378\ : Span4Mux_v
    port map (
            O => \N__29908\,
            I => \N__29902\
        );

    \I__5377\ : Span4Mux_v
    port map (
            O => \N__29905\,
            I => \N__29899\
        );

    \I__5376\ : Odrv4
    port map (
            O => \N__29902\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_30\
        );

    \I__5375\ : Odrv4
    port map (
            O => \N__29899\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_30\
        );

    \I__5374\ : CascadeMux
    port map (
            O => \N__29894\,
            I => \N__29890\
        );

    \I__5373\ : CascadeMux
    port map (
            O => \N__29893\,
            I => \N__29886\
        );

    \I__5372\ : InMux
    port map (
            O => \N__29890\,
            I => \N__29879\
        );

    \I__5371\ : InMux
    port map (
            O => \N__29889\,
            I => \N__29879\
        );

    \I__5370\ : InMux
    port map (
            O => \N__29886\,
            I => \N__29879\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__29879\,
            I => \N__29876\
        );

    \I__5368\ : Span4Mux_v
    port map (
            O => \N__29876\,
            I => \N__29873\
        );

    \I__5367\ : Odrv4
    port map (
            O => \N__29873\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\
        );

    \I__5366\ : InMux
    port map (
            O => \N__29870\,
            I => \N__29867\
        );

    \I__5365\ : LocalMux
    port map (
            O => \N__29867\,
            I => \N__29864\
        );

    \I__5364\ : Odrv4
    port map (
            O => \N__29864\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\
        );

    \I__5363\ : InMux
    port map (
            O => \N__29861\,
            I => \N__29855\
        );

    \I__5362\ : InMux
    port map (
            O => \N__29860\,
            I => \N__29855\
        );

    \I__5361\ : LocalMux
    port map (
            O => \N__29855\,
            I => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\
        );

    \I__5360\ : InMux
    port map (
            O => \N__29852\,
            I => \N__29849\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__29849\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\
        );

    \I__5358\ : CascadeMux
    port map (
            O => \N__29846\,
            I => \N__29842\
        );

    \I__5357\ : CascadeMux
    port map (
            O => \N__29845\,
            I => \N__29839\
        );

    \I__5356\ : InMux
    port map (
            O => \N__29842\,
            I => \N__29835\
        );

    \I__5355\ : InMux
    port map (
            O => \N__29839\,
            I => \N__29832\
        );

    \I__5354\ : InMux
    port map (
            O => \N__29838\,
            I => \N__29829\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__29835\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__29832\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__29829\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__5350\ : InMux
    port map (
            O => \N__29822\,
            I => \N__29818\
        );

    \I__5349\ : InMux
    port map (
            O => \N__29821\,
            I => \N__29815\
        );

    \I__5348\ : LocalMux
    port map (
            O => \N__29818\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__5347\ : LocalMux
    port map (
            O => \N__29815\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__5346\ : InMux
    port map (
            O => \N__29810\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\
        );

    \I__5345\ : InMux
    port map (
            O => \N__29807\,
            I => \N__29802\
        );

    \I__5344\ : InMux
    port map (
            O => \N__29806\,
            I => \N__29799\
        );

    \I__5343\ : InMux
    port map (
            O => \N__29805\,
            I => \N__29796\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__29802\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__29799\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__5340\ : LocalMux
    port map (
            O => \N__29796\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__5339\ : InMux
    port map (
            O => \N__29789\,
            I => \pwm_generator_inst.counter_cry_5\
        );

    \I__5338\ : InMux
    port map (
            O => \N__29786\,
            I => \pwm_generator_inst.counter_cry_6\
        );

    \I__5337\ : InMux
    port map (
            O => \N__29783\,
            I => \bfn_10_25_0_\
        );

    \I__5336\ : InMux
    port map (
            O => \N__29780\,
            I => \N__29766\
        );

    \I__5335\ : InMux
    port map (
            O => \N__29779\,
            I => \N__29766\
        );

    \I__5334\ : InMux
    port map (
            O => \N__29778\,
            I => \N__29757\
        );

    \I__5333\ : InMux
    port map (
            O => \N__29777\,
            I => \N__29757\
        );

    \I__5332\ : InMux
    port map (
            O => \N__29776\,
            I => \N__29757\
        );

    \I__5331\ : InMux
    port map (
            O => \N__29775\,
            I => \N__29757\
        );

    \I__5330\ : InMux
    port map (
            O => \N__29774\,
            I => \N__29748\
        );

    \I__5329\ : InMux
    port map (
            O => \N__29773\,
            I => \N__29748\
        );

    \I__5328\ : InMux
    port map (
            O => \N__29772\,
            I => \N__29748\
        );

    \I__5327\ : InMux
    port map (
            O => \N__29771\,
            I => \N__29748\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__29766\,
            I => \N__29745\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__29757\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__29748\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__5323\ : Odrv4
    port map (
            O => \N__29745\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__5322\ : InMux
    port map (
            O => \N__29738\,
            I => \pwm_generator_inst.counter_cry_8\
        );

    \I__5321\ : InMux
    port map (
            O => \N__29735\,
            I => \N__29731\
        );

    \I__5320\ : InMux
    port map (
            O => \N__29734\,
            I => \N__29727\
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__29731\,
            I => \N__29724\
        );

    \I__5318\ : InMux
    port map (
            O => \N__29730\,
            I => \N__29721\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__29727\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16\
        );

    \I__5316\ : Odrv4
    port map (
            O => \N__29724\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__29721\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16\
        );

    \I__5314\ : InMux
    port map (
            O => \N__29714\,
            I => \N__29710\
        );

    \I__5313\ : InMux
    port map (
            O => \N__29713\,
            I => \N__29707\
        );

    \I__5312\ : LocalMux
    port map (
            O => \N__29710\,
            I => \N__29703\
        );

    \I__5311\ : LocalMux
    port map (
            O => \N__29707\,
            I => \N__29700\
        );

    \I__5310\ : InMux
    port map (
            O => \N__29706\,
            I => \N__29697\
        );

    \I__5309\ : Span4Mux_h
    port map (
            O => \N__29703\,
            I => \N__29693\
        );

    \I__5308\ : Sp12to4
    port map (
            O => \N__29700\,
            I => \N__29688\
        );

    \I__5307\ : LocalMux
    port map (
            O => \N__29697\,
            I => \N__29688\
        );

    \I__5306\ : CascadeMux
    port map (
            O => \N__29696\,
            I => \N__29685\
        );

    \I__5305\ : Span4Mux_v
    port map (
            O => \N__29693\,
            I => \N__29682\
        );

    \I__5304\ : Span12Mux_s5_v
    port map (
            O => \N__29688\,
            I => \N__29679\
        );

    \I__5303\ : InMux
    port map (
            O => \N__29685\,
            I => \N__29676\
        );

    \I__5302\ : Odrv4
    port map (
            O => \N__29682\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__5301\ : Odrv12
    port map (
            O => \N__29679\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__29676\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__5299\ : CascadeMux
    port map (
            O => \N__29669\,
            I => \N__29666\
        );

    \I__5298\ : InMux
    port map (
            O => \N__29666\,
            I => \N__29663\
        );

    \I__5297\ : LocalMux
    port map (
            O => \N__29663\,
            I => \N__29660\
        );

    \I__5296\ : Span4Mux_h
    port map (
            O => \N__29660\,
            I => \N__29657\
        );

    \I__5295\ : Odrv4
    port map (
            O => \N__29657\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt16\
        );

    \I__5294\ : InMux
    port map (
            O => \N__29654\,
            I => \N__29648\
        );

    \I__5293\ : InMux
    port map (
            O => \N__29653\,
            I => \N__29648\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__29648\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\
        );

    \I__5291\ : InMux
    port map (
            O => \N__29645\,
            I => \N__29641\
        );

    \I__5290\ : InMux
    port map (
            O => \N__29644\,
            I => \N__29638\
        );

    \I__5289\ : LocalMux
    port map (
            O => \N__29641\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__29638\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\
        );

    \I__5287\ : InMux
    port map (
            O => \N__29633\,
            I => \N__29630\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__29630\,
            I => \N__29627\
        );

    \I__5285\ : Odrv4
    port map (
            O => \N__29627\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\
        );

    \I__5284\ : InMux
    port map (
            O => \N__29624\,
            I => \N__29621\
        );

    \I__5283\ : LocalMux
    port map (
            O => \N__29621\,
            I => \N__29616\
        );

    \I__5282\ : InMux
    port map (
            O => \N__29620\,
            I => \N__29611\
        );

    \I__5281\ : InMux
    port map (
            O => \N__29619\,
            I => \N__29611\
        );

    \I__5280\ : Span4Mux_v
    port map (
            O => \N__29616\,
            I => \N__29608\
        );

    \I__5279\ : LocalMux
    port map (
            O => \N__29611\,
            I => \N__29605\
        );

    \I__5278\ : Span4Mux_v
    port map (
            O => \N__29608\,
            I => \N__29601\
        );

    \I__5277\ : Sp12to4
    port map (
            O => \N__29605\,
            I => \N__29598\
        );

    \I__5276\ : InMux
    port map (
            O => \N__29604\,
            I => \N__29595\
        );

    \I__5275\ : Odrv4
    port map (
            O => \N__29601\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__5274\ : Odrv12
    port map (
            O => \N__29598\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__5273\ : LocalMux
    port map (
            O => \N__29595\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__5272\ : InMux
    port map (
            O => \N__29588\,
            I => \N__29585\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__29585\,
            I => \N__29581\
        );

    \I__5270\ : InMux
    port map (
            O => \N__29584\,
            I => \N__29578\
        );

    \I__5269\ : Odrv12
    port map (
            O => \N__29581\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15\
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__29578\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15\
        );

    \I__5267\ : InMux
    port map (
            O => \N__29573\,
            I => \N__29570\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__29570\,
            I => \N__29567\
        );

    \I__5265\ : Odrv4
    port map (
            O => \N__29567\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\
        );

    \I__5264\ : CascadeMux
    port map (
            O => \N__29564\,
            I => \pwm_generator_inst.un1_counterlto2_0_cascade_\
        );

    \I__5263\ : CascadeMux
    port map (
            O => \N__29561\,
            I => \pwm_generator_inst.un1_counterlt9_cascade_\
        );

    \I__5262\ : InMux
    port map (
            O => \N__29558\,
            I => \N__29553\
        );

    \I__5261\ : InMux
    port map (
            O => \N__29557\,
            I => \N__29550\
        );

    \I__5260\ : InMux
    port map (
            O => \N__29556\,
            I => \N__29547\
        );

    \I__5259\ : LocalMux
    port map (
            O => \N__29553\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__5258\ : LocalMux
    port map (
            O => \N__29550\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__29547\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__5256\ : InMux
    port map (
            O => \N__29540\,
            I => \bfn_10_24_0_\
        );

    \I__5255\ : InMux
    port map (
            O => \N__29537\,
            I => \N__29532\
        );

    \I__5254\ : InMux
    port map (
            O => \N__29536\,
            I => \N__29529\
        );

    \I__5253\ : InMux
    port map (
            O => \N__29535\,
            I => \N__29526\
        );

    \I__5252\ : LocalMux
    port map (
            O => \N__29532\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__29529\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__5250\ : LocalMux
    port map (
            O => \N__29526\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__5249\ : InMux
    port map (
            O => \N__29519\,
            I => \pwm_generator_inst.counter_cry_0\
        );

    \I__5248\ : InMux
    port map (
            O => \N__29516\,
            I => \N__29511\
        );

    \I__5247\ : InMux
    port map (
            O => \N__29515\,
            I => \N__29508\
        );

    \I__5246\ : InMux
    port map (
            O => \N__29514\,
            I => \N__29505\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__29511\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__29508\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__5243\ : LocalMux
    port map (
            O => \N__29505\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__5242\ : InMux
    port map (
            O => \N__29498\,
            I => \pwm_generator_inst.counter_cry_1\
        );

    \I__5241\ : InMux
    port map (
            O => \N__29495\,
            I => \N__29490\
        );

    \I__5240\ : InMux
    port map (
            O => \N__29494\,
            I => \N__29487\
        );

    \I__5239\ : InMux
    port map (
            O => \N__29493\,
            I => \N__29484\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__29490\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__5237\ : LocalMux
    port map (
            O => \N__29487\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__5236\ : LocalMux
    port map (
            O => \N__29484\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__5235\ : InMux
    port map (
            O => \N__29477\,
            I => \pwm_generator_inst.counter_cry_2\
        );

    \I__5234\ : InMux
    port map (
            O => \N__29474\,
            I => \N__29469\
        );

    \I__5233\ : InMux
    port map (
            O => \N__29473\,
            I => \N__29466\
        );

    \I__5232\ : InMux
    port map (
            O => \N__29472\,
            I => \N__29463\
        );

    \I__5231\ : LocalMux
    port map (
            O => \N__29469\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__29466\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__29463\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__5228\ : InMux
    port map (
            O => \N__29456\,
            I => \pwm_generator_inst.counter_cry_3\
        );

    \I__5227\ : InMux
    port map (
            O => \N__29453\,
            I => \N__29448\
        );

    \I__5226\ : InMux
    port map (
            O => \N__29452\,
            I => \N__29445\
        );

    \I__5225\ : InMux
    port map (
            O => \N__29451\,
            I => \N__29442\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__29448\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__29445\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__29442\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__5221\ : InMux
    port map (
            O => \N__29435\,
            I => \pwm_generator_inst.counter_cry_4\
        );

    \I__5220\ : InMux
    port map (
            O => \N__29432\,
            I => \N__29429\
        );

    \I__5219\ : LocalMux
    port map (
            O => \N__29429\,
            I => \N__29425\
        );

    \I__5218\ : InMux
    port map (
            O => \N__29428\,
            I => \N__29421\
        );

    \I__5217\ : Span4Mux_h
    port map (
            O => \N__29425\,
            I => \N__29418\
        );

    \I__5216\ : InMux
    port map (
            O => \N__29424\,
            I => \N__29415\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__29421\,
            I => \elapsed_time_ns_1_RNIK63T9_0_8\
        );

    \I__5214\ : Odrv4
    port map (
            O => \N__29418\,
            I => \elapsed_time_ns_1_RNIK63T9_0_8\
        );

    \I__5213\ : LocalMux
    port map (
            O => \N__29415\,
            I => \elapsed_time_ns_1_RNIK63T9_0_8\
        );

    \I__5212\ : InMux
    port map (
            O => \N__29408\,
            I => \N__29404\
        );

    \I__5211\ : InMux
    port map (
            O => \N__29407\,
            I => \N__29401\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__29404\,
            I => \N__29397\
        );

    \I__5209\ : LocalMux
    port map (
            O => \N__29401\,
            I => \N__29393\
        );

    \I__5208\ : InMux
    port map (
            O => \N__29400\,
            I => \N__29390\
        );

    \I__5207\ : Span4Mux_v
    port map (
            O => \N__29397\,
            I => \N__29387\
        );

    \I__5206\ : InMux
    port map (
            O => \N__29396\,
            I => \N__29384\
        );

    \I__5205\ : Span4Mux_v
    port map (
            O => \N__29393\,
            I => \N__29379\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__29390\,
            I => \N__29379\
        );

    \I__5203\ : Odrv4
    port map (
            O => \N__29387\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__29384\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__5201\ : Odrv4
    port map (
            O => \N__29379\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__5200\ : CascadeMux
    port map (
            O => \N__29372\,
            I => \N__29369\
        );

    \I__5199\ : InMux
    port map (
            O => \N__29369\,
            I => \N__29366\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__29366\,
            I => \N__29363\
        );

    \I__5197\ : Span12Mux_v
    port map (
            O => \N__29363\,
            I => \N__29360\
        );

    \I__5196\ : Odrv12
    port map (
            O => \N__29360\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\
        );

    \I__5195\ : CEMux
    port map (
            O => \N__29357\,
            I => \N__29353\
        );

    \I__5194\ : CEMux
    port map (
            O => \N__29356\,
            I => \N__29350\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__29353\,
            I => \N__29345\
        );

    \I__5192\ : LocalMux
    port map (
            O => \N__29350\,
            I => \N__29342\
        );

    \I__5191\ : CEMux
    port map (
            O => \N__29349\,
            I => \N__29339\
        );

    \I__5190\ : CEMux
    port map (
            O => \N__29348\,
            I => \N__29336\
        );

    \I__5189\ : Span4Mux_v
    port map (
            O => \N__29345\,
            I => \N__29331\
        );

    \I__5188\ : Span4Mux_v
    port map (
            O => \N__29342\,
            I => \N__29331\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__29339\,
            I => \N__29326\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__29336\,
            I => \N__29326\
        );

    \I__5185\ : Span4Mux_h
    port map (
            O => \N__29331\,
            I => \N__29321\
        );

    \I__5184\ : Span4Mux_v
    port map (
            O => \N__29326\,
            I => \N__29321\
        );

    \I__5183\ : Odrv4
    port map (
            O => \N__29321\,
            I => \delay_measurement_inst.delay_hc_timer.N_203_i\
        );

    \I__5182\ : InMux
    port map (
            O => \N__29318\,
            I => \N__29315\
        );

    \I__5181\ : LocalMux
    port map (
            O => \N__29315\,
            I => \N__29312\
        );

    \I__5180\ : Span4Mux_h
    port map (
            O => \N__29312\,
            I => \N__29309\
        );

    \I__5179\ : Sp12to4
    port map (
            O => \N__29309\,
            I => \N__29306\
        );

    \I__5178\ : Span12Mux_v
    port map (
            O => \N__29306\,
            I => \N__29303\
        );

    \I__5177\ : Odrv12
    port map (
            O => \N__29303\,
            I => \il_max_comp1_D1\
        );

    \I__5176\ : InMux
    port map (
            O => \N__29300\,
            I => \N__29296\
        );

    \I__5175\ : InMux
    port map (
            O => \N__29299\,
            I => \N__29293\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__29296\,
            I => \N__29290\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__29293\,
            I => \N__29287\
        );

    \I__5172\ : Span4Mux_h
    port map (
            O => \N__29290\,
            I => \N__29282\
        );

    \I__5171\ : Span4Mux_v
    port map (
            O => \N__29287\,
            I => \N__29282\
        );

    \I__5170\ : Odrv4
    port map (
            O => \N__29282\,
            I => \current_shift_inst.control_input_axb_0\
        );

    \I__5169\ : InMux
    port map (
            O => \N__29279\,
            I => \N__29271\
        );

    \I__5168\ : InMux
    port map (
            O => \N__29278\,
            I => \N__29271\
        );

    \I__5167\ : InMux
    port map (
            O => \N__29277\,
            I => \N__29268\
        );

    \I__5166\ : InMux
    port map (
            O => \N__29276\,
            I => \N__29265\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__29271\,
            I => \N__29262\
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__29268\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__5163\ : LocalMux
    port map (
            O => \N__29265\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__5162\ : Odrv12
    port map (
            O => \N__29262\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__5161\ : InMux
    port map (
            O => \N__29255\,
            I => \N__29239\
        );

    \I__5160\ : InMux
    port map (
            O => \N__29254\,
            I => \N__29239\
        );

    \I__5159\ : InMux
    port map (
            O => \N__29253\,
            I => \N__29239\
        );

    \I__5158\ : InMux
    port map (
            O => \N__29252\,
            I => \N__29239\
        );

    \I__5157\ : InMux
    port map (
            O => \N__29251\,
            I => \N__29208\
        );

    \I__5156\ : InMux
    port map (
            O => \N__29250\,
            I => \N__29208\
        );

    \I__5155\ : InMux
    port map (
            O => \N__29249\,
            I => \N__29208\
        );

    \I__5154\ : InMux
    port map (
            O => \N__29248\,
            I => \N__29208\
        );

    \I__5153\ : LocalMux
    port map (
            O => \N__29239\,
            I => \N__29205\
        );

    \I__5152\ : InMux
    port map (
            O => \N__29238\,
            I => \N__29196\
        );

    \I__5151\ : InMux
    port map (
            O => \N__29237\,
            I => \N__29196\
        );

    \I__5150\ : InMux
    port map (
            O => \N__29236\,
            I => \N__29196\
        );

    \I__5149\ : InMux
    port map (
            O => \N__29235\,
            I => \N__29196\
        );

    \I__5148\ : InMux
    port map (
            O => \N__29234\,
            I => \N__29191\
        );

    \I__5147\ : InMux
    port map (
            O => \N__29233\,
            I => \N__29191\
        );

    \I__5146\ : InMux
    port map (
            O => \N__29232\,
            I => \N__29182\
        );

    \I__5145\ : InMux
    port map (
            O => \N__29231\,
            I => \N__29182\
        );

    \I__5144\ : InMux
    port map (
            O => \N__29230\,
            I => \N__29182\
        );

    \I__5143\ : InMux
    port map (
            O => \N__29229\,
            I => \N__29182\
        );

    \I__5142\ : InMux
    port map (
            O => \N__29228\,
            I => \N__29173\
        );

    \I__5141\ : InMux
    port map (
            O => \N__29227\,
            I => \N__29173\
        );

    \I__5140\ : InMux
    port map (
            O => \N__29226\,
            I => \N__29173\
        );

    \I__5139\ : InMux
    port map (
            O => \N__29225\,
            I => \N__29173\
        );

    \I__5138\ : InMux
    port map (
            O => \N__29224\,
            I => \N__29164\
        );

    \I__5137\ : InMux
    port map (
            O => \N__29223\,
            I => \N__29164\
        );

    \I__5136\ : InMux
    port map (
            O => \N__29222\,
            I => \N__29164\
        );

    \I__5135\ : InMux
    port map (
            O => \N__29221\,
            I => \N__29164\
        );

    \I__5134\ : InMux
    port map (
            O => \N__29220\,
            I => \N__29155\
        );

    \I__5133\ : InMux
    port map (
            O => \N__29219\,
            I => \N__29155\
        );

    \I__5132\ : InMux
    port map (
            O => \N__29218\,
            I => \N__29155\
        );

    \I__5131\ : InMux
    port map (
            O => \N__29217\,
            I => \N__29155\
        );

    \I__5130\ : LocalMux
    port map (
            O => \N__29208\,
            I => \N__29150\
        );

    \I__5129\ : Span4Mux_v
    port map (
            O => \N__29205\,
            I => \N__29150\
        );

    \I__5128\ : LocalMux
    port map (
            O => \N__29196\,
            I => \N__29147\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__29191\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__5126\ : LocalMux
    port map (
            O => \N__29182\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__29173\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__29164\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__5123\ : LocalMux
    port map (
            O => \N__29155\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__5122\ : Odrv4
    port map (
            O => \N__29150\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__5121\ : Odrv4
    port map (
            O => \N__29147\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__5120\ : InMux
    port map (
            O => \N__29132\,
            I => \N__29129\
        );

    \I__5119\ : LocalMux
    port map (
            O => \N__29129\,
            I => \current_shift_inst.control_input_axb_12\
        );

    \I__5118\ : InMux
    port map (
            O => \N__29126\,
            I => \N__29123\
        );

    \I__5117\ : LocalMux
    port map (
            O => \N__29123\,
            I => \N__29119\
        );

    \I__5116\ : CascadeMux
    port map (
            O => \N__29122\,
            I => \N__29115\
        );

    \I__5115\ : Span4Mux_v
    port map (
            O => \N__29119\,
            I => \N__29112\
        );

    \I__5114\ : InMux
    port map (
            O => \N__29118\,
            I => \N__29109\
        );

    \I__5113\ : InMux
    port map (
            O => \N__29115\,
            I => \N__29106\
        );

    \I__5112\ : Odrv4
    port map (
            O => \N__29112\,
            I => \current_shift_inst.N_1304_i\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__29109\,
            I => \current_shift_inst.N_1304_i\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__29106\,
            I => \current_shift_inst.N_1304_i\
        );

    \I__5109\ : CascadeMux
    port map (
            O => \N__29099\,
            I => \N__29096\
        );

    \I__5108\ : InMux
    port map (
            O => \N__29096\,
            I => \N__29091\
        );

    \I__5107\ : InMux
    port map (
            O => \N__29095\,
            I => \N__29088\
        );

    \I__5106\ : InMux
    port map (
            O => \N__29094\,
            I => \N__29085\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__29091\,
            I => \N__29080\
        );

    \I__5104\ : LocalMux
    port map (
            O => \N__29088\,
            I => \N__29080\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__29085\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__5102\ : Odrv4
    port map (
            O => \N__29080\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__5101\ : InMux
    port map (
            O => \N__29075\,
            I => \N__29071\
        );

    \I__5100\ : InMux
    port map (
            O => \N__29074\,
            I => \N__29068\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__29071\,
            I => \N__29065\
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__29068\,
            I => \N__29062\
        );

    \I__5097\ : Span4Mux_h
    port map (
            O => \N__29065\,
            I => \N__29057\
        );

    \I__5096\ : Span4Mux_v
    port map (
            O => \N__29062\,
            I => \N__29057\
        );

    \I__5095\ : Span4Mux_v
    port map (
            O => \N__29057\,
            I => \N__29052\
        );

    \I__5094\ : InMux
    port map (
            O => \N__29056\,
            I => \N__29049\
        );

    \I__5093\ : InMux
    port map (
            O => \N__29055\,
            I => \N__29046\
        );

    \I__5092\ : Odrv4
    port map (
            O => \N__29052\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__29049\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__29046\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__5089\ : InMux
    port map (
            O => \N__29039\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__5088\ : CascadeMux
    port map (
            O => \N__29036\,
            I => \N__29033\
        );

    \I__5087\ : InMux
    port map (
            O => \N__29033\,
            I => \N__29029\
        );

    \I__5086\ : InMux
    port map (
            O => \N__29032\,
            I => \N__29026\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__29029\,
            I => \N__29020\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__29026\,
            I => \N__29020\
        );

    \I__5083\ : InMux
    port map (
            O => \N__29025\,
            I => \N__29017\
        );

    \I__5082\ : Span4Mux_h
    port map (
            O => \N__29020\,
            I => \N__29014\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__29017\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__5080\ : Odrv4
    port map (
            O => \N__29014\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__5079\ : InMux
    port map (
            O => \N__29009\,
            I => \N__29004\
        );

    \I__5078\ : InMux
    port map (
            O => \N__29008\,
            I => \N__29001\
        );

    \I__5077\ : InMux
    port map (
            O => \N__29007\,
            I => \N__28998\
        );

    \I__5076\ : LocalMux
    port map (
            O => \N__29004\,
            I => \N__28995\
        );

    \I__5075\ : LocalMux
    port map (
            O => \N__29001\,
            I => \N__28992\
        );

    \I__5074\ : LocalMux
    port map (
            O => \N__28998\,
            I => \N__28989\
        );

    \I__5073\ : Span4Mux_h
    port map (
            O => \N__28995\,
            I => \N__28984\
        );

    \I__5072\ : Span4Mux_h
    port map (
            O => \N__28992\,
            I => \N__28984\
        );

    \I__5071\ : Span12Mux_s10_h
    port map (
            O => \N__28989\,
            I => \N__28978\
        );

    \I__5070\ : Sp12to4
    port map (
            O => \N__28984\,
            I => \N__28978\
        );

    \I__5069\ : InMux
    port map (
            O => \N__28983\,
            I => \N__28975\
        );

    \I__5068\ : Odrv12
    port map (
            O => \N__28978\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__5067\ : LocalMux
    port map (
            O => \N__28975\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__5066\ : InMux
    port map (
            O => \N__28970\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__5065\ : CascadeMux
    port map (
            O => \N__28967\,
            I => \N__28964\
        );

    \I__5064\ : InMux
    port map (
            O => \N__28964\,
            I => \N__28960\
        );

    \I__5063\ : InMux
    port map (
            O => \N__28963\,
            I => \N__28957\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__28960\,
            I => \N__28951\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__28957\,
            I => \N__28951\
        );

    \I__5060\ : InMux
    port map (
            O => \N__28956\,
            I => \N__28948\
        );

    \I__5059\ : Span4Mux_h
    port map (
            O => \N__28951\,
            I => \N__28945\
        );

    \I__5058\ : LocalMux
    port map (
            O => \N__28948\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__5057\ : Odrv4
    port map (
            O => \N__28945\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__5056\ : InMux
    port map (
            O => \N__28940\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__5055\ : CascadeMux
    port map (
            O => \N__28937\,
            I => \N__28934\
        );

    \I__5054\ : InMux
    port map (
            O => \N__28934\,
            I => \N__28930\
        );

    \I__5053\ : InMux
    port map (
            O => \N__28933\,
            I => \N__28927\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__28930\,
            I => \N__28923\
        );

    \I__5051\ : LocalMux
    port map (
            O => \N__28927\,
            I => \N__28920\
        );

    \I__5050\ : InMux
    port map (
            O => \N__28926\,
            I => \N__28917\
        );

    \I__5049\ : Span4Mux_h
    port map (
            O => \N__28923\,
            I => \N__28914\
        );

    \I__5048\ : Span4Mux_h
    port map (
            O => \N__28920\,
            I => \N__28911\
        );

    \I__5047\ : LocalMux
    port map (
            O => \N__28917\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__5046\ : Odrv4
    port map (
            O => \N__28914\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__5045\ : Odrv4
    port map (
            O => \N__28911\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__5044\ : InMux
    port map (
            O => \N__28904\,
            I => \N__28896\
        );

    \I__5043\ : InMux
    port map (
            O => \N__28903\,
            I => \N__28896\
        );

    \I__5042\ : InMux
    port map (
            O => \N__28902\,
            I => \N__28893\
        );

    \I__5041\ : InMux
    port map (
            O => \N__28901\,
            I => \N__28890\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__28896\,
            I => \N__28885\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__28893\,
            I => \N__28885\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__28890\,
            I => \N__28882\
        );

    \I__5037\ : Span4Mux_h
    port map (
            O => \N__28885\,
            I => \N__28879\
        );

    \I__5036\ : Odrv12
    port map (
            O => \N__28882\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__5035\ : Odrv4
    port map (
            O => \N__28879\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__5034\ : InMux
    port map (
            O => \N__28874\,
            I => \bfn_10_15_0_\
        );

    \I__5033\ : InMux
    port map (
            O => \N__28871\,
            I => \N__28867\
        );

    \I__5032\ : InMux
    port map (
            O => \N__28870\,
            I => \N__28864\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__28867\,
            I => \N__28860\
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__28864\,
            I => \N__28857\
        );

    \I__5029\ : InMux
    port map (
            O => \N__28863\,
            I => \N__28854\
        );

    \I__5028\ : Span4Mux_h
    port map (
            O => \N__28860\,
            I => \N__28851\
        );

    \I__5027\ : Odrv4
    port map (
            O => \N__28857\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__28854\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__5025\ : Odrv4
    port map (
            O => \N__28851\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__5024\ : InMux
    port map (
            O => \N__28844\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__5023\ : InMux
    port map (
            O => \N__28841\,
            I => \N__28834\
        );

    \I__5022\ : InMux
    port map (
            O => \N__28840\,
            I => \N__28834\
        );

    \I__5021\ : InMux
    port map (
            O => \N__28839\,
            I => \N__28831\
        );

    \I__5020\ : LocalMux
    port map (
            O => \N__28834\,
            I => \N__28828\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__28831\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__5018\ : Odrv4
    port map (
            O => \N__28828\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__5017\ : CascadeMux
    port map (
            O => \N__28823\,
            I => \N__28820\
        );

    \I__5016\ : InMux
    port map (
            O => \N__28820\,
            I => \N__28816\
        );

    \I__5015\ : InMux
    port map (
            O => \N__28819\,
            I => \N__28813\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__28816\,
            I => \N__28810\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__28813\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__5012\ : Odrv4
    port map (
            O => \N__28810\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__5011\ : InMux
    port map (
            O => \N__28805\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__5010\ : InMux
    port map (
            O => \N__28802\,
            I => \N__28799\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__28799\,
            I => \N__28795\
        );

    \I__5008\ : InMux
    port map (
            O => \N__28798\,
            I => \N__28792\
        );

    \I__5007\ : Span4Mux_v
    port map (
            O => \N__28795\,
            I => \N__28789\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__28792\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__5005\ : Odrv4
    port map (
            O => \N__28789\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__5004\ : CascadeMux
    port map (
            O => \N__28784\,
            I => \N__28779\
        );

    \I__5003\ : CascadeMux
    port map (
            O => \N__28783\,
            I => \N__28776\
        );

    \I__5002\ : InMux
    port map (
            O => \N__28782\,
            I => \N__28773\
        );

    \I__5001\ : InMux
    port map (
            O => \N__28779\,
            I => \N__28768\
        );

    \I__5000\ : InMux
    port map (
            O => \N__28776\,
            I => \N__28768\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__28773\,
            I => \N__28763\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__28768\,
            I => \N__28763\
        );

    \I__4997\ : Odrv4
    port map (
            O => \N__28763\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__4996\ : InMux
    port map (
            O => \N__28760\,
            I => \N__28755\
        );

    \I__4995\ : InMux
    port map (
            O => \N__28759\,
            I => \N__28752\
        );

    \I__4994\ : CascadeMux
    port map (
            O => \N__28758\,
            I => \N__28749\
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__28755\,
            I => \N__28746\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__28752\,
            I => \N__28743\
        );

    \I__4991\ : InMux
    port map (
            O => \N__28749\,
            I => \N__28740\
        );

    \I__4990\ : Span4Mux_h
    port map (
            O => \N__28746\,
            I => \N__28732\
        );

    \I__4989\ : Span4Mux_h
    port map (
            O => \N__28743\,
            I => \N__28732\
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__28740\,
            I => \N__28732\
        );

    \I__4987\ : InMux
    port map (
            O => \N__28739\,
            I => \N__28729\
        );

    \I__4986\ : Odrv4
    port map (
            O => \N__28732\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__4985\ : LocalMux
    port map (
            O => \N__28729\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__4984\ : InMux
    port map (
            O => \N__28724\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__4983\ : InMux
    port map (
            O => \N__28721\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__4982\ : InMux
    port map (
            O => \N__28718\,
            I => \N__28714\
        );

    \I__4981\ : InMux
    port map (
            O => \N__28717\,
            I => \N__28711\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__28714\,
            I => \N__28706\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__28711\,
            I => \N__28703\
        );

    \I__4978\ : InMux
    port map (
            O => \N__28710\,
            I => \N__28698\
        );

    \I__4977\ : InMux
    port map (
            O => \N__28709\,
            I => \N__28698\
        );

    \I__4976\ : Span4Mux_h
    port map (
            O => \N__28706\,
            I => \N__28695\
        );

    \I__4975\ : Span4Mux_v
    port map (
            O => \N__28703\,
            I => \N__28690\
        );

    \I__4974\ : LocalMux
    port map (
            O => \N__28698\,
            I => \N__28690\
        );

    \I__4973\ : Odrv4
    port map (
            O => \N__28695\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__4972\ : Odrv4
    port map (
            O => \N__28690\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__4971\ : CEMux
    port map (
            O => \N__28685\,
            I => \N__28680\
        );

    \I__4970\ : CEMux
    port map (
            O => \N__28684\,
            I => \N__28677\
        );

    \I__4969\ : CEMux
    port map (
            O => \N__28683\,
            I => \N__28672\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__28680\,
            I => \N__28668\
        );

    \I__4967\ : LocalMux
    port map (
            O => \N__28677\,
            I => \N__28665\
        );

    \I__4966\ : CEMux
    port map (
            O => \N__28676\,
            I => \N__28662\
        );

    \I__4965\ : CEMux
    port map (
            O => \N__28675\,
            I => \N__28659\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__28672\,
            I => \N__28656\
        );

    \I__4963\ : CEMux
    port map (
            O => \N__28671\,
            I => \N__28653\
        );

    \I__4962\ : Span4Mux_v
    port map (
            O => \N__28668\,
            I => \N__28650\
        );

    \I__4961\ : Span4Mux_h
    port map (
            O => \N__28665\,
            I => \N__28645\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__28662\,
            I => \N__28645\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__28659\,
            I => \N__28638\
        );

    \I__4958\ : Span4Mux_v
    port map (
            O => \N__28656\,
            I => \N__28638\
        );

    \I__4957\ : LocalMux
    port map (
            O => \N__28653\,
            I => \N__28638\
        );

    \I__4956\ : Span4Mux_h
    port map (
            O => \N__28650\,
            I => \N__28633\
        );

    \I__4955\ : Span4Mux_v
    port map (
            O => \N__28645\,
            I => \N__28633\
        );

    \I__4954\ : Span4Mux_h
    port map (
            O => \N__28638\,
            I => \N__28630\
        );

    \I__4953\ : Odrv4
    port map (
            O => \N__28633\,
            I => \delay_measurement_inst.delay_hc_timer.N_202_i\
        );

    \I__4952\ : Odrv4
    port map (
            O => \N__28630\,
            I => \delay_measurement_inst.delay_hc_timer.N_202_i\
        );

    \I__4951\ : CascadeMux
    port map (
            O => \N__28625\,
            I => \N__28621\
        );

    \I__4950\ : CascadeMux
    port map (
            O => \N__28624\,
            I => \N__28618\
        );

    \I__4949\ : InMux
    port map (
            O => \N__28621\,
            I => \N__28612\
        );

    \I__4948\ : InMux
    port map (
            O => \N__28618\,
            I => \N__28612\
        );

    \I__4947\ : InMux
    port map (
            O => \N__28617\,
            I => \N__28609\
        );

    \I__4946\ : LocalMux
    port map (
            O => \N__28612\,
            I => \N__28606\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__28609\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__4944\ : Odrv4
    port map (
            O => \N__28606\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__4943\ : InMux
    port map (
            O => \N__28601\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__4942\ : CascadeMux
    port map (
            O => \N__28598\,
            I => \N__28595\
        );

    \I__4941\ : InMux
    port map (
            O => \N__28595\,
            I => \N__28591\
        );

    \I__4940\ : InMux
    port map (
            O => \N__28594\,
            I => \N__28588\
        );

    \I__4939\ : LocalMux
    port map (
            O => \N__28591\,
            I => \N__28582\
        );

    \I__4938\ : LocalMux
    port map (
            O => \N__28588\,
            I => \N__28582\
        );

    \I__4937\ : InMux
    port map (
            O => \N__28587\,
            I => \N__28579\
        );

    \I__4936\ : Span4Mux_h
    port map (
            O => \N__28582\,
            I => \N__28576\
        );

    \I__4935\ : LocalMux
    port map (
            O => \N__28579\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__4934\ : Odrv4
    port map (
            O => \N__28576\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__4933\ : InMux
    port map (
            O => \N__28571\,
            I => \N__28566\
        );

    \I__4932\ : InMux
    port map (
            O => \N__28570\,
            I => \N__28563\
        );

    \I__4931\ : InMux
    port map (
            O => \N__28569\,
            I => \N__28560\
        );

    \I__4930\ : LocalMux
    port map (
            O => \N__28566\,
            I => \N__28557\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__28563\,
            I => \N__28552\
        );

    \I__4928\ : LocalMux
    port map (
            O => \N__28560\,
            I => \N__28552\
        );

    \I__4927\ : Span4Mux_v
    port map (
            O => \N__28557\,
            I => \N__28547\
        );

    \I__4926\ : Span4Mux_v
    port map (
            O => \N__28552\,
            I => \N__28547\
        );

    \I__4925\ : Span4Mux_v
    port map (
            O => \N__28547\,
            I => \N__28543\
        );

    \I__4924\ : InMux
    port map (
            O => \N__28546\,
            I => \N__28540\
        );

    \I__4923\ : Odrv4
    port map (
            O => \N__28543\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__4922\ : LocalMux
    port map (
            O => \N__28540\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__4921\ : InMux
    port map (
            O => \N__28535\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__4920\ : CascadeMux
    port map (
            O => \N__28532\,
            I => \N__28529\
        );

    \I__4919\ : InMux
    port map (
            O => \N__28529\,
            I => \N__28525\
        );

    \I__4918\ : InMux
    port map (
            O => \N__28528\,
            I => \N__28522\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__28525\,
            I => \N__28516\
        );

    \I__4916\ : LocalMux
    port map (
            O => \N__28522\,
            I => \N__28516\
        );

    \I__4915\ : InMux
    port map (
            O => \N__28521\,
            I => \N__28513\
        );

    \I__4914\ : Span4Mux_h
    port map (
            O => \N__28516\,
            I => \N__28510\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__28513\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__4912\ : Odrv4
    port map (
            O => \N__28510\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__4911\ : InMux
    port map (
            O => \N__28505\,
            I => \N__28500\
        );

    \I__4910\ : InMux
    port map (
            O => \N__28504\,
            I => \N__28495\
        );

    \I__4909\ : InMux
    port map (
            O => \N__28503\,
            I => \N__28495\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__28500\,
            I => \N__28492\
        );

    \I__4907\ : LocalMux
    port map (
            O => \N__28495\,
            I => \N__28489\
        );

    \I__4906\ : Span4Mux_h
    port map (
            O => \N__28492\,
            I => \N__28484\
        );

    \I__4905\ : Span4Mux_h
    port map (
            O => \N__28489\,
            I => \N__28484\
        );

    \I__4904\ : Span4Mux_v
    port map (
            O => \N__28484\,
            I => \N__28480\
        );

    \I__4903\ : InMux
    port map (
            O => \N__28483\,
            I => \N__28477\
        );

    \I__4902\ : Odrv4
    port map (
            O => \N__28480\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__28477\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__4900\ : InMux
    port map (
            O => \N__28472\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__4899\ : CascadeMux
    port map (
            O => \N__28469\,
            I => \N__28466\
        );

    \I__4898\ : InMux
    port map (
            O => \N__28466\,
            I => \N__28462\
        );

    \I__4897\ : InMux
    port map (
            O => \N__28465\,
            I => \N__28459\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__28462\,
            I => \N__28455\
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__28459\,
            I => \N__28452\
        );

    \I__4894\ : InMux
    port map (
            O => \N__28458\,
            I => \N__28449\
        );

    \I__4893\ : Span4Mux_h
    port map (
            O => \N__28455\,
            I => \N__28446\
        );

    \I__4892\ : Span4Mux_h
    port map (
            O => \N__28452\,
            I => \N__28443\
        );

    \I__4891\ : LocalMux
    port map (
            O => \N__28449\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__4890\ : Odrv4
    port map (
            O => \N__28446\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__4889\ : Odrv4
    port map (
            O => \N__28443\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__4888\ : InMux
    port map (
            O => \N__28436\,
            I => \N__28430\
        );

    \I__4887\ : InMux
    port map (
            O => \N__28435\,
            I => \N__28427\
        );

    \I__4886\ : CascadeMux
    port map (
            O => \N__28434\,
            I => \N__28424\
        );

    \I__4885\ : InMux
    port map (
            O => \N__28433\,
            I => \N__28421\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__28430\,
            I => \N__28418\
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__28427\,
            I => \N__28415\
        );

    \I__4882\ : InMux
    port map (
            O => \N__28424\,
            I => \N__28412\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__28421\,
            I => \N__28409\
        );

    \I__4880\ : Span4Mux_v
    port map (
            O => \N__28418\,
            I => \N__28404\
        );

    \I__4879\ : Span4Mux_h
    port map (
            O => \N__28415\,
            I => \N__28404\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__28412\,
            I => \N__28401\
        );

    \I__4877\ : Span4Mux_v
    port map (
            O => \N__28409\,
            I => \N__28396\
        );

    \I__4876\ : Span4Mux_v
    port map (
            O => \N__28404\,
            I => \N__28396\
        );

    \I__4875\ : Span4Mux_h
    port map (
            O => \N__28401\,
            I => \N__28393\
        );

    \I__4874\ : Odrv4
    port map (
            O => \N__28396\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__4873\ : Odrv4
    port map (
            O => \N__28393\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__4872\ : InMux
    port map (
            O => \N__28388\,
            I => \bfn_10_14_0_\
        );

    \I__4871\ : InMux
    port map (
            O => \N__28385\,
            I => \N__28381\
        );

    \I__4870\ : InMux
    port map (
            O => \N__28384\,
            I => \N__28378\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__28381\,
            I => \N__28374\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__28378\,
            I => \N__28371\
        );

    \I__4867\ : InMux
    port map (
            O => \N__28377\,
            I => \N__28368\
        );

    \I__4866\ : Span4Mux_h
    port map (
            O => \N__28374\,
            I => \N__28365\
        );

    \I__4865\ : Span4Mux_h
    port map (
            O => \N__28371\,
            I => \N__28362\
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__28368\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__4863\ : Odrv4
    port map (
            O => \N__28365\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__4862\ : Odrv4
    port map (
            O => \N__28362\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__4861\ : InMux
    port map (
            O => \N__28355\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__4860\ : InMux
    port map (
            O => \N__28352\,
            I => \N__28345\
        );

    \I__4859\ : InMux
    port map (
            O => \N__28351\,
            I => \N__28345\
        );

    \I__4858\ : InMux
    port map (
            O => \N__28350\,
            I => \N__28342\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__28345\,
            I => \N__28339\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__28342\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__4855\ : Odrv4
    port map (
            O => \N__28339\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__4854\ : InMux
    port map (
            O => \N__28334\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__4853\ : CascadeMux
    port map (
            O => \N__28331\,
            I => \N__28327\
        );

    \I__4852\ : CascadeMux
    port map (
            O => \N__28330\,
            I => \N__28324\
        );

    \I__4851\ : InMux
    port map (
            O => \N__28327\,
            I => \N__28318\
        );

    \I__4850\ : InMux
    port map (
            O => \N__28324\,
            I => \N__28318\
        );

    \I__4849\ : InMux
    port map (
            O => \N__28323\,
            I => \N__28315\
        );

    \I__4848\ : LocalMux
    port map (
            O => \N__28318\,
            I => \N__28312\
        );

    \I__4847\ : LocalMux
    port map (
            O => \N__28315\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__4846\ : Odrv4
    port map (
            O => \N__28312\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__4845\ : InMux
    port map (
            O => \N__28307\,
            I => \N__28302\
        );

    \I__4844\ : InMux
    port map (
            O => \N__28306\,
            I => \N__28297\
        );

    \I__4843\ : InMux
    port map (
            O => \N__28305\,
            I => \N__28297\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__28302\,
            I => \N__28291\
        );

    \I__4841\ : LocalMux
    port map (
            O => \N__28297\,
            I => \N__28291\
        );

    \I__4840\ : CascadeMux
    port map (
            O => \N__28296\,
            I => \N__28288\
        );

    \I__4839\ : Span4Mux_v
    port map (
            O => \N__28291\,
            I => \N__28285\
        );

    \I__4838\ : InMux
    port map (
            O => \N__28288\,
            I => \N__28282\
        );

    \I__4837\ : Odrv4
    port map (
            O => \N__28285\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__28282\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__4835\ : InMux
    port map (
            O => \N__28277\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__4834\ : CascadeMux
    port map (
            O => \N__28274\,
            I => \N__28270\
        );

    \I__4833\ : CascadeMux
    port map (
            O => \N__28273\,
            I => \N__28267\
        );

    \I__4832\ : InMux
    port map (
            O => \N__28270\,
            I => \N__28261\
        );

    \I__4831\ : InMux
    port map (
            O => \N__28267\,
            I => \N__28261\
        );

    \I__4830\ : InMux
    port map (
            O => \N__28266\,
            I => \N__28258\
        );

    \I__4829\ : LocalMux
    port map (
            O => \N__28261\,
            I => \N__28255\
        );

    \I__4828\ : LocalMux
    port map (
            O => \N__28258\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__4827\ : Odrv4
    port map (
            O => \N__28255\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__4826\ : InMux
    port map (
            O => \N__28250\,
            I => \N__28245\
        );

    \I__4825\ : InMux
    port map (
            O => \N__28249\,
            I => \N__28240\
        );

    \I__4824\ : InMux
    port map (
            O => \N__28248\,
            I => \N__28240\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__28245\,
            I => \N__28237\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__28240\,
            I => \N__28234\
        );

    \I__4821\ : Span4Mux_v
    port map (
            O => \N__28237\,
            I => \N__28230\
        );

    \I__4820\ : Sp12to4
    port map (
            O => \N__28234\,
            I => \N__28227\
        );

    \I__4819\ : InMux
    port map (
            O => \N__28233\,
            I => \N__28224\
        );

    \I__4818\ : Odrv4
    port map (
            O => \N__28230\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__4817\ : Odrv12
    port map (
            O => \N__28227\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__4816\ : LocalMux
    port map (
            O => \N__28224\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__4815\ : InMux
    port map (
            O => \N__28217\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__4814\ : CascadeMux
    port map (
            O => \N__28214\,
            I => \N__28210\
        );

    \I__4813\ : CascadeMux
    port map (
            O => \N__28213\,
            I => \N__28207\
        );

    \I__4812\ : InMux
    port map (
            O => \N__28210\,
            I => \N__28201\
        );

    \I__4811\ : InMux
    port map (
            O => \N__28207\,
            I => \N__28201\
        );

    \I__4810\ : InMux
    port map (
            O => \N__28206\,
            I => \N__28198\
        );

    \I__4809\ : LocalMux
    port map (
            O => \N__28201\,
            I => \N__28195\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__28198\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__4807\ : Odrv4
    port map (
            O => \N__28195\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__4806\ : InMux
    port map (
            O => \N__28190\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__4805\ : CascadeMux
    port map (
            O => \N__28187\,
            I => \N__28184\
        );

    \I__4804\ : InMux
    port map (
            O => \N__28184\,
            I => \N__28180\
        );

    \I__4803\ : InMux
    port map (
            O => \N__28183\,
            I => \N__28177\
        );

    \I__4802\ : LocalMux
    port map (
            O => \N__28180\,
            I => \N__28171\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__28177\,
            I => \N__28171\
        );

    \I__4800\ : InMux
    port map (
            O => \N__28176\,
            I => \N__28168\
        );

    \I__4799\ : Span4Mux_h
    port map (
            O => \N__28171\,
            I => \N__28165\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__28168\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__4797\ : Odrv4
    port map (
            O => \N__28165\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__4796\ : InMux
    port map (
            O => \N__28160\,
            I => \N__28157\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__28157\,
            I => \N__28151\
        );

    \I__4794\ : InMux
    port map (
            O => \N__28156\,
            I => \N__28144\
        );

    \I__4793\ : InMux
    port map (
            O => \N__28155\,
            I => \N__28144\
        );

    \I__4792\ : InMux
    port map (
            O => \N__28154\,
            I => \N__28144\
        );

    \I__4791\ : Span4Mux_v
    port map (
            O => \N__28151\,
            I => \N__28139\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__28144\,
            I => \N__28139\
        );

    \I__4789\ : Odrv4
    port map (
            O => \N__28139\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__4788\ : InMux
    port map (
            O => \N__28136\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__4787\ : InMux
    port map (
            O => \N__28133\,
            I => \N__28127\
        );

    \I__4786\ : InMux
    port map (
            O => \N__28132\,
            I => \N__28127\
        );

    \I__4785\ : LocalMux
    port map (
            O => \N__28127\,
            I => \N__28123\
        );

    \I__4784\ : InMux
    port map (
            O => \N__28126\,
            I => \N__28120\
        );

    \I__4783\ : Span4Mux_h
    port map (
            O => \N__28123\,
            I => \N__28117\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__28120\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__4781\ : Odrv4
    port map (
            O => \N__28117\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__4780\ : InMux
    port map (
            O => \N__28112\,
            I => \N__28108\
        );

    \I__4779\ : CascadeMux
    port map (
            O => \N__28111\,
            I => \N__28103\
        );

    \I__4778\ : LocalMux
    port map (
            O => \N__28108\,
            I => \N__28100\
        );

    \I__4777\ : InMux
    port map (
            O => \N__28107\,
            I => \N__28093\
        );

    \I__4776\ : InMux
    port map (
            O => \N__28106\,
            I => \N__28093\
        );

    \I__4775\ : InMux
    port map (
            O => \N__28103\,
            I => \N__28093\
        );

    \I__4774\ : Span4Mux_h
    port map (
            O => \N__28100\,
            I => \N__28088\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__28093\,
            I => \N__28088\
        );

    \I__4772\ : Odrv4
    port map (
            O => \N__28088\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__4771\ : InMux
    port map (
            O => \N__28085\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__4770\ : CascadeMux
    port map (
            O => \N__28082\,
            I => \N__28079\
        );

    \I__4769\ : InMux
    port map (
            O => \N__28079\,
            I => \N__28075\
        );

    \I__4768\ : InMux
    port map (
            O => \N__28078\,
            I => \N__28072\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__28075\,
            I => \N__28068\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__28072\,
            I => \N__28065\
        );

    \I__4765\ : InMux
    port map (
            O => \N__28071\,
            I => \N__28062\
        );

    \I__4764\ : Span4Mux_h
    port map (
            O => \N__28068\,
            I => \N__28059\
        );

    \I__4763\ : Span4Mux_h
    port map (
            O => \N__28065\,
            I => \N__28056\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__28062\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__4761\ : Odrv4
    port map (
            O => \N__28059\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__4760\ : Odrv4
    port map (
            O => \N__28056\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__4759\ : InMux
    port map (
            O => \N__28049\,
            I => \N__28046\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__28046\,
            I => \N__28040\
        );

    \I__4757\ : InMux
    port map (
            O => \N__28045\,
            I => \N__28035\
        );

    \I__4756\ : InMux
    port map (
            O => \N__28044\,
            I => \N__28035\
        );

    \I__4755\ : InMux
    port map (
            O => \N__28043\,
            I => \N__28032\
        );

    \I__4754\ : Span4Mux_h
    port map (
            O => \N__28040\,
            I => \N__28027\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__28035\,
            I => \N__28027\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__28032\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__4751\ : Odrv4
    port map (
            O => \N__28027\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__4750\ : InMux
    port map (
            O => \N__28022\,
            I => \bfn_10_13_0_\
        );

    \I__4749\ : CascadeMux
    port map (
            O => \N__28019\,
            I => \N__28015\
        );

    \I__4748\ : CascadeMux
    port map (
            O => \N__28018\,
            I => \N__28012\
        );

    \I__4747\ : InMux
    port map (
            O => \N__28015\,
            I => \N__28009\
        );

    \I__4746\ : InMux
    port map (
            O => \N__28012\,
            I => \N__28006\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__28009\,
            I => \N__28002\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__28006\,
            I => \N__27999\
        );

    \I__4743\ : InMux
    port map (
            O => \N__28005\,
            I => \N__27996\
        );

    \I__4742\ : Span4Mux_h
    port map (
            O => \N__28002\,
            I => \N__27993\
        );

    \I__4741\ : Span4Mux_h
    port map (
            O => \N__27999\,
            I => \N__27990\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__27996\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__4739\ : Odrv4
    port map (
            O => \N__27993\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__4738\ : Odrv4
    port map (
            O => \N__27990\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__4737\ : InMux
    port map (
            O => \N__27983\,
            I => \N__27977\
        );

    \I__4736\ : InMux
    port map (
            O => \N__27982\,
            I => \N__27974\
        );

    \I__4735\ : InMux
    port map (
            O => \N__27981\,
            I => \N__27971\
        );

    \I__4734\ : InMux
    port map (
            O => \N__27980\,
            I => \N__27968\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__27977\,
            I => \N__27961\
        );

    \I__4732\ : LocalMux
    port map (
            O => \N__27974\,
            I => \N__27961\
        );

    \I__4731\ : LocalMux
    port map (
            O => \N__27971\,
            I => \N__27961\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__27968\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__4729\ : Odrv4
    port map (
            O => \N__27961\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__4728\ : InMux
    port map (
            O => \N__27956\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__4727\ : InMux
    port map (
            O => \N__27953\,
            I => \N__27946\
        );

    \I__4726\ : InMux
    port map (
            O => \N__27952\,
            I => \N__27946\
        );

    \I__4725\ : InMux
    port map (
            O => \N__27951\,
            I => \N__27943\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__27946\,
            I => \N__27940\
        );

    \I__4723\ : LocalMux
    port map (
            O => \N__27943\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__4722\ : Odrv4
    port map (
            O => \N__27940\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__4721\ : InMux
    port map (
            O => \N__27935\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__4720\ : InMux
    port map (
            O => \N__27932\,
            I => \N__27926\
        );

    \I__4719\ : InMux
    port map (
            O => \N__27931\,
            I => \N__27926\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__27926\,
            I => \N__27922\
        );

    \I__4717\ : InMux
    port map (
            O => \N__27925\,
            I => \N__27919\
        );

    \I__4716\ : Span4Mux_h
    port map (
            O => \N__27922\,
            I => \N__27916\
        );

    \I__4715\ : LocalMux
    port map (
            O => \N__27919\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__4714\ : Odrv4
    port map (
            O => \N__27916\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__4713\ : InMux
    port map (
            O => \N__27911\,
            I => \N__27906\
        );

    \I__4712\ : InMux
    port map (
            O => \N__27910\,
            I => \N__27903\
        );

    \I__4711\ : InMux
    port map (
            O => \N__27909\,
            I => \N__27900\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__27906\,
            I => \N__27895\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__27903\,
            I => \N__27895\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__27900\,
            I => \N__27889\
        );

    \I__4707\ : Sp12to4
    port map (
            O => \N__27895\,
            I => \N__27889\
        );

    \I__4706\ : InMux
    port map (
            O => \N__27894\,
            I => \N__27886\
        );

    \I__4705\ : Odrv12
    port map (
            O => \N__27889\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__4704\ : LocalMux
    port map (
            O => \N__27886\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__4703\ : InMux
    port map (
            O => \N__27881\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__4702\ : CascadeMux
    port map (
            O => \N__27878\,
            I => \N__27874\
        );

    \I__4701\ : CascadeMux
    port map (
            O => \N__27877\,
            I => \N__27871\
        );

    \I__4700\ : InMux
    port map (
            O => \N__27874\,
            I => \N__27865\
        );

    \I__4699\ : InMux
    port map (
            O => \N__27871\,
            I => \N__27865\
        );

    \I__4698\ : InMux
    port map (
            O => \N__27870\,
            I => \N__27862\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__27865\,
            I => \N__27859\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__27862\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__4695\ : Odrv4
    port map (
            O => \N__27859\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__4694\ : InMux
    port map (
            O => \N__27854\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__4693\ : InMux
    port map (
            O => \N__27851\,
            I => \N__27845\
        );

    \I__4692\ : InMux
    port map (
            O => \N__27850\,
            I => \N__27845\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__27845\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_28\
        );

    \I__4690\ : CascadeMux
    port map (
            O => \N__27842\,
            I => \N__27839\
        );

    \I__4689\ : InMux
    port map (
            O => \N__27839\,
            I => \N__27836\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__27836\,
            I => \N__27833\
        );

    \I__4687\ : Odrv4
    port map (
            O => \N__27833\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt28\
        );

    \I__4686\ : CascadeMux
    port map (
            O => \N__27830\,
            I => \N__27827\
        );

    \I__4685\ : InMux
    port map (
            O => \N__27827\,
            I => \N__27821\
        );

    \I__4684\ : InMux
    port map (
            O => \N__27826\,
            I => \N__27821\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__27821\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_29\
        );

    \I__4682\ : InMux
    port map (
            O => \N__27818\,
            I => \N__27814\
        );

    \I__4681\ : InMux
    port map (
            O => \N__27817\,
            I => \N__27811\
        );

    \I__4680\ : LocalMux
    port map (
            O => \N__27814\,
            I => \N__27807\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__27811\,
            I => \N__27804\
        );

    \I__4678\ : InMux
    port map (
            O => \N__27810\,
            I => \N__27801\
        );

    \I__4677\ : Span4Mux_v
    port map (
            O => \N__27807\,
            I => \N__27796\
        );

    \I__4676\ : Span4Mux_v
    port map (
            O => \N__27804\,
            I => \N__27796\
        );

    \I__4675\ : LocalMux
    port map (
            O => \N__27801\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__4674\ : Odrv4
    port map (
            O => \N__27796\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__4673\ : InMux
    port map (
            O => \N__27791\,
            I => \N__27786\
        );

    \I__4672\ : InMux
    port map (
            O => \N__27790\,
            I => \N__27783\
        );

    \I__4671\ : InMux
    port map (
            O => \N__27789\,
            I => \N__27780\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__27786\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__27783\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__27780\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30\
        );

    \I__4667\ : InMux
    port map (
            O => \N__27773\,
            I => \N__27769\
        );

    \I__4666\ : InMux
    port map (
            O => \N__27772\,
            I => \N__27765\
        );

    \I__4665\ : LocalMux
    port map (
            O => \N__27769\,
            I => \N__27762\
        );

    \I__4664\ : InMux
    port map (
            O => \N__27768\,
            I => \N__27759\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__27765\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__4662\ : Odrv4
    port map (
            O => \N__27762\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__27759\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__4660\ : InMux
    port map (
            O => \N__27752\,
            I => \N__27747\
        );

    \I__4659\ : InMux
    port map (
            O => \N__27751\,
            I => \N__27744\
        );

    \I__4658\ : InMux
    port map (
            O => \N__27750\,
            I => \N__27741\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__27747\,
            I => \N__27736\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__27744\,
            I => \N__27736\
        );

    \I__4655\ : LocalMux
    port map (
            O => \N__27741\,
            I => \N__27732\
        );

    \I__4654\ : Span4Mux_v
    port map (
            O => \N__27736\,
            I => \N__27729\
        );

    \I__4653\ : InMux
    port map (
            O => \N__27735\,
            I => \N__27726\
        );

    \I__4652\ : Span4Mux_v
    port map (
            O => \N__27732\,
            I => \N__27723\
        );

    \I__4651\ : Span4Mux_h
    port map (
            O => \N__27729\,
            I => \N__27720\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__27726\,
            I => \N__27717\
        );

    \I__4649\ : Odrv4
    port map (
            O => \N__27723\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__4648\ : Odrv4
    port map (
            O => \N__27720\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__4647\ : Odrv12
    port map (
            O => \N__27717\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__4646\ : CascadeMux
    port map (
            O => \N__27710\,
            I => \N__27707\
        );

    \I__4645\ : InMux
    port map (
            O => \N__27707\,
            I => \N__27704\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__27704\,
            I => \N__27699\
        );

    \I__4643\ : InMux
    port map (
            O => \N__27703\,
            I => \N__27696\
        );

    \I__4642\ : InMux
    port map (
            O => \N__27702\,
            I => \N__27693\
        );

    \I__4641\ : Span4Mux_h
    port map (
            O => \N__27699\,
            I => \N__27690\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__27696\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__27693\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__4638\ : Odrv4
    port map (
            O => \N__27690\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__4637\ : InMux
    port map (
            O => \N__27683\,
            I => \N__27678\
        );

    \I__4636\ : InMux
    port map (
            O => \N__27682\,
            I => \N__27674\
        );

    \I__4635\ : InMux
    port map (
            O => \N__27681\,
            I => \N__27671\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__27678\,
            I => \N__27668\
        );

    \I__4633\ : CascadeMux
    port map (
            O => \N__27677\,
            I => \N__27665\
        );

    \I__4632\ : LocalMux
    port map (
            O => \N__27674\,
            I => \N__27662\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__27671\,
            I => \N__27659\
        );

    \I__4630\ : Span4Mux_v
    port map (
            O => \N__27668\,
            I => \N__27656\
        );

    \I__4629\ : InMux
    port map (
            O => \N__27665\,
            I => \N__27653\
        );

    \I__4628\ : Span4Mux_h
    port map (
            O => \N__27662\,
            I => \N__27648\
        );

    \I__4627\ : Span4Mux_v
    port map (
            O => \N__27659\,
            I => \N__27648\
        );

    \I__4626\ : Span4Mux_h
    port map (
            O => \N__27656\,
            I => \N__27645\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__27653\,
            I => \N__27642\
        );

    \I__4624\ : Odrv4
    port map (
            O => \N__27648\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__4623\ : Odrv4
    port map (
            O => \N__27645\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__4622\ : Odrv12
    port map (
            O => \N__27642\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__4621\ : InMux
    port map (
            O => \N__27635\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__4620\ : CascadeMux
    port map (
            O => \N__27632\,
            I => \N__27628\
        );

    \I__4619\ : InMux
    port map (
            O => \N__27631\,
            I => \N__27624\
        );

    \I__4618\ : InMux
    port map (
            O => \N__27628\,
            I => \N__27621\
        );

    \I__4617\ : InMux
    port map (
            O => \N__27627\,
            I => \N__27618\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__27624\,
            I => \N__27613\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__27621\,
            I => \N__27613\
        );

    \I__4614\ : LocalMux
    port map (
            O => \N__27618\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__4613\ : Odrv4
    port map (
            O => \N__27613\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__4612\ : InMux
    port map (
            O => \N__27608\,
            I => \N__27601\
        );

    \I__4611\ : InMux
    port map (
            O => \N__27607\,
            I => \N__27601\
        );

    \I__4610\ : InMux
    port map (
            O => \N__27606\,
            I => \N__27598\
        );

    \I__4609\ : LocalMux
    port map (
            O => \N__27601\,
            I => \N__27594\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__27598\,
            I => \N__27591\
        );

    \I__4607\ : InMux
    port map (
            O => \N__27597\,
            I => \N__27588\
        );

    \I__4606\ : Span4Mux_h
    port map (
            O => \N__27594\,
            I => \N__27585\
        );

    \I__4605\ : Span4Mux_v
    port map (
            O => \N__27591\,
            I => \N__27580\
        );

    \I__4604\ : LocalMux
    port map (
            O => \N__27588\,
            I => \N__27580\
        );

    \I__4603\ : Odrv4
    port map (
            O => \N__27585\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__4602\ : Odrv4
    port map (
            O => \N__27580\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__4601\ : InMux
    port map (
            O => \N__27575\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__4600\ : InMux
    port map (
            O => \N__27572\,
            I => \N__27565\
        );

    \I__4599\ : InMux
    port map (
            O => \N__27571\,
            I => \N__27565\
        );

    \I__4598\ : InMux
    port map (
            O => \N__27570\,
            I => \N__27562\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__27565\,
            I => \N__27559\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__27562\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__4595\ : Odrv4
    port map (
            O => \N__27559\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__4594\ : InMux
    port map (
            O => \N__27554\,
            I => \N__27551\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__27551\,
            I => \N__27545\
        );

    \I__4592\ : InMux
    port map (
            O => \N__27550\,
            I => \N__27542\
        );

    \I__4591\ : InMux
    port map (
            O => \N__27549\,
            I => \N__27539\
        );

    \I__4590\ : InMux
    port map (
            O => \N__27548\,
            I => \N__27536\
        );

    \I__4589\ : Span4Mux_v
    port map (
            O => \N__27545\,
            I => \N__27531\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__27542\,
            I => \N__27531\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__27539\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__27536\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__4585\ : Odrv4
    port map (
            O => \N__27531\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__4584\ : InMux
    port map (
            O => \N__27524\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__4583\ : CascadeMux
    port map (
            O => \N__27521\,
            I => \N__27517\
        );

    \I__4582\ : CascadeMux
    port map (
            O => \N__27520\,
            I => \N__27514\
        );

    \I__4581\ : InMux
    port map (
            O => \N__27517\,
            I => \N__27508\
        );

    \I__4580\ : InMux
    port map (
            O => \N__27514\,
            I => \N__27508\
        );

    \I__4579\ : InMux
    port map (
            O => \N__27513\,
            I => \N__27505\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__27508\,
            I => \N__27502\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__27505\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__4576\ : Odrv4
    port map (
            O => \N__27502\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__4575\ : InMux
    port map (
            O => \N__27497\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__4574\ : InMux
    port map (
            O => \N__27494\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_30\
        );

    \I__4573\ : CascadeMux
    port map (
            O => \N__27491\,
            I => \N__27488\
        );

    \I__4572\ : InMux
    port map (
            O => \N__27488\,
            I => \N__27485\
        );

    \I__4571\ : LocalMux
    port map (
            O => \N__27485\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt24\
        );

    \I__4570\ : InMux
    port map (
            O => \N__27482\,
            I => \N__27476\
        );

    \I__4569\ : InMux
    port map (
            O => \N__27481\,
            I => \N__27476\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__27476\,
            I => \N__27473\
        );

    \I__4567\ : Odrv12
    port map (
            O => \N__27473\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_24\
        );

    \I__4566\ : CascadeMux
    port map (
            O => \N__27470\,
            I => \N__27466\
        );

    \I__4565\ : InMux
    port map (
            O => \N__27469\,
            I => \N__27461\
        );

    \I__4564\ : InMux
    port map (
            O => \N__27466\,
            I => \N__27461\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__27461\,
            I => \N__27458\
        );

    \I__4562\ : Odrv12
    port map (
            O => \N__27458\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_25\
        );

    \I__4561\ : InMux
    port map (
            O => \N__27455\,
            I => \N__27452\
        );

    \I__4560\ : LocalMux
    port map (
            O => \N__27452\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24\
        );

    \I__4559\ : InMux
    port map (
            O => \N__27449\,
            I => \N__27446\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__27446\,
            I => \N__27442\
        );

    \I__4557\ : InMux
    port map (
            O => \N__27445\,
            I => \N__27438\
        );

    \I__4556\ : Span4Mux_h
    port map (
            O => \N__27442\,
            I => \N__27435\
        );

    \I__4555\ : InMux
    port map (
            O => \N__27441\,
            I => \N__27432\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__27438\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12\
        );

    \I__4553\ : Odrv4
    port map (
            O => \N__27435\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__27432\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12\
        );

    \I__4551\ : InMux
    port map (
            O => \N__27425\,
            I => \N__27422\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__27422\,
            I => \N__27419\
        );

    \I__4549\ : Odrv4
    port map (
            O => \N__27419\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\
        );

    \I__4548\ : InMux
    port map (
            O => \N__27416\,
            I => \N__27413\
        );

    \I__4547\ : LocalMux
    port map (
            O => \N__27413\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26\
        );

    \I__4546\ : CascadeMux
    port map (
            O => \N__27410\,
            I => \N__27407\
        );

    \I__4545\ : InMux
    port map (
            O => \N__27407\,
            I => \N__27404\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__27404\,
            I => \N__27401\
        );

    \I__4543\ : Odrv4
    port map (
            O => \N__27401\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt26\
        );

    \I__4542\ : InMux
    port map (
            O => \N__27398\,
            I => \N__27395\
        );

    \I__4541\ : LocalMux
    port map (
            O => \N__27395\,
            I => \N__27392\
        );

    \I__4540\ : Span4Mux_h
    port map (
            O => \N__27392\,
            I => \N__27388\
        );

    \I__4539\ : InMux
    port map (
            O => \N__27391\,
            I => \N__27385\
        );

    \I__4538\ : Odrv4
    port map (
            O => \N__27388\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__27385\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27\
        );

    \I__4536\ : InMux
    port map (
            O => \N__27380\,
            I => \N__27376\
        );

    \I__4535\ : InMux
    port map (
            O => \N__27379\,
            I => \N__27373\
        );

    \I__4534\ : LocalMux
    port map (
            O => \N__27376\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__27373\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\
        );

    \I__4532\ : InMux
    port map (
            O => \N__27368\,
            I => \N__27365\
        );

    \I__4531\ : LocalMux
    port map (
            O => \N__27365\,
            I => \N__27362\
        );

    \I__4530\ : Odrv4
    port map (
            O => \N__27362\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28\
        );

    \I__4529\ : InMux
    port map (
            O => \N__27359\,
            I => \N__27356\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__27356\,
            I => \N__27353\
        );

    \I__4527\ : Odrv4
    port map (
            O => \N__27353\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\
        );

    \I__4526\ : CascadeMux
    port map (
            O => \N__27350\,
            I => \N__27347\
        );

    \I__4525\ : InMux
    port map (
            O => \N__27347\,
            I => \N__27344\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__27344\,
            I => \N__27341\
        );

    \I__4523\ : Span4Mux_h
    port map (
            O => \N__27341\,
            I => \N__27338\
        );

    \I__4522\ : Odrv4
    port map (
            O => \N__27338\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt18\
        );

    \I__4521\ : InMux
    port map (
            O => \N__27335\,
            I => \N__27332\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__27332\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22\
        );

    \I__4519\ : CascadeMux
    port map (
            O => \N__27329\,
            I => \N__27326\
        );

    \I__4518\ : InMux
    port map (
            O => \N__27326\,
            I => \N__27323\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__27323\,
            I => \N__27320\
        );

    \I__4516\ : Odrv4
    port map (
            O => \N__27320\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt22\
        );

    \I__4515\ : InMux
    port map (
            O => \N__27317\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_28\
        );

    \I__4514\ : InMux
    port map (
            O => \N__27314\,
            I => \N__27311\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__27311\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\
        );

    \I__4512\ : InMux
    port map (
            O => \N__27308\,
            I => \N__27305\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__27305\,
            I => \N__27302\
        );

    \I__4510\ : Odrv4
    port map (
            O => \N__27302\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\
        );

    \I__4509\ : CascadeMux
    port map (
            O => \N__27299\,
            I => \N__27296\
        );

    \I__4508\ : InMux
    port map (
            O => \N__27296\,
            I => \N__27293\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__27293\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\
        );

    \I__4506\ : InMux
    port map (
            O => \N__27290\,
            I => \N__27287\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__27287\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\
        );

    \I__4504\ : CascadeMux
    port map (
            O => \N__27284\,
            I => \N__27281\
        );

    \I__4503\ : InMux
    port map (
            O => \N__27281\,
            I => \N__27278\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__27278\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\
        );

    \I__4501\ : CascadeMux
    port map (
            O => \N__27275\,
            I => \N__27272\
        );

    \I__4500\ : InMux
    port map (
            O => \N__27272\,
            I => \N__27269\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__27269\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\
        );

    \I__4498\ : InMux
    port map (
            O => \N__27266\,
            I => \N__27263\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__27263\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\
        );

    \I__4496\ : CascadeMux
    port map (
            O => \N__27260\,
            I => \N__27257\
        );

    \I__4495\ : InMux
    port map (
            O => \N__27257\,
            I => \N__27254\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__27254\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\
        );

    \I__4493\ : CascadeMux
    port map (
            O => \N__27251\,
            I => \N__27248\
        );

    \I__4492\ : InMux
    port map (
            O => \N__27248\,
            I => \N__27245\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__27245\,
            I => \N__27242\
        );

    \I__4490\ : Odrv4
    port map (
            O => \N__27242\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\
        );

    \I__4489\ : InMux
    port map (
            O => \N__27239\,
            I => \N__27236\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__27236\,
            I => \N__27233\
        );

    \I__4487\ : Odrv4
    port map (
            O => \N__27233\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\
        );

    \I__4486\ : CascadeMux
    port map (
            O => \N__27230\,
            I => \N__27227\
        );

    \I__4485\ : InMux
    port map (
            O => \N__27227\,
            I => \N__27224\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__27224\,
            I => \N__27221\
        );

    \I__4483\ : Odrv4
    port map (
            O => \N__27221\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\
        );

    \I__4482\ : CascadeMux
    port map (
            O => \N__27218\,
            I => \N__27215\
        );

    \I__4481\ : InMux
    port map (
            O => \N__27215\,
            I => \N__27212\
        );

    \I__4480\ : LocalMux
    port map (
            O => \N__27212\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\
        );

    \I__4479\ : InMux
    port map (
            O => \N__27209\,
            I => \N__27204\
        );

    \I__4478\ : InMux
    port map (
            O => \N__27208\,
            I => \N__27201\
        );

    \I__4477\ : InMux
    port map (
            O => \N__27207\,
            I => \N__27198\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__27204\,
            I => \N__27195\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__27201\,
            I => \N__27192\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__27198\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__4473\ : Odrv12
    port map (
            O => \N__27195\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__4472\ : Odrv4
    port map (
            O => \N__27192\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__4471\ : CascadeMux
    port map (
            O => \N__27185\,
            I => \N__27182\
        );

    \I__4470\ : InMux
    port map (
            O => \N__27182\,
            I => \N__27179\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__27179\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\
        );

    \I__4468\ : InMux
    port map (
            O => \N__27176\,
            I => \N__27173\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__27173\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\
        );

    \I__4466\ : InMux
    port map (
            O => \N__27170\,
            I => \N__27167\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__27167\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\
        );

    \I__4464\ : CascadeMux
    port map (
            O => \N__27164\,
            I => \N__27161\
        );

    \I__4463\ : InMux
    port map (
            O => \N__27161\,
            I => \N__27158\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__27158\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\
        );

    \I__4461\ : InMux
    port map (
            O => \N__27155\,
            I => \N__27152\
        );

    \I__4460\ : LocalMux
    port map (
            O => \N__27152\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\
        );

    \I__4459\ : CascadeMux
    port map (
            O => \N__27149\,
            I => \N__27146\
        );

    \I__4458\ : InMux
    port map (
            O => \N__27146\,
            I => \N__27143\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__27143\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\
        );

    \I__4456\ : InMux
    port map (
            O => \N__27140\,
            I => \N__27137\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__27137\,
            I => \N__27134\
        );

    \I__4454\ : Odrv4
    port map (
            O => \N__27134\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\
        );

    \I__4453\ : CascadeMux
    port map (
            O => \N__27131\,
            I => \N__27128\
        );

    \I__4452\ : InMux
    port map (
            O => \N__27128\,
            I => \N__27125\
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__27125\,
            I => \N__27122\
        );

    \I__4450\ : Odrv4
    port map (
            O => \N__27122\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\
        );

    \I__4449\ : InMux
    port map (
            O => \N__27119\,
            I => \N__27116\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__27116\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\
        );

    \I__4447\ : CascadeMux
    port map (
            O => \N__27113\,
            I => \N__27110\
        );

    \I__4446\ : InMux
    port map (
            O => \N__27110\,
            I => \N__27107\
        );

    \I__4445\ : LocalMux
    port map (
            O => \N__27107\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\
        );

    \I__4444\ : InMux
    port map (
            O => \N__27104\,
            I => \N__27101\
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__27101\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\
        );

    \I__4442\ : CascadeMux
    port map (
            O => \N__27098\,
            I => \N__27095\
        );

    \I__4441\ : InMux
    port map (
            O => \N__27095\,
            I => \N__27092\
        );

    \I__4440\ : LocalMux
    port map (
            O => \N__27092\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\
        );

    \I__4439\ : CascadeMux
    port map (
            O => \N__27089\,
            I => \N__27086\
        );

    \I__4438\ : InMux
    port map (
            O => \N__27086\,
            I => \N__27083\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__27083\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\
        );

    \I__4436\ : InMux
    port map (
            O => \N__27080\,
            I => \N__27076\
        );

    \I__4435\ : InMux
    port map (
            O => \N__27079\,
            I => \N__27072\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__27076\,
            I => \N__27069\
        );

    \I__4433\ : InMux
    port map (
            O => \N__27075\,
            I => \N__27066\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__27072\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19\
        );

    \I__4431\ : Odrv4
    port map (
            O => \N__27069\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__27066\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19\
        );

    \I__4429\ : CascadeMux
    port map (
            O => \N__27059\,
            I => \N__27055\
        );

    \I__4428\ : CascadeMux
    port map (
            O => \N__27058\,
            I => \N__27052\
        );

    \I__4427\ : InMux
    port map (
            O => \N__27055\,
            I => \N__27047\
        );

    \I__4426\ : InMux
    port map (
            O => \N__27052\,
            I => \N__27047\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__27047\,
            I => \N__27044\
        );

    \I__4424\ : Odrv4
    port map (
            O => \N__27044\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\
        );

    \I__4423\ : CascadeMux
    port map (
            O => \N__27041\,
            I => \N__27038\
        );

    \I__4422\ : InMux
    port map (
            O => \N__27038\,
            I => \N__27035\
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__27035\,
            I => \N__27032\
        );

    \I__4420\ : Span4Mux_v
    port map (
            O => \N__27032\,
            I => \N__27029\
        );

    \I__4419\ : Span4Mux_v
    port map (
            O => \N__27029\,
            I => \N__27026\
        );

    \I__4418\ : Odrv4
    port map (
            O => \N__27026\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\
        );

    \I__4417\ : InMux
    port map (
            O => \N__27023\,
            I => \N__27020\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__27020\,
            I => \N__27016\
        );

    \I__4415\ : InMux
    port map (
            O => \N__27019\,
            I => \N__27013\
        );

    \I__4414\ : Span4Mux_h
    port map (
            O => \N__27016\,
            I => \N__27010\
        );

    \I__4413\ : LocalMux
    port map (
            O => \N__27013\,
            I => \elapsed_time_ns_1_RNIL73T9_0_9\
        );

    \I__4412\ : Odrv4
    port map (
            O => \N__27010\,
            I => \elapsed_time_ns_1_RNIL73T9_0_9\
        );

    \I__4411\ : InMux
    port map (
            O => \N__27005\,
            I => \N__27001\
        );

    \I__4410\ : InMux
    port map (
            O => \N__27004\,
            I => \N__26998\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__27001\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__26998\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18\
        );

    \I__4407\ : InMux
    port map (
            O => \N__26993\,
            I => \N__26987\
        );

    \I__4406\ : InMux
    port map (
            O => \N__26992\,
            I => \N__26987\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__26987\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\
        );

    \I__4404\ : InMux
    port map (
            O => \N__26984\,
            I => \N__26981\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__26981\,
            I => \N__26977\
        );

    \I__4402\ : InMux
    port map (
            O => \N__26980\,
            I => \N__26973\
        );

    \I__4401\ : Span4Mux_h
    port map (
            O => \N__26977\,
            I => \N__26970\
        );

    \I__4400\ : InMux
    port map (
            O => \N__26976\,
            I => \N__26967\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__26973\,
            I => \elapsed_time_ns_1_RNIDV2T9_0_1\
        );

    \I__4398\ : Odrv4
    port map (
            O => \N__26970\,
            I => \elapsed_time_ns_1_RNIDV2T9_0_1\
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__26967\,
            I => \elapsed_time_ns_1_RNIDV2T9_0_1\
        );

    \I__4396\ : InMux
    port map (
            O => \N__26960\,
            I => \N__26955\
        );

    \I__4395\ : InMux
    port map (
            O => \N__26959\,
            I => \N__26952\
        );

    \I__4394\ : InMux
    port map (
            O => \N__26958\,
            I => \N__26949\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__26955\,
            I => \N__26946\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__26952\,
            I => \N__26942\
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__26949\,
            I => \N__26937\
        );

    \I__4390\ : Span4Mux_h
    port map (
            O => \N__26946\,
            I => \N__26937\
        );

    \I__4389\ : InMux
    port map (
            O => \N__26945\,
            I => \N__26934\
        );

    \I__4388\ : Span12Mux_v
    port map (
            O => \N__26942\,
            I => \N__26931\
        );

    \I__4387\ : Span4Mux_v
    port map (
            O => \N__26937\,
            I => \N__26926\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__26934\,
            I => \N__26926\
        );

    \I__4385\ : Odrv12
    port map (
            O => \N__26931\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__4384\ : Odrv4
    port map (
            O => \N__26926\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__4383\ : InMux
    port map (
            O => \N__26921\,
            I => \N__26918\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__26918\,
            I => \N__26914\
        );

    \I__4381\ : InMux
    port map (
            O => \N__26917\,
            I => \N__26910\
        );

    \I__4380\ : Span4Mux_v
    port map (
            O => \N__26914\,
            I => \N__26907\
        );

    \I__4379\ : InMux
    port map (
            O => \N__26913\,
            I => \N__26904\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__26910\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24\
        );

    \I__4377\ : Odrv4
    port map (
            O => \N__26907\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__26904\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24\
        );

    \I__4375\ : InMux
    port map (
            O => \N__26897\,
            I => \N__26892\
        );

    \I__4374\ : InMux
    port map (
            O => \N__26896\,
            I => \N__26889\
        );

    \I__4373\ : InMux
    port map (
            O => \N__26895\,
            I => \N__26886\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__26892\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__26889\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17\
        );

    \I__4370\ : LocalMux
    port map (
            O => \N__26886\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17\
        );

    \I__4369\ : InMux
    port map (
            O => \N__26879\,
            I => \N__26876\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__26876\,
            I => \N__26873\
        );

    \I__4367\ : Span4Mux_h
    port map (
            O => \N__26873\,
            I => \N__26868\
        );

    \I__4366\ : InMux
    port map (
            O => \N__26872\,
            I => \N__26865\
        );

    \I__4365\ : InMux
    port map (
            O => \N__26871\,
            I => \N__26862\
        );

    \I__4364\ : Span4Mux_v
    port map (
            O => \N__26868\,
            I => \N__26859\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__26865\,
            I => \elapsed_time_ns_1_RNII43T9_0_6\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__26862\,
            I => \elapsed_time_ns_1_RNII43T9_0_6\
        );

    \I__4361\ : Odrv4
    port map (
            O => \N__26859\,
            I => \elapsed_time_ns_1_RNII43T9_0_6\
        );

    \I__4360\ : InMux
    port map (
            O => \N__26852\,
            I => \N__26848\
        );

    \I__4359\ : InMux
    port map (
            O => \N__26851\,
            I => \N__26844\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__26848\,
            I => \N__26841\
        );

    \I__4357\ : InMux
    port map (
            O => \N__26847\,
            I => \N__26838\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__26844\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14\
        );

    \I__4355\ : Odrv4
    port map (
            O => \N__26841\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__26838\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14\
        );

    \I__4353\ : InMux
    port map (
            O => \N__26831\,
            I => \N__26828\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__26828\,
            I => \pwm_generator_inst.counter_i_4\
        );

    \I__4351\ : CascadeMux
    port map (
            O => \N__26825\,
            I => \N__26822\
        );

    \I__4350\ : InMux
    port map (
            O => \N__26822\,
            I => \N__26819\
        );

    \I__4349\ : LocalMux
    port map (
            O => \N__26819\,
            I => \N__26816\
        );

    \I__4348\ : Odrv4
    port map (
            O => \N__26816\,
            I => \pwm_generator_inst.threshold_5\
        );

    \I__4347\ : InMux
    port map (
            O => \N__26813\,
            I => \N__26810\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__26810\,
            I => \pwm_generator_inst.counter_i_5\
        );

    \I__4345\ : CascadeMux
    port map (
            O => \N__26807\,
            I => \N__26804\
        );

    \I__4344\ : InMux
    port map (
            O => \N__26804\,
            I => \N__26801\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__26801\,
            I => \N__26798\
        );

    \I__4342\ : Span4Mux_h
    port map (
            O => \N__26798\,
            I => \N__26795\
        );

    \I__4341\ : Odrv4
    port map (
            O => \N__26795\,
            I => \pwm_generator_inst.un14_counter_6\
        );

    \I__4340\ : InMux
    port map (
            O => \N__26792\,
            I => \N__26789\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__26789\,
            I => \pwm_generator_inst.counter_i_6\
        );

    \I__4338\ : CascadeMux
    port map (
            O => \N__26786\,
            I => \N__26783\
        );

    \I__4337\ : InMux
    port map (
            O => \N__26783\,
            I => \N__26780\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__26780\,
            I => \pwm_generator_inst.un14_counter_7\
        );

    \I__4335\ : InMux
    port map (
            O => \N__26777\,
            I => \N__26774\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__26774\,
            I => \pwm_generator_inst.counter_i_7\
        );

    \I__4333\ : CascadeMux
    port map (
            O => \N__26771\,
            I => \N__26768\
        );

    \I__4332\ : InMux
    port map (
            O => \N__26768\,
            I => \N__26765\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__26765\,
            I => \N__26762\
        );

    \I__4330\ : Odrv4
    port map (
            O => \N__26762\,
            I => \pwm_generator_inst.un14_counter_8\
        );

    \I__4329\ : InMux
    port map (
            O => \N__26759\,
            I => \N__26756\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__26756\,
            I => \pwm_generator_inst.counter_i_8\
        );

    \I__4327\ : CascadeMux
    port map (
            O => \N__26753\,
            I => \N__26750\
        );

    \I__4326\ : InMux
    port map (
            O => \N__26750\,
            I => \N__26747\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__26747\,
            I => \pwm_generator_inst.threshold_9\
        );

    \I__4324\ : InMux
    port map (
            O => \N__26744\,
            I => \N__26741\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__26741\,
            I => \pwm_generator_inst.counter_i_9\
        );

    \I__4322\ : InMux
    port map (
            O => \N__26738\,
            I => \pwm_generator_inst.un14_counter_cry_9\
        );

    \I__4321\ : IoInMux
    port map (
            O => \N__26735\,
            I => \N__26732\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__26732\,
            I => \N__26729\
        );

    \I__4319\ : Span4Mux_s2_v
    port map (
            O => \N__26729\,
            I => \N__26726\
        );

    \I__4318\ : Sp12to4
    port map (
            O => \N__26726\,
            I => \N__26723\
        );

    \I__4317\ : Span12Mux_h
    port map (
            O => \N__26723\,
            I => \N__26720\
        );

    \I__4316\ : Span12Mux_v
    port map (
            O => \N__26720\,
            I => \N__26717\
        );

    \I__4315\ : Odrv12
    port map (
            O => \N__26717\,
            I => pwm_output_c
        );

    \I__4314\ : IoInMux
    port map (
            O => \N__26714\,
            I => \N__26711\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__26711\,
            I => s3_phy_c
        );

    \I__4312\ : InMux
    port map (
            O => \N__26708\,
            I => \N__26705\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__26705\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\
        );

    \I__4310\ : InMux
    port map (
            O => \N__26702\,
            I => \current_shift_inst.control_input_cry_10\
        );

    \I__4309\ : InMux
    port map (
            O => \N__26699\,
            I => \N__26696\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__26696\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\
        );

    \I__4307\ : InMux
    port map (
            O => \N__26693\,
            I => \current_shift_inst.control_input_cry_11\
        );

    \I__4306\ : InMux
    port map (
            O => \N__26690\,
            I => \current_shift_inst.control_input_cry_12\
        );

    \I__4305\ : InMux
    port map (
            O => \N__26687\,
            I => \N__26683\
        );

    \I__4304\ : InMux
    port map (
            O => \N__26686\,
            I => \N__26680\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__26683\,
            I => \current_shift_inst.control_input_31\
        );

    \I__4302\ : LocalMux
    port map (
            O => \N__26680\,
            I => \current_shift_inst.control_input_31\
        );

    \I__4301\ : InMux
    port map (
            O => \N__26675\,
            I => \N__26672\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__26672\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\
        );

    \I__4299\ : CascadeMux
    port map (
            O => \N__26669\,
            I => \N__26666\
        );

    \I__4298\ : InMux
    port map (
            O => \N__26666\,
            I => \N__26663\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__26663\,
            I => \N__26660\
        );

    \I__4296\ : Odrv4
    port map (
            O => \N__26660\,
            I => \pwm_generator_inst.threshold_0\
        );

    \I__4295\ : InMux
    port map (
            O => \N__26657\,
            I => \N__26654\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__26654\,
            I => \pwm_generator_inst.counter_i_0\
        );

    \I__4293\ : CascadeMux
    port map (
            O => \N__26651\,
            I => \N__26648\
        );

    \I__4292\ : InMux
    port map (
            O => \N__26648\,
            I => \N__26645\
        );

    \I__4291\ : LocalMux
    port map (
            O => \N__26645\,
            I => \pwm_generator_inst.un14_counter_1\
        );

    \I__4290\ : InMux
    port map (
            O => \N__26642\,
            I => \N__26639\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__26639\,
            I => \pwm_generator_inst.counter_i_1\
        );

    \I__4288\ : CascadeMux
    port map (
            O => \N__26636\,
            I => \N__26633\
        );

    \I__4287\ : InMux
    port map (
            O => \N__26633\,
            I => \N__26630\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__26630\,
            I => \pwm_generator_inst.threshold_2\
        );

    \I__4285\ : InMux
    port map (
            O => \N__26627\,
            I => \N__26624\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__26624\,
            I => \pwm_generator_inst.counter_i_2\
        );

    \I__4283\ : CascadeMux
    port map (
            O => \N__26621\,
            I => \N__26618\
        );

    \I__4282\ : InMux
    port map (
            O => \N__26618\,
            I => \N__26615\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__26615\,
            I => \pwm_generator_inst.threshold_3\
        );

    \I__4280\ : InMux
    port map (
            O => \N__26612\,
            I => \N__26609\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__26609\,
            I => \pwm_generator_inst.counter_i_3\
        );

    \I__4278\ : CascadeMux
    port map (
            O => \N__26606\,
            I => \N__26603\
        );

    \I__4277\ : InMux
    port map (
            O => \N__26603\,
            I => \N__26600\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__26600\,
            I => \N__26597\
        );

    \I__4275\ : Odrv4
    port map (
            O => \N__26597\,
            I => \pwm_generator_inst.threshold_4\
        );

    \I__4274\ : InMux
    port map (
            O => \N__26594\,
            I => \N__26591\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__26591\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\
        );

    \I__4272\ : InMux
    port map (
            O => \N__26588\,
            I => \current_shift_inst.control_input_cry_2\
        );

    \I__4271\ : InMux
    port map (
            O => \N__26585\,
            I => \N__26582\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__26582\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\
        );

    \I__4269\ : InMux
    port map (
            O => \N__26579\,
            I => \current_shift_inst.control_input_cry_3\
        );

    \I__4268\ : InMux
    port map (
            O => \N__26576\,
            I => \N__26573\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__26573\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\
        );

    \I__4266\ : InMux
    port map (
            O => \N__26570\,
            I => \current_shift_inst.control_input_cry_4\
        );

    \I__4265\ : InMux
    port map (
            O => \N__26567\,
            I => \N__26564\
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__26564\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\
        );

    \I__4263\ : InMux
    port map (
            O => \N__26561\,
            I => \current_shift_inst.control_input_cry_5\
        );

    \I__4262\ : InMux
    port map (
            O => \N__26558\,
            I => \N__26555\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__26555\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\
        );

    \I__4260\ : InMux
    port map (
            O => \N__26552\,
            I => \current_shift_inst.control_input_cry_6\
        );

    \I__4259\ : InMux
    port map (
            O => \N__26549\,
            I => \N__26546\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__26546\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\
        );

    \I__4257\ : InMux
    port map (
            O => \N__26543\,
            I => \bfn_9_20_0_\
        );

    \I__4256\ : InMux
    port map (
            O => \N__26540\,
            I => \N__26537\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__26537\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\
        );

    \I__4254\ : InMux
    port map (
            O => \N__26534\,
            I => \current_shift_inst.control_input_cry_8\
        );

    \I__4253\ : InMux
    port map (
            O => \N__26531\,
            I => \N__26528\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__26528\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\
        );

    \I__4251\ : InMux
    port map (
            O => \N__26525\,
            I => \current_shift_inst.control_input_cry_9\
        );

    \I__4250\ : InMux
    port map (
            O => \N__26522\,
            I => \bfn_9_18_0_\
        );

    \I__4249\ : InMux
    port map (
            O => \N__26519\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_24\
        );

    \I__4248\ : InMux
    port map (
            O => \N__26516\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_25\
        );

    \I__4247\ : InMux
    port map (
            O => \N__26513\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_26\
        );

    \I__4246\ : InMux
    port map (
            O => \N__26510\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_27\
        );

    \I__4245\ : InMux
    port map (
            O => \N__26507\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_28\
        );

    \I__4244\ : InMux
    port map (
            O => \N__26504\,
            I => \N__26501\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__26501\,
            I => \current_shift_inst.control_input_18\
        );

    \I__4242\ : InMux
    port map (
            O => \N__26498\,
            I => \N__26495\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__26495\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\
        );

    \I__4240\ : InMux
    port map (
            O => \N__26492\,
            I => \current_shift_inst.control_input_cry_0\
        );

    \I__4239\ : InMux
    port map (
            O => \N__26489\,
            I => \N__26486\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__26486\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\
        );

    \I__4237\ : InMux
    port map (
            O => \N__26483\,
            I => \current_shift_inst.control_input_cry_1\
        );

    \I__4236\ : InMux
    port map (
            O => \N__26480\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_14\
        );

    \I__4235\ : InMux
    port map (
            O => \N__26477\,
            I => \bfn_9_17_0_\
        );

    \I__4234\ : InMux
    port map (
            O => \N__26474\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_16\
        );

    \I__4233\ : InMux
    port map (
            O => \N__26471\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_17\
        );

    \I__4232\ : InMux
    port map (
            O => \N__26468\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_18\
        );

    \I__4231\ : InMux
    port map (
            O => \N__26465\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_19\
        );

    \I__4230\ : InMux
    port map (
            O => \N__26462\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_20\
        );

    \I__4229\ : InMux
    port map (
            O => \N__26459\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_21\
        );

    \I__4228\ : InMux
    port map (
            O => \N__26456\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_22\
        );

    \I__4227\ : InMux
    port map (
            O => \N__26453\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_5\
        );

    \I__4226\ : InMux
    port map (
            O => \N__26450\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_6\
        );

    \I__4225\ : InMux
    port map (
            O => \N__26447\,
            I => \bfn_9_16_0_\
        );

    \I__4224\ : InMux
    port map (
            O => \N__26444\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_8\
        );

    \I__4223\ : InMux
    port map (
            O => \N__26441\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_9\
        );

    \I__4222\ : InMux
    port map (
            O => \N__26438\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_10\
        );

    \I__4221\ : InMux
    port map (
            O => \N__26435\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_11\
        );

    \I__4220\ : InMux
    port map (
            O => \N__26432\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_12\
        );

    \I__4219\ : InMux
    port map (
            O => \N__26429\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_13\
        );

    \I__4218\ : InMux
    port map (
            O => \N__26426\,
            I => \N__26423\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__26423\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20\
        );

    \I__4216\ : InMux
    port map (
            O => \N__26420\,
            I => \N__26417\
        );

    \I__4215\ : LocalMux
    port map (
            O => \N__26417\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\
        );

    \I__4214\ : InMux
    port map (
            O => \N__26414\,
            I => \bfn_9_15_0_\
        );

    \I__4213\ : InMux
    port map (
            O => \N__26411\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_0\
        );

    \I__4212\ : InMux
    port map (
            O => \N__26408\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_1\
        );

    \I__4211\ : InMux
    port map (
            O => \N__26405\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_2\
        );

    \I__4210\ : InMux
    port map (
            O => \N__26402\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_3\
        );

    \I__4209\ : InMux
    port map (
            O => \N__26399\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_4\
        );

    \I__4208\ : InMux
    port map (
            O => \N__26396\,
            I => \N__26393\
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__26393\,
            I => \N__26390\
        );

    \I__4206\ : Odrv4
    port map (
            O => \N__26390\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15\
        );

    \I__4205\ : InMux
    port map (
            O => \N__26387\,
            I => \N__26384\
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__26384\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\
        );

    \I__4203\ : CascadeMux
    port map (
            O => \N__26381\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18_cascade_\
        );

    \I__4202\ : InMux
    port map (
            O => \N__26378\,
            I => \N__26375\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__26375\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19\
        );

    \I__4200\ : CascadeMux
    port map (
            O => \N__26372\,
            I => \N__26369\
        );

    \I__4199\ : InMux
    port map (
            O => \N__26369\,
            I => \N__26366\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__26366\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\
        );

    \I__4197\ : InMux
    port map (
            O => \N__26363\,
            I => \N__26360\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__26360\,
            I => \N__26355\
        );

    \I__4195\ : InMux
    port map (
            O => \N__26359\,
            I => \N__26352\
        );

    \I__4194\ : InMux
    port map (
            O => \N__26358\,
            I => \N__26349\
        );

    \I__4193\ : Span4Mux_h
    port map (
            O => \N__26355\,
            I => \N__26344\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__26352\,
            I => \N__26344\
        );

    \I__4191\ : LocalMux
    port map (
            O => \N__26349\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11\
        );

    \I__4190\ : Odrv4
    port map (
            O => \N__26344\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11\
        );

    \I__4189\ : InMux
    port map (
            O => \N__26339\,
            I => \N__26336\
        );

    \I__4188\ : LocalMux
    port map (
            O => \N__26336\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\
        );

    \I__4187\ : InMux
    port map (
            O => \N__26333\,
            I => \N__26324\
        );

    \I__4186\ : InMux
    port map (
            O => \N__26332\,
            I => \N__26324\
        );

    \I__4185\ : InMux
    port map (
            O => \N__26331\,
            I => \N__26324\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__26324\,
            I => \N__26321\
        );

    \I__4183\ : Span4Mux_h
    port map (
            O => \N__26321\,
            I => \N__26318\
        );

    \I__4182\ : Odrv4
    port map (
            O => \N__26318\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_30\
        );

    \I__4181\ : InMux
    port map (
            O => \N__26315\,
            I => \N__26312\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__26312\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\
        );

    \I__4179\ : InMux
    port map (
            O => \N__26309\,
            I => \N__26303\
        );

    \I__4178\ : InMux
    port map (
            O => \N__26308\,
            I => \N__26303\
        );

    \I__4177\ : LocalMux
    port map (
            O => \N__26303\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_26\
        );

    \I__4176\ : CascadeMux
    port map (
            O => \N__26300\,
            I => \N__26297\
        );

    \I__4175\ : InMux
    port map (
            O => \N__26297\,
            I => \N__26294\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__26294\,
            I => \N__26291\
        );

    \I__4173\ : Span4Mux_v
    port map (
            O => \N__26291\,
            I => \N__26288\
        );

    \I__4172\ : Odrv4
    port map (
            O => \N__26288\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\
        );

    \I__4171\ : InMux
    port map (
            O => \N__26285\,
            I => \N__26282\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__26282\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\
        );

    \I__4169\ : InMux
    port map (
            O => \N__26279\,
            I => \N__26276\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__26276\,
            I => \N__26273\
        );

    \I__4167\ : Odrv4
    port map (
            O => \N__26273\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\
        );

    \I__4166\ : CascadeMux
    port map (
            O => \N__26270\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\
        );

    \I__4165\ : CascadeMux
    port map (
            O => \N__26267\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_\
        );

    \I__4164\ : InMux
    port map (
            O => \N__26264\,
            I => \N__26260\
        );

    \I__4163\ : InMux
    port map (
            O => \N__26263\,
            I => \N__26257\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__26260\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10\
        );

    \I__4161\ : LocalMux
    port map (
            O => \N__26257\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10\
        );

    \I__4160\ : CascadeMux
    port map (
            O => \N__26252\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10_cascade_\
        );

    \I__4159\ : InMux
    port map (
            O => \N__26249\,
            I => \N__26246\
        );

    \I__4158\ : LocalMux
    port map (
            O => \N__26246\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\
        );

    \I__4157\ : InMux
    port map (
            O => \N__26243\,
            I => \N__26240\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__26240\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3\
        );

    \I__4155\ : CascadeMux
    port map (
            O => \N__26237\,
            I => \elapsed_time_ns_1_RNIL73T9_0_9_cascade_\
        );

    \I__4154\ : InMux
    port map (
            O => \N__26234\,
            I => \N__26231\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__26231\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\
        );

    \I__4152\ : InMux
    port map (
            O => \N__26228\,
            I => \N__26225\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__26225\,
            I => \N__26222\
        );

    \I__4150\ : Span4Mux_v
    port map (
            O => \N__26222\,
            I => \N__26219\
        );

    \I__4149\ : Odrv4
    port map (
            O => \N__26219\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22\
        );

    \I__4148\ : CascadeMux
    port map (
            O => \N__26216\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23_cascade_\
        );

    \I__4147\ : CascadeMux
    port map (
            O => \N__26213\,
            I => \N__26210\
        );

    \I__4146\ : InMux
    port map (
            O => \N__26210\,
            I => \N__26204\
        );

    \I__4145\ : InMux
    port map (
            O => \N__26209\,
            I => \N__26204\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__26204\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_23\
        );

    \I__4143\ : CascadeMux
    port map (
            O => \N__26201\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22_cascade_\
        );

    \I__4142\ : InMux
    port map (
            O => \N__26198\,
            I => \N__26192\
        );

    \I__4141\ : InMux
    port map (
            O => \N__26197\,
            I => \N__26192\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__26192\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_22\
        );

    \I__4139\ : InMux
    port map (
            O => \N__26189\,
            I => \N__26186\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__26186\,
            I => \N__26181\
        );

    \I__4137\ : InMux
    port map (
            O => \N__26185\,
            I => \N__26178\
        );

    \I__4136\ : InMux
    port map (
            O => \N__26184\,
            I => \N__26175\
        );

    \I__4135\ : Span4Mux_v
    port map (
            O => \N__26181\,
            I => \N__26170\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__26178\,
            I => \N__26170\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__26175\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4\
        );

    \I__4132\ : Odrv4
    port map (
            O => \N__26170\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4\
        );

    \I__4131\ : InMux
    port map (
            O => \N__26165\,
            I => \N__26162\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__26162\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\
        );

    \I__4129\ : InMux
    port map (
            O => \N__26159\,
            I => \N__26155\
        );

    \I__4128\ : InMux
    port map (
            O => \N__26158\,
            I => \N__26152\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__26155\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22\
        );

    \I__4126\ : LocalMux
    port map (
            O => \N__26152\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22\
        );

    \I__4125\ : InMux
    port map (
            O => \N__26147\,
            I => \N__26141\
        );

    \I__4124\ : InMux
    port map (
            O => \N__26146\,
            I => \N__26141\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__26141\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_22\
        );

    \I__4122\ : InMux
    port map (
            O => \N__26138\,
            I => \N__26134\
        );

    \I__4121\ : InMux
    port map (
            O => \N__26137\,
            I => \N__26131\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__26134\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__26131\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23\
        );

    \I__4118\ : CascadeMux
    port map (
            O => \N__26126\,
            I => \N__26123\
        );

    \I__4117\ : InMux
    port map (
            O => \N__26123\,
            I => \N__26117\
        );

    \I__4116\ : InMux
    port map (
            O => \N__26122\,
            I => \N__26117\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__26117\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_23\
        );

    \I__4114\ : CascadeMux
    port map (
            O => \N__26114\,
            I => \N__26111\
        );

    \I__4113\ : InMux
    port map (
            O => \N__26111\,
            I => \N__26105\
        );

    \I__4112\ : InMux
    port map (
            O => \N__26110\,
            I => \N__26105\
        );

    \I__4111\ : LocalMux
    port map (
            O => \N__26105\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\
        );

    \I__4110\ : InMux
    port map (
            O => \N__26102\,
            I => \N__26097\
        );

    \I__4109\ : InMux
    port map (
            O => \N__26101\,
            I => \N__26094\
        );

    \I__4108\ : InMux
    port map (
            O => \N__26100\,
            I => \N__26091\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__26097\,
            I => \N__26088\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__26094\,
            I => \N__26085\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__26091\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__4104\ : Odrv4
    port map (
            O => \N__26088\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__4103\ : Odrv4
    port map (
            O => \N__26085\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__4102\ : InMux
    port map (
            O => \N__26078\,
            I => \N__26074\
        );

    \I__4101\ : InMux
    port map (
            O => \N__26077\,
            I => \N__26070\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__26074\,
            I => \N__26067\
        );

    \I__4099\ : InMux
    port map (
            O => \N__26073\,
            I => \N__26064\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__26070\,
            I => \N__26061\
        );

    \I__4097\ : Span4Mux_h
    port map (
            O => \N__26067\,
            I => \N__26053\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__26064\,
            I => \N__26053\
        );

    \I__4095\ : Span4Mux_h
    port map (
            O => \N__26061\,
            I => \N__26053\
        );

    \I__4094\ : InMux
    port map (
            O => \N__26060\,
            I => \N__26050\
        );

    \I__4093\ : Span4Mux_v
    port map (
            O => \N__26053\,
            I => \N__26045\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__26050\,
            I => \N__26045\
        );

    \I__4091\ : Odrv4
    port map (
            O => \N__26045\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__4090\ : InMux
    port map (
            O => \N__26042\,
            I => \N__26038\
        );

    \I__4089\ : InMux
    port map (
            O => \N__26041\,
            I => \N__26034\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__26038\,
            I => \N__26031\
        );

    \I__4087\ : InMux
    port map (
            O => \N__26037\,
            I => \N__26028\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__26034\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3\
        );

    \I__4085\ : Odrv4
    port map (
            O => \N__26031\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__26028\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3\
        );

    \I__4083\ : InMux
    port map (
            O => \N__26021\,
            I => \N__26018\
        );

    \I__4082\ : LocalMux
    port map (
            O => \N__26018\,
            I => \N__26015\
        );

    \I__4081\ : Span4Mux_v
    port map (
            O => \N__26015\,
            I => \N__26011\
        );

    \I__4080\ : InMux
    port map (
            O => \N__26014\,
            I => \N__26008\
        );

    \I__4079\ : Odrv4
    port map (
            O => \N__26011\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__26008\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5\
        );

    \I__4077\ : CascadeMux
    port map (
            O => \N__26003\,
            I => \N__26000\
        );

    \I__4076\ : InMux
    port map (
            O => \N__26000\,
            I => \N__25997\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__25997\,
            I => \N__25994\
        );

    \I__4074\ : Span4Mux_v
    port map (
            O => \N__25994\,
            I => \N__25991\
        );

    \I__4073\ : Odrv4
    port map (
            O => \N__25991\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt22\
        );

    \I__4072\ : CascadeMux
    port map (
            O => \N__25988\,
            I => \N__25983\
        );

    \I__4071\ : InMux
    port map (
            O => \N__25987\,
            I => \N__25980\
        );

    \I__4070\ : InMux
    port map (
            O => \N__25986\,
            I => \N__25975\
        );

    \I__4069\ : InMux
    port map (
            O => \N__25983\,
            I => \N__25975\
        );

    \I__4068\ : LocalMux
    port map (
            O => \N__25980\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__25975\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__4066\ : InMux
    port map (
            O => \N__25970\,
            I => \N__25965\
        );

    \I__4065\ : InMux
    port map (
            O => \N__25969\,
            I => \N__25960\
        );

    \I__4064\ : InMux
    port map (
            O => \N__25968\,
            I => \N__25960\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__25965\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__25960\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__4061\ : InMux
    port map (
            O => \N__25955\,
            I => \N__25950\
        );

    \I__4060\ : InMux
    port map (
            O => \N__25954\,
            I => \N__25947\
        );

    \I__4059\ : InMux
    port map (
            O => \N__25953\,
            I => \N__25944\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__25950\,
            I => \N__25941\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__25947\,
            I => \N__25938\
        );

    \I__4056\ : LocalMux
    port map (
            O => \N__25944\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__4055\ : Odrv4
    port map (
            O => \N__25941\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__4054\ : Odrv4
    port map (
            O => \N__25938\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__4053\ : CascadeMux
    port map (
            O => \N__25931\,
            I => \N__25928\
        );

    \I__4052\ : InMux
    port map (
            O => \N__25928\,
            I => \N__25923\
        );

    \I__4051\ : InMux
    port map (
            O => \N__25927\,
            I => \N__25920\
        );

    \I__4050\ : InMux
    port map (
            O => \N__25926\,
            I => \N__25917\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__25923\,
            I => \N__25914\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__25920\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__4047\ : LocalMux
    port map (
            O => \N__25917\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__4046\ : Odrv4
    port map (
            O => \N__25914\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__4045\ : CascadeMux
    port map (
            O => \N__25907\,
            I => \N__25904\
        );

    \I__4044\ : InMux
    port map (
            O => \N__25904\,
            I => \N__25900\
        );

    \I__4043\ : InMux
    port map (
            O => \N__25903\,
            I => \N__25897\
        );

    \I__4042\ : LocalMux
    port map (
            O => \N__25900\,
            I => \N__25894\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__25897\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\
        );

    \I__4040\ : Odrv4
    port map (
            O => \N__25894\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\
        );

    \I__4039\ : InMux
    port map (
            O => \N__25889\,
            I => \N__25885\
        );

    \I__4038\ : InMux
    port map (
            O => \N__25888\,
            I => \N__25882\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__25885\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__25882\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\
        );

    \I__4035\ : CascadeMux
    port map (
            O => \N__25877\,
            I => \N__25874\
        );

    \I__4034\ : InMux
    port map (
            O => \N__25874\,
            I => \N__25871\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__25871\,
            I => \N__25868\
        );

    \I__4032\ : Sp12to4
    port map (
            O => \N__25868\,
            I => \N__25865\
        );

    \I__4031\ : Odrv12
    port map (
            O => \N__25865\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt16\
        );

    \I__4030\ : InMux
    port map (
            O => \N__25862\,
            I => \N__25859\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__25859\,
            I => \N__25856\
        );

    \I__4028\ : Span4Mux_v
    port map (
            O => \N__25856\,
            I => \N__25853\
        );

    \I__4027\ : Odrv4
    port map (
            O => \N__25853\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt18\
        );

    \I__4026\ : CascadeMux
    port map (
            O => \N__25850\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18_cascade_\
        );

    \I__4025\ : InMux
    port map (
            O => \N__25847\,
            I => \N__25841\
        );

    \I__4024\ : InMux
    port map (
            O => \N__25846\,
            I => \N__25841\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__25841\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\
        );

    \I__4022\ : InMux
    port map (
            O => \N__25838\,
            I => \N__25833\
        );

    \I__4021\ : InMux
    port map (
            O => \N__25837\,
            I => \N__25828\
        );

    \I__4020\ : InMux
    port map (
            O => \N__25836\,
            I => \N__25828\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__25833\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__25828\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__4017\ : InMux
    port map (
            O => \N__25823\,
            I => \N__25818\
        );

    \I__4016\ : InMux
    port map (
            O => \N__25822\,
            I => \N__25813\
        );

    \I__4015\ : InMux
    port map (
            O => \N__25821\,
            I => \N__25813\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__25818\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__25813\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__4012\ : CascadeMux
    port map (
            O => \N__25808\,
            I => \N__25805\
        );

    \I__4011\ : InMux
    port map (
            O => \N__25805\,
            I => \N__25802\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__25802\,
            I => \N__25799\
        );

    \I__4009\ : Span4Mux_v
    port map (
            O => \N__25799\,
            I => \N__25796\
        );

    \I__4008\ : Odrv4
    port map (
            O => \N__25796\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\
        );

    \I__4007\ : CascadeMux
    port map (
            O => \N__25793\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15_cascade_\
        );

    \I__4006\ : InMux
    port map (
            O => \N__25790\,
            I => \N__25787\
        );

    \I__4005\ : LocalMux
    port map (
            O => \N__25787\,
            I => \N__25784\
        );

    \I__4004\ : Span4Mux_v
    port map (
            O => \N__25784\,
            I => \N__25781\
        );

    \I__4003\ : Odrv4
    port map (
            O => \N__25781\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\
        );

    \I__4002\ : CascadeMux
    port map (
            O => \N__25778\,
            I => \N__25775\
        );

    \I__4001\ : InMux
    port map (
            O => \N__25775\,
            I => \N__25772\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__25772\,
            I => \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2\
        );

    \I__3999\ : InMux
    port map (
            O => \N__25769\,
            I => \N__25766\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__25766\,
            I => \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2\
        );

    \I__3997\ : InMux
    port map (
            O => \N__25763\,
            I => \N__25760\
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__25760\,
            I => \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033\
        );

    \I__3995\ : CascadeMux
    port map (
            O => \N__25757\,
            I => \N__25754\
        );

    \I__3994\ : InMux
    port map (
            O => \N__25754\,
            I => \N__25751\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__25751\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433\
        );

    \I__3992\ : InMux
    port map (
            O => \N__25748\,
            I => \N__25745\
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__25745\,
            I => \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2\
        );

    \I__3990\ : InMux
    port map (
            O => \N__25742\,
            I => \N__25739\
        );

    \I__3989\ : LocalMux
    port map (
            O => \N__25739\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93\
        );

    \I__3988\ : InMux
    port map (
            O => \N__25736\,
            I => \N__25721\
        );

    \I__3987\ : InMux
    port map (
            O => \N__25735\,
            I => \N__25721\
        );

    \I__3986\ : InMux
    port map (
            O => \N__25734\,
            I => \N__25721\
        );

    \I__3985\ : InMux
    port map (
            O => \N__25733\,
            I => \N__25721\
        );

    \I__3984\ : InMux
    port map (
            O => \N__25732\,
            I => \N__25721\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__25721\,
            I => \N__25713\
        );

    \I__3982\ : InMux
    port map (
            O => \N__25720\,
            I => \N__25702\
        );

    \I__3981\ : InMux
    port map (
            O => \N__25719\,
            I => \N__25702\
        );

    \I__3980\ : InMux
    port map (
            O => \N__25718\,
            I => \N__25702\
        );

    \I__3979\ : InMux
    port map (
            O => \N__25717\,
            I => \N__25702\
        );

    \I__3978\ : InMux
    port map (
            O => \N__25716\,
            I => \N__25702\
        );

    \I__3977\ : Sp12to4
    port map (
            O => \N__25713\,
            I => \N__25697\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__25702\,
            I => \N__25697\
        );

    \I__3975\ : Span12Mux_s7_v
    port map (
            O => \N__25697\,
            I => \N__25694\
        );

    \I__3974\ : Odrv12
    port map (
            O => \N__25694\,
            I => \pwm_generator_inst.N_17\
        );

    \I__3973\ : InMux
    port map (
            O => \N__25691\,
            I => \N__25671\
        );

    \I__3972\ : InMux
    port map (
            O => \N__25690\,
            I => \N__25671\
        );

    \I__3971\ : InMux
    port map (
            O => \N__25689\,
            I => \N__25671\
        );

    \I__3970\ : InMux
    port map (
            O => \N__25688\,
            I => \N__25671\
        );

    \I__3969\ : InMux
    port map (
            O => \N__25687\,
            I => \N__25671\
        );

    \I__3968\ : InMux
    port map (
            O => \N__25686\,
            I => \N__25660\
        );

    \I__3967\ : InMux
    port map (
            O => \N__25685\,
            I => \N__25660\
        );

    \I__3966\ : InMux
    port map (
            O => \N__25684\,
            I => \N__25660\
        );

    \I__3965\ : InMux
    port map (
            O => \N__25683\,
            I => \N__25660\
        );

    \I__3964\ : InMux
    port map (
            O => \N__25682\,
            I => \N__25660\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__25671\,
            I => \N__25657\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__25660\,
            I => \N__25654\
        );

    \I__3961\ : Span4Mux_h
    port map (
            O => \N__25657\,
            I => \N__25649\
        );

    \I__3960\ : Span4Mux_v
    port map (
            O => \N__25654\,
            I => \N__25649\
        );

    \I__3959\ : Span4Mux_h
    port map (
            O => \N__25649\,
            I => \N__25646\
        );

    \I__3958\ : Odrv4
    port map (
            O => \N__25646\,
            I => \pwm_generator_inst.N_16\
        );

    \I__3957\ : CascadeMux
    port map (
            O => \N__25643\,
            I => \N__25640\
        );

    \I__3956\ : InMux
    port map (
            O => \N__25640\,
            I => \N__25637\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__25637\,
            I => \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2\
        );

    \I__3954\ : InMux
    port map (
            O => \N__25634\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_8\
        );

    \I__3953\ : InMux
    port map (
            O => \N__25631\,
            I => \N__25628\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__25628\,
            I => \N__25624\
        );

    \I__3951\ : InMux
    port map (
            O => \N__25627\,
            I => \N__25621\
        );

    \I__3950\ : Span4Mux_v
    port map (
            O => \N__25624\,
            I => \N__25618\
        );

    \I__3949\ : LocalMux
    port map (
            O => \N__25621\,
            I => \N__25615\
        );

    \I__3948\ : Sp12to4
    port map (
            O => \N__25618\,
            I => \N__25612\
        );

    \I__3947\ : Span4Mux_h
    port map (
            O => \N__25615\,
            I => \N__25609\
        );

    \I__3946\ : Span12Mux_s8_h
    port map (
            O => \N__25612\,
            I => \N__25606\
        );

    \I__3945\ : Odrv4
    port map (
            O => \N__25609\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__3944\ : Odrv12
    port map (
            O => \N__25606\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__3943\ : InMux
    port map (
            O => \N__25601\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_9\
        );

    \I__3942\ : InMux
    port map (
            O => \N__25598\,
            I => \N__25594\
        );

    \I__3941\ : InMux
    port map (
            O => \N__25597\,
            I => \N__25591\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__25594\,
            I => \N__25588\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__25591\,
            I => \N__25585\
        );

    \I__3938\ : Span12Mux_s8_h
    port map (
            O => \N__25588\,
            I => \N__25582\
        );

    \I__3937\ : Span4Mux_v
    port map (
            O => \N__25585\,
            I => \N__25579\
        );

    \I__3936\ : Span12Mux_v
    port map (
            O => \N__25582\,
            I => \N__25576\
        );

    \I__3935\ : Odrv4
    port map (
            O => \N__25579\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__3934\ : Odrv12
    port map (
            O => \N__25576\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__3933\ : InMux
    port map (
            O => \N__25571\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_10\
        );

    \I__3932\ : InMux
    port map (
            O => \N__25568\,
            I => \N__25564\
        );

    \I__3931\ : InMux
    port map (
            O => \N__25567\,
            I => \N__25561\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__25564\,
            I => \N__25558\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__25561\,
            I => \N__25555\
        );

    \I__3928\ : Span12Mux_s7_v
    port map (
            O => \N__25558\,
            I => \N__25552\
        );

    \I__3927\ : Span4Mux_h
    port map (
            O => \N__25555\,
            I => \N__25549\
        );

    \I__3926\ : Span12Mux_v
    port map (
            O => \N__25552\,
            I => \N__25546\
        );

    \I__3925\ : Odrv4
    port map (
            O => \N__25549\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__3924\ : Odrv12
    port map (
            O => \N__25546\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__3923\ : InMux
    port map (
            O => \N__25541\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_11\
        );

    \I__3922\ : InMux
    port map (
            O => \N__25538\,
            I => \N__25535\
        );

    \I__3921\ : LocalMux
    port map (
            O => \N__25535\,
            I => \N__25532\
        );

    \I__3920\ : Span4Mux_v
    port map (
            O => \N__25532\,
            I => \N__25528\
        );

    \I__3919\ : InMux
    port map (
            O => \N__25531\,
            I => \N__25525\
        );

    \I__3918\ : Span4Mux_v
    port map (
            O => \N__25528\,
            I => \N__25522\
        );

    \I__3917\ : LocalMux
    port map (
            O => \N__25525\,
            I => \N__25519\
        );

    \I__3916\ : Sp12to4
    port map (
            O => \N__25522\,
            I => \N__25516\
        );

    \I__3915\ : Span4Mux_h
    port map (
            O => \N__25519\,
            I => \N__25513\
        );

    \I__3914\ : Span12Mux_s8_h
    port map (
            O => \N__25516\,
            I => \N__25510\
        );

    \I__3913\ : Odrv4
    port map (
            O => \N__25513\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_13\
        );

    \I__3912\ : Odrv12
    port map (
            O => \N__25510\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_13\
        );

    \I__3911\ : InMux
    port map (
            O => \N__25505\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_12\
        );

    \I__3910\ : InMux
    port map (
            O => \N__25502\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_13\
        );

    \I__3909\ : InMux
    port map (
            O => \N__25499\,
            I => \N__25480\
        );

    \I__3908\ : InMux
    port map (
            O => \N__25498\,
            I => \N__25463\
        );

    \I__3907\ : InMux
    port map (
            O => \N__25497\,
            I => \N__25463\
        );

    \I__3906\ : InMux
    port map (
            O => \N__25496\,
            I => \N__25463\
        );

    \I__3905\ : InMux
    port map (
            O => \N__25495\,
            I => \N__25463\
        );

    \I__3904\ : InMux
    port map (
            O => \N__25494\,
            I => \N__25463\
        );

    \I__3903\ : InMux
    port map (
            O => \N__25493\,
            I => \N__25463\
        );

    \I__3902\ : InMux
    port map (
            O => \N__25492\,
            I => \N__25463\
        );

    \I__3901\ : InMux
    port map (
            O => \N__25491\,
            I => \N__25463\
        );

    \I__3900\ : InMux
    port map (
            O => \N__25490\,
            I => \N__25446\
        );

    \I__3899\ : InMux
    port map (
            O => \N__25489\,
            I => \N__25446\
        );

    \I__3898\ : InMux
    port map (
            O => \N__25488\,
            I => \N__25446\
        );

    \I__3897\ : InMux
    port map (
            O => \N__25487\,
            I => \N__25446\
        );

    \I__3896\ : InMux
    port map (
            O => \N__25486\,
            I => \N__25446\
        );

    \I__3895\ : InMux
    port map (
            O => \N__25485\,
            I => \N__25446\
        );

    \I__3894\ : InMux
    port map (
            O => \N__25484\,
            I => \N__25446\
        );

    \I__3893\ : InMux
    port map (
            O => \N__25483\,
            I => \N__25446\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__25480\,
            I => \N__25443\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__25463\,
            I => \N__25435\
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__25446\,
            I => \N__25435\
        );

    \I__3889\ : Span4Mux_v
    port map (
            O => \N__25443\,
            I => \N__25435\
        );

    \I__3888\ : InMux
    port map (
            O => \N__25442\,
            I => \N__25432\
        );

    \I__3887\ : Span4Mux_v
    port map (
            O => \N__25435\,
            I => \N__25429\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__25432\,
            I => \N__25426\
        );

    \I__3885\ : Sp12to4
    port map (
            O => \N__25429\,
            I => \N__25423\
        );

    \I__3884\ : Span4Mux_h
    port map (
            O => \N__25426\,
            I => \N__25420\
        );

    \I__3883\ : Span12Mux_s8_h
    port map (
            O => \N__25423\,
            I => \N__25417\
        );

    \I__3882\ : Odrv4
    port map (
            O => \N__25420\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__3881\ : Odrv12
    port map (
            O => \N__25417\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__3880\ : CascadeMux
    port map (
            O => \N__25412\,
            I => \N__25409\
        );

    \I__3879\ : InMux
    port map (
            O => \N__25409\,
            I => \N__25406\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__25406\,
            I => \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23\
        );

    \I__3877\ : CascadeMux
    port map (
            O => \N__25403\,
            I => \N__25400\
        );

    \I__3876\ : InMux
    port map (
            O => \N__25400\,
            I => \N__25397\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__25397\,
            I => \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23\
        );

    \I__3874\ : CascadeMux
    port map (
            O => \N__25394\,
            I => \N__25391\
        );

    \I__3873\ : InMux
    port map (
            O => \N__25391\,
            I => \N__25388\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__25388\,
            I => \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2\
        );

    \I__3871\ : InMux
    port map (
            O => \N__25385\,
            I => \N__25381\
        );

    \I__3870\ : InMux
    port map (
            O => \N__25384\,
            I => \N__25378\
        );

    \I__3869\ : LocalMux
    port map (
            O => \N__25381\,
            I => \N__25375\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__25378\,
            I => \N__25372\
        );

    \I__3867\ : Span4Mux_v
    port map (
            O => \N__25375\,
            I => \N__25369\
        );

    \I__3866\ : Span12Mux_s3_h
    port map (
            O => \N__25372\,
            I => \N__25366\
        );

    \I__3865\ : Sp12to4
    port map (
            O => \N__25369\,
            I => \N__25361\
        );

    \I__3864\ : Span12Mux_v
    port map (
            O => \N__25366\,
            I => \N__25361\
        );

    \I__3863\ : Odrv12
    port map (
            O => \N__25361\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_1\
        );

    \I__3862\ : InMux
    port map (
            O => \N__25358\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_0\
        );

    \I__3861\ : InMux
    port map (
            O => \N__25355\,
            I => \N__25351\
        );

    \I__3860\ : InMux
    port map (
            O => \N__25354\,
            I => \N__25348\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__25351\,
            I => \N__25345\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__25348\,
            I => \N__25342\
        );

    \I__3857\ : Span12Mux_s2_h
    port map (
            O => \N__25345\,
            I => \N__25339\
        );

    \I__3856\ : Span4Mux_v
    port map (
            O => \N__25342\,
            I => \N__25336\
        );

    \I__3855\ : Span12Mux_v
    port map (
            O => \N__25339\,
            I => \N__25333\
        );

    \I__3854\ : Odrv4
    port map (
            O => \N__25336\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__3853\ : Odrv12
    port map (
            O => \N__25333\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__3852\ : InMux
    port map (
            O => \N__25328\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_1\
        );

    \I__3851\ : InMux
    port map (
            O => \N__25325\,
            I => \N__25321\
        );

    \I__3850\ : InMux
    port map (
            O => \N__25324\,
            I => \N__25318\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__25321\,
            I => \N__25315\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__25318\,
            I => \N__25312\
        );

    \I__3847\ : Span12Mux_s1_h
    port map (
            O => \N__25315\,
            I => \N__25309\
        );

    \I__3846\ : Span4Mux_v
    port map (
            O => \N__25312\,
            I => \N__25306\
        );

    \I__3845\ : Span12Mux_v
    port map (
            O => \N__25309\,
            I => \N__25303\
        );

    \I__3844\ : Odrv4
    port map (
            O => \N__25306\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__3843\ : Odrv12
    port map (
            O => \N__25303\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__3842\ : InMux
    port map (
            O => \N__25298\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_2\
        );

    \I__3841\ : InMux
    port map (
            O => \N__25295\,
            I => \N__25291\
        );

    \I__3840\ : InMux
    port map (
            O => \N__25294\,
            I => \N__25288\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__25291\,
            I => \N__25285\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__25288\,
            I => \N__25282\
        );

    \I__3837\ : Span12Mux_s8_h
    port map (
            O => \N__25285\,
            I => \N__25279\
        );

    \I__3836\ : Span4Mux_h
    port map (
            O => \N__25282\,
            I => \N__25276\
        );

    \I__3835\ : Span12Mux_v
    port map (
            O => \N__25279\,
            I => \N__25273\
        );

    \I__3834\ : Odrv4
    port map (
            O => \N__25276\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__3833\ : Odrv12
    port map (
            O => \N__25273\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__3832\ : InMux
    port map (
            O => \N__25268\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_3\
        );

    \I__3831\ : InMux
    port map (
            O => \N__25265\,
            I => \N__25262\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__25262\,
            I => \N__25258\
        );

    \I__3829\ : InMux
    port map (
            O => \N__25261\,
            I => \N__25255\
        );

    \I__3828\ : Sp12to4
    port map (
            O => \N__25258\,
            I => \N__25252\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__25255\,
            I => \N__25249\
        );

    \I__3826\ : Span12Mux_s11_h
    port map (
            O => \N__25252\,
            I => \N__25246\
        );

    \I__3825\ : Span4Mux_h
    port map (
            O => \N__25249\,
            I => \N__25243\
        );

    \I__3824\ : Span12Mux_v
    port map (
            O => \N__25246\,
            I => \N__25240\
        );

    \I__3823\ : Odrv4
    port map (
            O => \N__25243\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__3822\ : Odrv12
    port map (
            O => \N__25240\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__3821\ : InMux
    port map (
            O => \N__25235\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_4\
        );

    \I__3820\ : InMux
    port map (
            O => \N__25232\,
            I => \N__25229\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__25229\,
            I => \N__25225\
        );

    \I__3818\ : InMux
    port map (
            O => \N__25228\,
            I => \N__25222\
        );

    \I__3817\ : Sp12to4
    port map (
            O => \N__25225\,
            I => \N__25219\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__25222\,
            I => \N__25216\
        );

    \I__3815\ : Span12Mux_s10_h
    port map (
            O => \N__25219\,
            I => \N__25213\
        );

    \I__3814\ : Span4Mux_h
    port map (
            O => \N__25216\,
            I => \N__25210\
        );

    \I__3813\ : Span12Mux_v
    port map (
            O => \N__25213\,
            I => \N__25207\
        );

    \I__3812\ : Odrv4
    port map (
            O => \N__25210\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__3811\ : Odrv12
    port map (
            O => \N__25207\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__3810\ : InMux
    port map (
            O => \N__25202\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_5\
        );

    \I__3809\ : InMux
    port map (
            O => \N__25199\,
            I => \N__25196\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__25196\,
            I => \N__25192\
        );

    \I__3807\ : InMux
    port map (
            O => \N__25195\,
            I => \N__25189\
        );

    \I__3806\ : Sp12to4
    port map (
            O => \N__25192\,
            I => \N__25186\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__25189\,
            I => \N__25183\
        );

    \I__3804\ : Span12Mux_s5_h
    port map (
            O => \N__25186\,
            I => \N__25180\
        );

    \I__3803\ : Span4Mux_h
    port map (
            O => \N__25183\,
            I => \N__25177\
        );

    \I__3802\ : Span12Mux_v
    port map (
            O => \N__25180\,
            I => \N__25174\
        );

    \I__3801\ : Odrv4
    port map (
            O => \N__25177\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__3800\ : Odrv12
    port map (
            O => \N__25174\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__3799\ : InMux
    port map (
            O => \N__25169\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_6\
        );

    \I__3798\ : InMux
    port map (
            O => \N__25166\,
            I => \N__25163\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__25163\,
            I => \N__25160\
        );

    \I__3796\ : Span4Mux_v
    port map (
            O => \N__25160\,
            I => \N__25156\
        );

    \I__3795\ : InMux
    port map (
            O => \N__25159\,
            I => \N__25153\
        );

    \I__3794\ : Sp12to4
    port map (
            O => \N__25156\,
            I => \N__25150\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__25153\,
            I => \N__25145\
        );

    \I__3792\ : Span12Mux_s4_h
    port map (
            O => \N__25150\,
            I => \N__25145\
        );

    \I__3791\ : Span12Mux_v
    port map (
            O => \N__25145\,
            I => \N__25142\
        );

    \I__3790\ : Odrv12
    port map (
            O => \N__25142\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__3789\ : InMux
    port map (
            O => \N__25139\,
            I => \bfn_8_20_0_\
        );

    \I__3788\ : InMux
    port map (
            O => \N__25136\,
            I => \N__25133\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__25133\,
            I => \N__25129\
        );

    \I__3786\ : InMux
    port map (
            O => \N__25132\,
            I => \N__25126\
        );

    \I__3785\ : Span4Mux_v
    port map (
            O => \N__25129\,
            I => \N__25123\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__25126\,
            I => \N__25120\
        );

    \I__3783\ : Sp12to4
    port map (
            O => \N__25123\,
            I => \N__25117\
        );

    \I__3782\ : Span4Mux_h
    port map (
            O => \N__25120\,
            I => \N__25114\
        );

    \I__3781\ : Span12Mux_s8_h
    port map (
            O => \N__25117\,
            I => \N__25111\
        );

    \I__3780\ : Odrv4
    port map (
            O => \N__25114\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__3779\ : Odrv12
    port map (
            O => \N__25111\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__3778\ : InMux
    port map (
            O => \N__25106\,
            I => \N__25100\
        );

    \I__3777\ : InMux
    port map (
            O => \N__25105\,
            I => \N__25100\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__25100\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_27\
        );

    \I__3775\ : CascadeMux
    port map (
            O => \N__25097\,
            I => \N__25094\
        );

    \I__3774\ : InMux
    port map (
            O => \N__25094\,
            I => \N__25087\
        );

    \I__3773\ : InMux
    port map (
            O => \N__25093\,
            I => \N__25087\
        );

    \I__3772\ : InMux
    port map (
            O => \N__25092\,
            I => \N__25084\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__25087\,
            I => \N__25081\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__25084\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__3769\ : Odrv12
    port map (
            O => \N__25081\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__3768\ : CascadeMux
    port map (
            O => \N__25076\,
            I => \N__25072\
        );

    \I__3767\ : InMux
    port map (
            O => \N__25075\,
            I => \N__25066\
        );

    \I__3766\ : InMux
    port map (
            O => \N__25072\,
            I => \N__25066\
        );

    \I__3765\ : InMux
    port map (
            O => \N__25071\,
            I => \N__25063\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__25066\,
            I => \N__25060\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__25063\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__3762\ : Odrv12
    port map (
            O => \N__25060\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__3761\ : CascadeMux
    port map (
            O => \N__25055\,
            I => \N__25052\
        );

    \I__3760\ : InMux
    port map (
            O => \N__25052\,
            I => \N__25049\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__25049\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt26\
        );

    \I__3758\ : InMux
    port map (
            O => \N__25046\,
            I => \N__25043\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__25043\,
            I => \N__25040\
        );

    \I__3756\ : Span4Mux_h
    port map (
            O => \N__25040\,
            I => \N__25037\
        );

    \I__3755\ : Odrv4
    port map (
            O => \N__25037\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\
        );

    \I__3754\ : CascadeMux
    port map (
            O => \N__25034\,
            I => \N__25031\
        );

    \I__3753\ : InMux
    port map (
            O => \N__25031\,
            I => \N__25025\
        );

    \I__3752\ : InMux
    port map (
            O => \N__25030\,
            I => \N__25025\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__25025\,
            I => \N__25022\
        );

    \I__3750\ : Odrv4
    port map (
            O => \N__25022\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_20\
        );

    \I__3749\ : CascadeMux
    port map (
            O => \N__25019\,
            I => \N__25016\
        );

    \I__3748\ : InMux
    port map (
            O => \N__25016\,
            I => \N__25013\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__25013\,
            I => \N__25009\
        );

    \I__3746\ : InMux
    port map (
            O => \N__25012\,
            I => \N__25006\
        );

    \I__3745\ : Span4Mux_h
    port map (
            O => \N__25009\,
            I => \N__25003\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__25006\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\
        );

    \I__3743\ : Odrv4
    port map (
            O => \N__25003\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\
        );

    \I__3742\ : InMux
    port map (
            O => \N__24998\,
            I => \N__24994\
        );

    \I__3741\ : InMux
    port map (
            O => \N__24997\,
            I => \N__24991\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__24994\,
            I => \N__24988\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__24991\,
            I => \N__24985\
        );

    \I__3738\ : Sp12to4
    port map (
            O => \N__24988\,
            I => \N__24982\
        );

    \I__3737\ : Span12Mux_v
    port map (
            O => \N__24985\,
            I => \N__24977\
        );

    \I__3736\ : Span12Mux_v
    port map (
            O => \N__24982\,
            I => \N__24977\
        );

    \I__3735\ : Odrv12
    port map (
            O => \N__24977\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__3734\ : InMux
    port map (
            O => \N__24974\,
            I => \N__24971\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__24971\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axb_0\
        );

    \I__3732\ : InMux
    port map (
            O => \N__24968\,
            I => \N__24965\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__24965\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt24\
        );

    \I__3730\ : CascadeMux
    port map (
            O => \N__24962\,
            I => \N__24959\
        );

    \I__3729\ : InMux
    port map (
            O => \N__24959\,
            I => \N__24956\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__24956\,
            I => \N__24953\
        );

    \I__3727\ : Odrv4
    port map (
            O => \N__24953\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24\
        );

    \I__3726\ : InMux
    port map (
            O => \N__24950\,
            I => \N__24947\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__24947\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\
        );

    \I__3724\ : CascadeMux
    port map (
            O => \N__24944\,
            I => \N__24941\
        );

    \I__3723\ : InMux
    port map (
            O => \N__24941\,
            I => \N__24938\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__24938\,
            I => \N__24934\
        );

    \I__3721\ : InMux
    port map (
            O => \N__24937\,
            I => \N__24931\
        );

    \I__3720\ : Odrv4
    port map (
            O => \N__24934\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt30\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__24931\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt30\
        );

    \I__3718\ : InMux
    port map (
            O => \N__24926\,
            I => \N__24923\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__24923\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO\
        );

    \I__3716\ : InMux
    port map (
            O => \N__24920\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_28\
        );

    \I__3715\ : InMux
    port map (
            O => \N__24917\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30\
        );

    \I__3714\ : InMux
    port map (
            O => \N__24914\,
            I => \N__24910\
        );

    \I__3713\ : InMux
    port map (
            O => \N__24913\,
            I => \N__24907\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__24910\,
            I => \N__24904\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__24907\,
            I => \N__24901\
        );

    \I__3710\ : Span4Mux_h
    port map (
            O => \N__24904\,
            I => \N__24898\
        );

    \I__3709\ : Span4Mux_h
    port map (
            O => \N__24901\,
            I => \N__24895\
        );

    \I__3708\ : Odrv4
    port map (
            O => \N__24898\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__3707\ : Odrv4
    port map (
            O => \N__24895\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__3706\ : CascadeMux
    port map (
            O => \N__24890\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27_cascade_\
        );

    \I__3705\ : InMux
    port map (
            O => \N__24887\,
            I => \N__24884\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__24884\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26\
        );

    \I__3703\ : InMux
    port map (
            O => \N__24881\,
            I => \N__24877\
        );

    \I__3702\ : InMux
    port map (
            O => \N__24880\,
            I => \N__24874\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__24877\,
            I => \N__24871\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__24874\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__3699\ : Odrv12
    port map (
            O => \N__24871\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__3698\ : CascadeMux
    port map (
            O => \N__24866\,
            I => \N__24863\
        );

    \I__3697\ : InMux
    port map (
            O => \N__24863\,
            I => \N__24860\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__24860\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\
        );

    \I__3695\ : InMux
    port map (
            O => \N__24857\,
            I => \N__24854\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__24854\,
            I => \N__24850\
        );

    \I__3693\ : InMux
    port map (
            O => \N__24853\,
            I => \N__24847\
        );

    \I__3692\ : Span4Mux_v
    port map (
            O => \N__24850\,
            I => \N__24844\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__24847\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__3690\ : Odrv4
    port map (
            O => \N__24844\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__3689\ : CascadeMux
    port map (
            O => \N__24839\,
            I => \N__24836\
        );

    \I__3688\ : InMux
    port map (
            O => \N__24836\,
            I => \N__24833\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__24833\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\
        );

    \I__3686\ : InMux
    port map (
            O => \N__24830\,
            I => \N__24826\
        );

    \I__3685\ : InMux
    port map (
            O => \N__24829\,
            I => \N__24823\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__24826\,
            I => \N__24820\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__24823\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__3682\ : Odrv12
    port map (
            O => \N__24820\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__3681\ : CascadeMux
    port map (
            O => \N__24815\,
            I => \N__24812\
        );

    \I__3680\ : InMux
    port map (
            O => \N__24812\,
            I => \N__24809\
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__24809\,
            I => \N__24806\
        );

    \I__3678\ : Odrv4
    port map (
            O => \N__24806\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\
        );

    \I__3677\ : InMux
    port map (
            O => \N__24803\,
            I => \N__24799\
        );

    \I__3676\ : InMux
    port map (
            O => \N__24802\,
            I => \N__24796\
        );

    \I__3675\ : LocalMux
    port map (
            O => \N__24799\,
            I => \N__24793\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__24796\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__3673\ : Odrv12
    port map (
            O => \N__24793\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__3672\ : InMux
    port map (
            O => \N__24788\,
            I => \N__24785\
        );

    \I__3671\ : LocalMux
    port map (
            O => \N__24785\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\
        );

    \I__3670\ : InMux
    port map (
            O => \N__24782\,
            I => \N__24778\
        );

    \I__3669\ : InMux
    port map (
            O => \N__24781\,
            I => \N__24775\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__24778\,
            I => \N__24772\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__24775\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__3666\ : Odrv12
    port map (
            O => \N__24772\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__3665\ : CascadeMux
    port map (
            O => \N__24767\,
            I => \N__24764\
        );

    \I__3664\ : InMux
    port map (
            O => \N__24764\,
            I => \N__24761\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__24761\,
            I => \N__24758\
        );

    \I__3662\ : Odrv4
    port map (
            O => \N__24758\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\
        );

    \I__3661\ : InMux
    port map (
            O => \N__24755\,
            I => \N__24752\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__24752\,
            I => \N__24749\
        );

    \I__3659\ : Span4Mux_v
    port map (
            O => \N__24749\,
            I => \N__24746\
        );

    \I__3658\ : Odrv4
    port map (
            O => \N__24746\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\
        );

    \I__3657\ : InMux
    port map (
            O => \N__24743\,
            I => \N__24740\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__24740\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20\
        );

    \I__3655\ : CascadeMux
    port map (
            O => \N__24737\,
            I => \N__24734\
        );

    \I__3654\ : InMux
    port map (
            O => \N__24734\,
            I => \N__24731\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__24731\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt20\
        );

    \I__3652\ : InMux
    port map (
            O => \N__24728\,
            I => \N__24725\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__24725\,
            I => \N__24721\
        );

    \I__3650\ : InMux
    port map (
            O => \N__24724\,
            I => \N__24718\
        );

    \I__3649\ : Span4Mux_v
    port map (
            O => \N__24721\,
            I => \N__24715\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__24718\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__3647\ : Odrv4
    port map (
            O => \N__24715\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__3646\ : CascadeMux
    port map (
            O => \N__24710\,
            I => \N__24707\
        );

    \I__3645\ : InMux
    port map (
            O => \N__24707\,
            I => \N__24704\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__24704\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\
        );

    \I__3643\ : InMux
    port map (
            O => \N__24701\,
            I => \N__24697\
        );

    \I__3642\ : InMux
    port map (
            O => \N__24700\,
            I => \N__24694\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__24697\,
            I => \N__24691\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__24694\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__3639\ : Odrv12
    port map (
            O => \N__24691\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__3638\ : CascadeMux
    port map (
            O => \N__24686\,
            I => \N__24683\
        );

    \I__3637\ : InMux
    port map (
            O => \N__24683\,
            I => \N__24680\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__24680\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\
        );

    \I__3635\ : InMux
    port map (
            O => \N__24677\,
            I => \N__24674\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__24674\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\
        );

    \I__3633\ : InMux
    port map (
            O => \N__24671\,
            I => \N__24667\
        );

    \I__3632\ : InMux
    port map (
            O => \N__24670\,
            I => \N__24664\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__24667\,
            I => \N__24661\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__24664\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__3629\ : Odrv12
    port map (
            O => \N__24661\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__3628\ : InMux
    port map (
            O => \N__24656\,
            I => \N__24653\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__24653\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\
        );

    \I__3626\ : InMux
    port map (
            O => \N__24650\,
            I => \N__24646\
        );

    \I__3625\ : InMux
    port map (
            O => \N__24649\,
            I => \N__24643\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__24646\,
            I => \N__24640\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__24643\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__3622\ : Odrv12
    port map (
            O => \N__24640\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__3621\ : CascadeMux
    port map (
            O => \N__24635\,
            I => \N__24632\
        );

    \I__3620\ : InMux
    port map (
            O => \N__24632\,
            I => \N__24629\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__24629\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\
        );

    \I__3618\ : InMux
    port map (
            O => \N__24626\,
            I => \N__24622\
        );

    \I__3617\ : InMux
    port map (
            O => \N__24625\,
            I => \N__24619\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__24622\,
            I => \N__24616\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__24619\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__3614\ : Odrv12
    port map (
            O => \N__24616\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__3613\ : CascadeMux
    port map (
            O => \N__24611\,
            I => \N__24608\
        );

    \I__3612\ : InMux
    port map (
            O => \N__24608\,
            I => \N__24605\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__24605\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\
        );

    \I__3610\ : InMux
    port map (
            O => \N__24602\,
            I => \N__24598\
        );

    \I__3609\ : InMux
    port map (
            O => \N__24601\,
            I => \N__24595\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__24598\,
            I => \N__24592\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__24595\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__3606\ : Odrv12
    port map (
            O => \N__24592\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__3605\ : CascadeMux
    port map (
            O => \N__24587\,
            I => \N__24584\
        );

    \I__3604\ : InMux
    port map (
            O => \N__24584\,
            I => \N__24581\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__24581\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\
        );

    \I__3602\ : InMux
    port map (
            O => \N__24578\,
            I => \N__24574\
        );

    \I__3601\ : InMux
    port map (
            O => \N__24577\,
            I => \N__24571\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__24574\,
            I => \N__24568\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__24571\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__3598\ : Odrv12
    port map (
            O => \N__24568\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__3597\ : CascadeMux
    port map (
            O => \N__24563\,
            I => \N__24560\
        );

    \I__3596\ : InMux
    port map (
            O => \N__24560\,
            I => \N__24557\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__24557\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\
        );

    \I__3594\ : InMux
    port map (
            O => \N__24554\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\
        );

    \I__3593\ : InMux
    port map (
            O => \N__24551\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\
        );

    \I__3592\ : InMux
    port map (
            O => \N__24548\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\
        );

    \I__3591\ : InMux
    port map (
            O => \N__24545\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\
        );

    \I__3590\ : InMux
    port map (
            O => \N__24542\,
            I => \N__24532\
        );

    \I__3589\ : InMux
    port map (
            O => \N__24541\,
            I => \N__24532\
        );

    \I__3588\ : InMux
    port map (
            O => \N__24540\,
            I => \N__24532\
        );

    \I__3587\ : InMux
    port map (
            O => \N__24539\,
            I => \N__24529\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__24532\,
            I => \N__24526\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__24529\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__3584\ : Odrv4
    port map (
            O => \N__24526\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__3583\ : InMux
    port map (
            O => \N__24521\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\
        );

    \I__3582\ : InMux
    port map (
            O => \N__24518\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\
        );

    \I__3581\ : InMux
    port map (
            O => \N__24515\,
            I => \N__24505\
        );

    \I__3580\ : InMux
    port map (
            O => \N__24514\,
            I => \N__24505\
        );

    \I__3579\ : InMux
    port map (
            O => \N__24513\,
            I => \N__24505\
        );

    \I__3578\ : InMux
    port map (
            O => \N__24512\,
            I => \N__24502\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__24505\,
            I => \N__24499\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__24502\,
            I => \N__24494\
        );

    \I__3575\ : Span4Mux_v
    port map (
            O => \N__24499\,
            I => \N__24494\
        );

    \I__3574\ : Odrv4
    port map (
            O => \N__24494\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__3573\ : InMux
    port map (
            O => \N__24491\,
            I => \N__24488\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__24488\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\
        );

    \I__3571\ : CascadeMux
    port map (
            O => \N__24485\,
            I => \N__24482\
        );

    \I__3570\ : InMux
    port map (
            O => \N__24482\,
            I => \N__24479\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__24479\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\
        );

    \I__3568\ : InMux
    port map (
            O => \N__24476\,
            I => \N__24473\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__24473\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\
        );

    \I__3566\ : InMux
    port map (
            O => \N__24470\,
            I => \N__24466\
        );

    \I__3565\ : InMux
    port map (
            O => \N__24469\,
            I => \N__24463\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__24466\,
            I => \N__24460\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__24463\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__3562\ : Odrv12
    port map (
            O => \N__24460\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__3561\ : CascadeMux
    port map (
            O => \N__24455\,
            I => \N__24452\
        );

    \I__3560\ : InMux
    port map (
            O => \N__24452\,
            I => \N__24449\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__24449\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\
        );

    \I__3558\ : InMux
    port map (
            O => \N__24446\,
            I => \N__24443\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__24443\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\
        );

    \I__3556\ : InMux
    port map (
            O => \N__24440\,
            I => \N__24436\
        );

    \I__3555\ : InMux
    port map (
            O => \N__24439\,
            I => \N__24433\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__24436\,
            I => \N__24430\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__24433\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__3552\ : Odrv12
    port map (
            O => \N__24430\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__3551\ : CascadeMux
    port map (
            O => \N__24425\,
            I => \N__24422\
        );

    \I__3550\ : InMux
    port map (
            O => \N__24422\,
            I => \N__24419\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__24419\,
            I => \N__24416\
        );

    \I__3548\ : Odrv4
    port map (
            O => \N__24416\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\
        );

    \I__3547\ : InMux
    port map (
            O => \N__24413\,
            I => \bfn_8_7_0_\
        );

    \I__3546\ : InMux
    port map (
            O => \N__24410\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\
        );

    \I__3545\ : InMux
    port map (
            O => \N__24407\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\
        );

    \I__3544\ : InMux
    port map (
            O => \N__24404\,
            I => \N__24397\
        );

    \I__3543\ : InMux
    port map (
            O => \N__24403\,
            I => \N__24397\
        );

    \I__3542\ : InMux
    port map (
            O => \N__24402\,
            I => \N__24394\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__24397\,
            I => \N__24391\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__24394\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__3539\ : Odrv4
    port map (
            O => \N__24391\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__3538\ : InMux
    port map (
            O => \N__24386\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\
        );

    \I__3537\ : CascadeMux
    port map (
            O => \N__24383\,
            I => \N__24380\
        );

    \I__3536\ : InMux
    port map (
            O => \N__24380\,
            I => \N__24374\
        );

    \I__3535\ : InMux
    port map (
            O => \N__24379\,
            I => \N__24374\
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__24374\,
            I => \N__24370\
        );

    \I__3533\ : InMux
    port map (
            O => \N__24373\,
            I => \N__24367\
        );

    \I__3532\ : Span4Mux_h
    port map (
            O => \N__24370\,
            I => \N__24364\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__24367\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__3530\ : Odrv4
    port map (
            O => \N__24364\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__3529\ : InMux
    port map (
            O => \N__24359\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__3528\ : InMux
    port map (
            O => \N__24356\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\
        );

    \I__3527\ : InMux
    port map (
            O => \N__24353\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\
        );

    \I__3526\ : InMux
    port map (
            O => \N__24350\,
            I => \N__24347\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__24347\,
            I => \N__24342\
        );

    \I__3524\ : InMux
    port map (
            O => \N__24346\,
            I => \N__24339\
        );

    \I__3523\ : InMux
    port map (
            O => \N__24345\,
            I => \N__24336\
        );

    \I__3522\ : Span4Mux_v
    port map (
            O => \N__24342\,
            I => \N__24331\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__24339\,
            I => \N__24331\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__24336\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__3519\ : Odrv4
    port map (
            O => \N__24331\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__3518\ : InMux
    port map (
            O => \N__24326\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\
        );

    \I__3517\ : CascadeMux
    port map (
            O => \N__24323\,
            I => \N__24320\
        );

    \I__3516\ : InMux
    port map (
            O => \N__24320\,
            I => \N__24317\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__24317\,
            I => \N__24312\
        );

    \I__3514\ : InMux
    port map (
            O => \N__24316\,
            I => \N__24309\
        );

    \I__3513\ : InMux
    port map (
            O => \N__24315\,
            I => \N__24306\
        );

    \I__3512\ : Span4Mux_v
    port map (
            O => \N__24312\,
            I => \N__24303\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__24309\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__24306\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__3509\ : Odrv4
    port map (
            O => \N__24303\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__3508\ : InMux
    port map (
            O => \N__24296\,
            I => \bfn_8_8_0_\
        );

    \I__3507\ : InMux
    port map (
            O => \N__24293\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\
        );

    \I__3506\ : InMux
    port map (
            O => \N__24290\,
            I => \bfn_8_6_0_\
        );

    \I__3505\ : InMux
    port map (
            O => \N__24287\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\
        );

    \I__3504\ : InMux
    port map (
            O => \N__24284\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\
        );

    \I__3503\ : InMux
    port map (
            O => \N__24281\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\
        );

    \I__3502\ : InMux
    port map (
            O => \N__24278\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\
        );

    \I__3501\ : InMux
    port map (
            O => \N__24275\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\
        );

    \I__3500\ : InMux
    port map (
            O => \N__24272\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\
        );

    \I__3499\ : InMux
    port map (
            O => \N__24269\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\
        );

    \I__3498\ : InMux
    port map (
            O => \N__24266\,
            I => \N__24263\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__24263\,
            I => \N__24260\
        );

    \I__3496\ : Odrv12
    port map (
            O => \N__24260\,
            I => il_max_comp1_c
        );

    \I__3495\ : InMux
    port map (
            O => \N__24257\,
            I => \N__24254\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__24254\,
            I => \N__24251\
        );

    \I__3493\ : Span4Mux_h
    port map (
            O => \N__24251\,
            I => \N__24248\
        );

    \I__3492\ : Span4Mux_v
    port map (
            O => \N__24248\,
            I => \N__24245\
        );

    \I__3491\ : Odrv4
    port map (
            O => \N__24245\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\
        );

    \I__3490\ : InMux
    port map (
            O => \N__24242\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\
        );

    \I__3489\ : CascadeMux
    port map (
            O => \N__24239\,
            I => \N__24236\
        );

    \I__3488\ : InMux
    port map (
            O => \N__24236\,
            I => \N__24233\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__24233\,
            I => \N__24230\
        );

    \I__3486\ : Span4Mux_v
    port map (
            O => \N__24230\,
            I => \N__24227\
        );

    \I__3485\ : Odrv4
    port map (
            O => \N__24227\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3Z0Z_28\
        );

    \I__3484\ : InMux
    port map (
            O => \N__24224\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\
        );

    \I__3483\ : InMux
    port map (
            O => \N__24221\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\
        );

    \I__3482\ : InMux
    port map (
            O => \N__24218\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\
        );

    \I__3481\ : InMux
    port map (
            O => \N__24215\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\
        );

    \I__3480\ : InMux
    port map (
            O => \N__24212\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\
        );

    \I__3479\ : InMux
    port map (
            O => \N__24209\,
            I => \N__24206\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__24206\,
            I => \N__24203\
        );

    \I__3477\ : Span4Mux_h
    port map (
            O => \N__24203\,
            I => \N__24200\
        );

    \I__3476\ : Odrv4
    port map (
            O => \N__24200\,
            I => \pwm_generator_inst.un19_threshold_axb_3\
        );

    \I__3475\ : InMux
    port map (
            O => \N__24197\,
            I => \pwm_generator_inst.un19_threshold_cry_2\
        );

    \I__3474\ : InMux
    port map (
            O => \N__24194\,
            I => \N__24191\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__24191\,
            I => \N__24188\
        );

    \I__3472\ : Span4Mux_h
    port map (
            O => \N__24188\,
            I => \N__24185\
        );

    \I__3471\ : Odrv4
    port map (
            O => \N__24185\,
            I => \pwm_generator_inst.un19_threshold_axb_4\
        );

    \I__3470\ : InMux
    port map (
            O => \N__24182\,
            I => \pwm_generator_inst.un19_threshold_cry_3\
        );

    \I__3469\ : InMux
    port map (
            O => \N__24179\,
            I => \N__24176\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__24176\,
            I => \N__24173\
        );

    \I__3467\ : Span4Mux_v
    port map (
            O => \N__24173\,
            I => \N__24170\
        );

    \I__3466\ : Odrv4
    port map (
            O => \N__24170\,
            I => \pwm_generator_inst.un19_threshold_axb_5\
        );

    \I__3465\ : InMux
    port map (
            O => \N__24167\,
            I => \pwm_generator_inst.un19_threshold_cry_4\
        );

    \I__3464\ : InMux
    port map (
            O => \N__24164\,
            I => \N__24161\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__24161\,
            I => \N__24158\
        );

    \I__3462\ : Span4Mux_h
    port map (
            O => \N__24158\,
            I => \N__24155\
        );

    \I__3461\ : Odrv4
    port map (
            O => \N__24155\,
            I => \pwm_generator_inst.un19_threshold_axb_6\
        );

    \I__3460\ : InMux
    port map (
            O => \N__24152\,
            I => \pwm_generator_inst.un19_threshold_cry_5\
        );

    \I__3459\ : InMux
    port map (
            O => \N__24149\,
            I => \N__24146\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__24146\,
            I => \N__24143\
        );

    \I__3457\ : Span4Mux_h
    port map (
            O => \N__24143\,
            I => \N__24140\
        );

    \I__3456\ : Odrv4
    port map (
            O => \N__24140\,
            I => \pwm_generator_inst.un19_threshold_axb_7\
        );

    \I__3455\ : InMux
    port map (
            O => \N__24137\,
            I => \pwm_generator_inst.un19_threshold_cry_6\
        );

    \I__3454\ : InMux
    port map (
            O => \N__24134\,
            I => \bfn_7_24_0_\
        );

    \I__3453\ : InMux
    port map (
            O => \N__24131\,
            I => \N__24128\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__24128\,
            I => \N__24125\
        );

    \I__3451\ : Span4Mux_h
    port map (
            O => \N__24125\,
            I => \N__24122\
        );

    \I__3450\ : Odrv4
    port map (
            O => \N__24122\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\
        );

    \I__3449\ : InMux
    port map (
            O => \N__24119\,
            I => \N__24116\
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__24116\,
            I => \N__24113\
        );

    \I__3447\ : Span4Mux_v
    port map (
            O => \N__24113\,
            I => \N__24110\
        );

    \I__3446\ : Odrv4
    port map (
            O => \N__24110\,
            I => \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11\
        );

    \I__3445\ : InMux
    port map (
            O => \N__24107\,
            I => \pwm_generator_inst.un19_threshold_cry_8\
        );

    \I__3444\ : InMux
    port map (
            O => \N__24104\,
            I => \N__24101\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__24101\,
            I => \N__24096\
        );

    \I__3442\ : InMux
    port map (
            O => \N__24100\,
            I => \N__24093\
        );

    \I__3441\ : InMux
    port map (
            O => \N__24099\,
            I => \N__24090\
        );

    \I__3440\ : Span4Mux_h
    port map (
            O => \N__24096\,
            I => \N__24087\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__24093\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__24090\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__3437\ : Odrv4
    port map (
            O => \N__24087\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__3436\ : InMux
    port map (
            O => \N__24080\,
            I => \N__24076\
        );

    \I__3435\ : InMux
    port map (
            O => \N__24079\,
            I => \N__24073\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__24076\,
            I => \N__24070\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__24073\,
            I => \N__24067\
        );

    \I__3432\ : Span4Mux_h
    port map (
            O => \N__24070\,
            I => \N__24064\
        );

    \I__3431\ : Span4Mux_v
    port map (
            O => \N__24067\,
            I => \N__24061\
        );

    \I__3430\ : Odrv4
    port map (
            O => \N__24064\,
            I => \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\
        );

    \I__3429\ : Odrv4
    port map (
            O => \N__24061\,
            I => \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\
        );

    \I__3428\ : CascadeMux
    port map (
            O => \N__24056\,
            I => \N__24050\
        );

    \I__3427\ : CascadeMux
    port map (
            O => \N__24055\,
            I => \N__24047\
        );

    \I__3426\ : CascadeMux
    port map (
            O => \N__24054\,
            I => \N__24044\
        );

    \I__3425\ : InMux
    port map (
            O => \N__24053\,
            I => \N__24041\
        );

    \I__3424\ : InMux
    port map (
            O => \N__24050\,
            I => \N__24038\
        );

    \I__3423\ : InMux
    port map (
            O => \N__24047\,
            I => \N__24035\
        );

    \I__3422\ : InMux
    port map (
            O => \N__24044\,
            I => \N__24032\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__24041\,
            I => \N__24027\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__24038\,
            I => \N__24020\
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__24035\,
            I => \N__24020\
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__24032\,
            I => \N__24020\
        );

    \I__3417\ : InMux
    port map (
            O => \N__24031\,
            I => \N__24015\
        );

    \I__3416\ : CascadeMux
    port map (
            O => \N__24030\,
            I => \N__24012\
        );

    \I__3415\ : Span4Mux_v
    port map (
            O => \N__24027\,
            I => \N__24004\
        );

    \I__3414\ : Span4Mux_v
    port map (
            O => \N__24020\,
            I => \N__24004\
        );

    \I__3413\ : InMux
    port map (
            O => \N__24019\,
            I => \N__24001\
        );

    \I__3412\ : InMux
    port map (
            O => \N__24018\,
            I => \N__23998\
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__24015\,
            I => \N__23995\
        );

    \I__3410\ : InMux
    port map (
            O => \N__24012\,
            I => \N__23986\
        );

    \I__3409\ : InMux
    port map (
            O => \N__24011\,
            I => \N__23986\
        );

    \I__3408\ : InMux
    port map (
            O => \N__24010\,
            I => \N__23986\
        );

    \I__3407\ : InMux
    port map (
            O => \N__24009\,
            I => \N__23986\
        );

    \I__3406\ : Odrv4
    port map (
            O => \N__24004\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__24001\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__23998\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__3403\ : Odrv4
    port map (
            O => \N__23995\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__23986\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__3401\ : InMux
    port map (
            O => \N__23975\,
            I => \N__23972\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__23972\,
            I => \N__23969\
        );

    \I__3399\ : Span4Mux_v
    port map (
            O => \N__23969\,
            I => \N__23966\
        );

    \I__3398\ : Odrv4
    port map (
            O => \N__23966\,
            I => \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\
        );

    \I__3397\ : InMux
    port map (
            O => \N__23963\,
            I => \N__23960\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__23960\,
            I => \pwm_generator_inst.un19_threshold_axb_8\
        );

    \I__3395\ : InMux
    port map (
            O => \N__23957\,
            I => \N__23954\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__23954\,
            I => \N__23950\
        );

    \I__3393\ : InMux
    port map (
            O => \N__23953\,
            I => \N__23947\
        );

    \I__3392\ : Odrv12
    port map (
            O => \N__23950\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__23947\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\
        );

    \I__3390\ : CascadeMux
    port map (
            O => \N__23942\,
            I => \N__23937\
        );

    \I__3389\ : CascadeMux
    port map (
            O => \N__23941\,
            I => \N__23934\
        );

    \I__3388\ : CascadeMux
    port map (
            O => \N__23940\,
            I => \N__23931\
        );

    \I__3387\ : InMux
    port map (
            O => \N__23937\,
            I => \N__23924\
        );

    \I__3386\ : InMux
    port map (
            O => \N__23934\,
            I => \N__23924\
        );

    \I__3385\ : InMux
    port map (
            O => \N__23931\,
            I => \N__23924\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__23924\,
            I => \N__23921\
        );

    \I__3383\ : Odrv4
    port map (
            O => \N__23921\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_31\
        );

    \I__3382\ : InMux
    port map (
            O => \N__23918\,
            I => \N__23912\
        );

    \I__3381\ : InMux
    port map (
            O => \N__23917\,
            I => \N__23909\
        );

    \I__3380\ : InMux
    port map (
            O => \N__23916\,
            I => \N__23904\
        );

    \I__3379\ : InMux
    port map (
            O => \N__23915\,
            I => \N__23904\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__23912\,
            I => \N__23896\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__23909\,
            I => \N__23896\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__23904\,
            I => \N__23896\
        );

    \I__3375\ : InMux
    port map (
            O => \N__23903\,
            I => \N__23893\
        );

    \I__3374\ : Span4Mux_v
    port map (
            O => \N__23896\,
            I => \N__23890\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__23893\,
            I => \N__23887\
        );

    \I__3372\ : Span4Mux_v
    port map (
            O => \N__23890\,
            I => \N__23884\
        );

    \I__3371\ : Odrv12
    port map (
            O => \N__23887\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__3370\ : Odrv4
    port map (
            O => \N__23884\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__3369\ : InMux
    port map (
            O => \N__23879\,
            I => \N__23876\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__23876\,
            I => \N__23873\
        );

    \I__3367\ : Span4Mux_h
    port map (
            O => \N__23873\,
            I => \N__23870\
        );

    \I__3366\ : Odrv4
    port map (
            O => \N__23870\,
            I => \pwm_generator_inst.un19_threshold_axb_0\
        );

    \I__3365\ : InMux
    port map (
            O => \N__23867\,
            I => \N__23864\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__23864\,
            I => \N__23861\
        );

    \I__3363\ : Span4Mux_h
    port map (
            O => \N__23861\,
            I => \N__23858\
        );

    \I__3362\ : Odrv4
    port map (
            O => \N__23858\,
            I => \pwm_generator_inst.un19_threshold_axb_1\
        );

    \I__3361\ : InMux
    port map (
            O => \N__23855\,
            I => \pwm_generator_inst.un19_threshold_cry_0\
        );

    \I__3360\ : InMux
    port map (
            O => \N__23852\,
            I => \N__23849\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__23849\,
            I => \N__23846\
        );

    \I__3358\ : Span4Mux_h
    port map (
            O => \N__23846\,
            I => \N__23843\
        );

    \I__3357\ : Odrv4
    port map (
            O => \N__23843\,
            I => \pwm_generator_inst.un19_threshold_axb_2\
        );

    \I__3356\ : InMux
    port map (
            O => \N__23840\,
            I => \pwm_generator_inst.un19_threshold_cry_1\
        );

    \I__3355\ : InMux
    port map (
            O => \N__23837\,
            I => \N__23831\
        );

    \I__3354\ : InMux
    port map (
            O => \N__23836\,
            I => \N__23831\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__23831\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_21\
        );

    \I__3352\ : CascadeMux
    port map (
            O => \N__23828\,
            I => \phase_controller_inst1.stoper_hc.un4_running_df30_cascade_\
        );

    \I__3351\ : CascadeMux
    port map (
            O => \N__23825\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_\
        );

    \I__3350\ : CascadeMux
    port map (
            O => \N__23822\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5_cascade_\
        );

    \I__3349\ : InMux
    port map (
            O => \N__23819\,
            I => \N__23814\
        );

    \I__3348\ : InMux
    port map (
            O => \N__23818\,
            I => \N__23811\
        );

    \I__3347\ : InMux
    port map (
            O => \N__23817\,
            I => \N__23808\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__23814\,
            I => \pwm_generator_inst.un15_threshold_1_axb_13\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__23811\,
            I => \pwm_generator_inst.un15_threshold_1_axb_13\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__23808\,
            I => \pwm_generator_inst.un15_threshold_1_axb_13\
        );

    \I__3343\ : InMux
    port map (
            O => \N__23801\,
            I => \N__23798\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__23798\,
            I => \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\
        );

    \I__3341\ : InMux
    port map (
            O => \N__23795\,
            I => \pwm_generator_inst.un15_threshold_1_cry_12\
        );

    \I__3340\ : CascadeMux
    port map (
            O => \N__23792\,
            I => \N__23787\
        );

    \I__3339\ : InMux
    port map (
            O => \N__23791\,
            I => \N__23784\
        );

    \I__3338\ : InMux
    port map (
            O => \N__23790\,
            I => \N__23781\
        );

    \I__3337\ : InMux
    port map (
            O => \N__23787\,
            I => \N__23778\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__23784\,
            I => \N__23775\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__23781\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__23778\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__3333\ : Odrv4
    port map (
            O => \N__23775\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__3332\ : InMux
    port map (
            O => \N__23768\,
            I => \N__23765\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__23765\,
            I => \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\
        );

    \I__3330\ : InMux
    port map (
            O => \N__23762\,
            I => \pwm_generator_inst.un15_threshold_1_cry_13\
        );

    \I__3329\ : InMux
    port map (
            O => \N__23759\,
            I => \N__23754\
        );

    \I__3328\ : InMux
    port map (
            O => \N__23758\,
            I => \N__23751\
        );

    \I__3327\ : InMux
    port map (
            O => \N__23757\,
            I => \N__23748\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__23754\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__23751\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__23748\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__3323\ : InMux
    port map (
            O => \N__23741\,
            I => \N__23738\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__23738\,
            I => \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\
        );

    \I__3321\ : InMux
    port map (
            O => \N__23735\,
            I => \pwm_generator_inst.un15_threshold_1_cry_14\
        );

    \I__3320\ : InMux
    port map (
            O => \N__23732\,
            I => \N__23728\
        );

    \I__3319\ : InMux
    port map (
            O => \N__23731\,
            I => \N__23725\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__23728\,
            I => \pwm_generator_inst.un15_threshold_1_axb_16\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__23725\,
            I => \pwm_generator_inst.un15_threshold_1_axb_16\
        );

    \I__3316\ : InMux
    port map (
            O => \N__23720\,
            I => \N__23717\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__23717\,
            I => \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\
        );

    \I__3314\ : InMux
    port map (
            O => \N__23714\,
            I => \bfn_5_27_0_\
        );

    \I__3313\ : InMux
    port map (
            O => \N__23711\,
            I => \N__23706\
        );

    \I__3312\ : InMux
    port map (
            O => \N__23710\,
            I => \N__23703\
        );

    \I__3311\ : InMux
    port map (
            O => \N__23709\,
            I => \N__23700\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__23706\,
            I => \pwm_generator_inst.un15_threshold_1_axb_17\
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__23703\,
            I => \pwm_generator_inst.un15_threshold_1_axb_17\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__23700\,
            I => \pwm_generator_inst.un15_threshold_1_axb_17\
        );

    \I__3307\ : InMux
    port map (
            O => \N__23693\,
            I => \N__23690\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__23690\,
            I => \N__23687\
        );

    \I__3305\ : Odrv4
    port map (
            O => \N__23687\,
            I => \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\
        );

    \I__3304\ : InMux
    port map (
            O => \N__23684\,
            I => \pwm_generator_inst.un15_threshold_1_cry_16\
        );

    \I__3303\ : InMux
    port map (
            O => \N__23681\,
            I => \pwm_generator_inst.un15_threshold_1_cry_17\
        );

    \I__3302\ : InMux
    port map (
            O => \N__23678\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18\
        );

    \I__3301\ : InMux
    port map (
            O => \N__23675\,
            I => \N__23672\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__23672\,
            I => \N__23669\
        );

    \I__3299\ : Span4Mux_h
    port map (
            O => \N__23669\,
            I => \N__23666\
        );

    \I__3298\ : Span4Mux_h
    port map (
            O => \N__23666\,
            I => \N__23663\
        );

    \I__3297\ : Odrv4
    port map (
            O => \N__23663\,
            I => \pwm_generator_inst.O_5\
        );

    \I__3296\ : InMux
    port map (
            O => \N__23660\,
            I => \N__23657\
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__23657\,
            I => \pwm_generator_inst.un15_threshold_1_axb_5\
        );

    \I__3294\ : InMux
    port map (
            O => \N__23654\,
            I => \N__23651\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__23651\,
            I => \N__23648\
        );

    \I__3292\ : Span4Mux_h
    port map (
            O => \N__23648\,
            I => \N__23645\
        );

    \I__3291\ : Span4Mux_h
    port map (
            O => \N__23645\,
            I => \N__23642\
        );

    \I__3290\ : Odrv4
    port map (
            O => \N__23642\,
            I => \pwm_generator_inst.O_6\
        );

    \I__3289\ : InMux
    port map (
            O => \N__23639\,
            I => \N__23636\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__23636\,
            I => \pwm_generator_inst.un15_threshold_1_axb_6\
        );

    \I__3287\ : InMux
    port map (
            O => \N__23633\,
            I => \N__23630\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__23630\,
            I => \N__23627\
        );

    \I__3285\ : Span4Mux_v
    port map (
            O => \N__23627\,
            I => \N__23624\
        );

    \I__3284\ : Span4Mux_h
    port map (
            O => \N__23624\,
            I => \N__23621\
        );

    \I__3283\ : Odrv4
    port map (
            O => \N__23621\,
            I => \pwm_generator_inst.O_7\
        );

    \I__3282\ : InMux
    port map (
            O => \N__23618\,
            I => \N__23615\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__23615\,
            I => \pwm_generator_inst.un15_threshold_1_axb_7\
        );

    \I__3280\ : InMux
    port map (
            O => \N__23612\,
            I => \N__23609\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__23609\,
            I => \N__23606\
        );

    \I__3278\ : Span4Mux_h
    port map (
            O => \N__23606\,
            I => \N__23603\
        );

    \I__3277\ : Span4Mux_h
    port map (
            O => \N__23603\,
            I => \N__23600\
        );

    \I__3276\ : Odrv4
    port map (
            O => \N__23600\,
            I => \pwm_generator_inst.O_8\
        );

    \I__3275\ : InMux
    port map (
            O => \N__23597\,
            I => \N__23594\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__23594\,
            I => \pwm_generator_inst.un15_threshold_1_axb_8\
        );

    \I__3273\ : InMux
    port map (
            O => \N__23591\,
            I => \N__23588\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__23588\,
            I => \N__23585\
        );

    \I__3271\ : Span4Mux_h
    port map (
            O => \N__23585\,
            I => \N__23582\
        );

    \I__3270\ : Span4Mux_h
    port map (
            O => \N__23582\,
            I => \N__23579\
        );

    \I__3269\ : Odrv4
    port map (
            O => \N__23579\,
            I => \pwm_generator_inst.O_9\
        );

    \I__3268\ : InMux
    port map (
            O => \N__23576\,
            I => \N__23573\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__23573\,
            I => \pwm_generator_inst.un15_threshold_1_axb_9\
        );

    \I__3266\ : InMux
    port map (
            O => \N__23570\,
            I => \N__23566\
        );

    \I__3265\ : InMux
    port map (
            O => \N__23569\,
            I => \N__23562\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__23566\,
            I => \N__23559\
        );

    \I__3263\ : InMux
    port map (
            O => \N__23565\,
            I => \N__23556\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__23562\,
            I => \N__23553\
        );

    \I__3261\ : Span4Mux_h
    port map (
            O => \N__23559\,
            I => \N__23550\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__23556\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__3259\ : Odrv4
    port map (
            O => \N__23553\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__3258\ : Odrv4
    port map (
            O => \N__23550\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__3257\ : InMux
    port map (
            O => \N__23543\,
            I => \N__23540\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__23540\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\
        );

    \I__3255\ : InMux
    port map (
            O => \N__23537\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9\
        );

    \I__3254\ : InMux
    port map (
            O => \N__23534\,
            I => \N__23531\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__23531\,
            I => \N__23527\
        );

    \I__3252\ : InMux
    port map (
            O => \N__23530\,
            I => \N__23524\
        );

    \I__3251\ : Span12Mux_s6_v
    port map (
            O => \N__23527\,
            I => \N__23521\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__23524\,
            I => \N__23518\
        );

    \I__3249\ : Odrv12
    port map (
            O => \N__23521\,
            I => \pwm_generator_inst.un3_threshold\
        );

    \I__3248\ : Odrv4
    port map (
            O => \N__23518\,
            I => \pwm_generator_inst.un3_threshold\
        );

    \I__3247\ : InMux
    port map (
            O => \N__23513\,
            I => \pwm_generator_inst.un15_threshold_1_cry_10\
        );

    \I__3246\ : InMux
    port map (
            O => \N__23510\,
            I => \N__23506\
        );

    \I__3245\ : InMux
    port map (
            O => \N__23509\,
            I => \N__23502\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__23506\,
            I => \N__23499\
        );

    \I__3243\ : InMux
    port map (
            O => \N__23505\,
            I => \N__23496\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__23502\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__3241\ : Odrv4
    port map (
            O => \N__23499\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__23496\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__3239\ : InMux
    port map (
            O => \N__23489\,
            I => \N__23486\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__23486\,
            I => \N__23483\
        );

    \I__3237\ : Odrv4
    port map (
            O => \N__23483\,
            I => \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\
        );

    \I__3236\ : InMux
    port map (
            O => \N__23480\,
            I => \pwm_generator_inst.un15_threshold_1_cry_11\
        );

    \I__3235\ : InMux
    port map (
            O => \N__23477\,
            I => \N__23474\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__23474\,
            I => \N__23471\
        );

    \I__3233\ : Span4Mux_h
    port map (
            O => \N__23471\,
            I => \N__23468\
        );

    \I__3232\ : Sp12to4
    port map (
            O => \N__23468\,
            I => \N__23465\
        );

    \I__3231\ : Span12Mux_s5_v
    port map (
            O => \N__23465\,
            I => \N__23462\
        );

    \I__3230\ : Span12Mux_h
    port map (
            O => \N__23462\,
            I => \N__23459\
        );

    \I__3229\ : Odrv12
    port map (
            O => \N__23459\,
            I => \pwm_generator_inst.un2_threshold_2_1_16\
        );

    \I__3228\ : InMux
    port map (
            O => \N__23456\,
            I => \N__23453\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__23453\,
            I => \N__23450\
        );

    \I__3226\ : Span4Mux_h
    port map (
            O => \N__23450\,
            I => \N__23447\
        );

    \I__3225\ : Odrv4
    port map (
            O => \N__23447\,
            I => \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\
        );

    \I__3224\ : CascadeMux
    port map (
            O => \N__23444\,
            I => \N__23440\
        );

    \I__3223\ : InMux
    port map (
            O => \N__23443\,
            I => \N__23437\
        );

    \I__3222\ : InMux
    port map (
            O => \N__23440\,
            I => \N__23434\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__23437\,
            I => \N__23431\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__23434\,
            I => \N__23428\
        );

    \I__3219\ : Span4Mux_h
    port map (
            O => \N__23431\,
            I => \N__23425\
        );

    \I__3218\ : Odrv4
    port map (
            O => \N__23428\,
            I => \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\
        );

    \I__3217\ : Odrv4
    port map (
            O => \N__23425\,
            I => \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\
        );

    \I__3216\ : InMux
    port map (
            O => \N__23420\,
            I => \N__23416\
        );

    \I__3215\ : InMux
    port map (
            O => \N__23419\,
            I => \N__23413\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__23416\,
            I => \N__23410\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__23413\,
            I => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\
        );

    \I__3212\ : Odrv4
    port map (
            O => \N__23410\,
            I => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\
        );

    \I__3211\ : InMux
    port map (
            O => \N__23405\,
            I => \N__23402\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__23402\,
            I => \N__23399\
        );

    \I__3209\ : Span4Mux_h
    port map (
            O => \N__23399\,
            I => \N__23396\
        );

    \I__3208\ : Span4Mux_h
    port map (
            O => \N__23396\,
            I => \N__23393\
        );

    \I__3207\ : Odrv4
    port map (
            O => \N__23393\,
            I => \pwm_generator_inst.O_0\
        );

    \I__3206\ : InMux
    port map (
            O => \N__23390\,
            I => \N__23387\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__23387\,
            I => \pwm_generator_inst.un15_threshold_1_axb_0\
        );

    \I__3204\ : InMux
    port map (
            O => \N__23384\,
            I => \N__23381\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__23381\,
            I => \N__23378\
        );

    \I__3202\ : Span4Mux_h
    port map (
            O => \N__23378\,
            I => \N__23375\
        );

    \I__3201\ : Span4Mux_h
    port map (
            O => \N__23375\,
            I => \N__23372\
        );

    \I__3200\ : Odrv4
    port map (
            O => \N__23372\,
            I => \pwm_generator_inst.O_1\
        );

    \I__3199\ : InMux
    port map (
            O => \N__23369\,
            I => \N__23366\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__23366\,
            I => \pwm_generator_inst.un15_threshold_1_axb_1\
        );

    \I__3197\ : InMux
    port map (
            O => \N__23363\,
            I => \N__23360\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__23360\,
            I => \N__23357\
        );

    \I__3195\ : Span12Mux_h
    port map (
            O => \N__23357\,
            I => \N__23354\
        );

    \I__3194\ : Odrv12
    port map (
            O => \N__23354\,
            I => \pwm_generator_inst.O_2\
        );

    \I__3193\ : InMux
    port map (
            O => \N__23351\,
            I => \N__23348\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__23348\,
            I => \pwm_generator_inst.un15_threshold_1_axb_2\
        );

    \I__3191\ : InMux
    port map (
            O => \N__23345\,
            I => \N__23342\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__23342\,
            I => \N__23339\
        );

    \I__3189\ : Span12Mux_s7_v
    port map (
            O => \N__23339\,
            I => \N__23336\
        );

    \I__3188\ : Odrv12
    port map (
            O => \N__23336\,
            I => \pwm_generator_inst.O_3\
        );

    \I__3187\ : InMux
    port map (
            O => \N__23333\,
            I => \N__23330\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__23330\,
            I => \pwm_generator_inst.un15_threshold_1_axb_3\
        );

    \I__3185\ : InMux
    port map (
            O => \N__23327\,
            I => \N__23324\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__23324\,
            I => \N__23321\
        );

    \I__3183\ : Span4Mux_h
    port map (
            O => \N__23321\,
            I => \N__23318\
        );

    \I__3182\ : Span4Mux_h
    port map (
            O => \N__23318\,
            I => \N__23315\
        );

    \I__3181\ : Odrv4
    port map (
            O => \N__23315\,
            I => \pwm_generator_inst.O_4\
        );

    \I__3180\ : InMux
    port map (
            O => \N__23312\,
            I => \N__23309\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__23309\,
            I => \pwm_generator_inst.un15_threshold_1_axb_4\
        );

    \I__3178\ : CascadeMux
    port map (
            O => \N__23306\,
            I => \N__23303\
        );

    \I__3177\ : InMux
    port map (
            O => \N__23303\,
            I => \N__23300\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__23300\,
            I => \N__23297\
        );

    \I__3175\ : Odrv4
    port map (
            O => \N__23297\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\
        );

    \I__3174\ : CascadeMux
    port map (
            O => \N__23294\,
            I => \N__23291\
        );

    \I__3173\ : InMux
    port map (
            O => \N__23291\,
            I => \N__23288\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__23288\,
            I => \N__23284\
        );

    \I__3171\ : InMux
    port map (
            O => \N__23287\,
            I => \N__23279\
        );

    \I__3170\ : Span4Mux_v
    port map (
            O => \N__23284\,
            I => \N__23276\
        );

    \I__3169\ : InMux
    port map (
            O => \N__23283\,
            I => \N__23271\
        );

    \I__3168\ : InMux
    port map (
            O => \N__23282\,
            I => \N__23271\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__23279\,
            I => \N__23268\
        );

    \I__3166\ : Odrv4
    port map (
            O => \N__23276\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__23271\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__3164\ : Odrv12
    port map (
            O => \N__23268\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__3163\ : InMux
    port map (
            O => \N__23261\,
            I => \N__23249\
        );

    \I__3162\ : InMux
    port map (
            O => \N__23260\,
            I => \N__23246\
        );

    \I__3161\ : CascadeMux
    port map (
            O => \N__23259\,
            I => \N__23242\
        );

    \I__3160\ : CascadeMux
    port map (
            O => \N__23258\,
            I => \N__23239\
        );

    \I__3159\ : CascadeMux
    port map (
            O => \N__23257\,
            I => \N__23236\
        );

    \I__3158\ : InMux
    port map (
            O => \N__23256\,
            I => \N__23224\
        );

    \I__3157\ : InMux
    port map (
            O => \N__23255\,
            I => \N__23217\
        );

    \I__3156\ : InMux
    port map (
            O => \N__23254\,
            I => \N__23217\
        );

    \I__3155\ : InMux
    port map (
            O => \N__23253\,
            I => \N__23212\
        );

    \I__3154\ : InMux
    port map (
            O => \N__23252\,
            I => \N__23212\
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__23249\,
            I => \N__23207\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__23246\,
            I => \N__23207\
        );

    \I__3151\ : InMux
    port map (
            O => \N__23245\,
            I => \N__23204\
        );

    \I__3150\ : InMux
    port map (
            O => \N__23242\,
            I => \N__23193\
        );

    \I__3149\ : InMux
    port map (
            O => \N__23239\,
            I => \N__23193\
        );

    \I__3148\ : InMux
    port map (
            O => \N__23236\,
            I => \N__23193\
        );

    \I__3147\ : InMux
    port map (
            O => \N__23235\,
            I => \N__23193\
        );

    \I__3146\ : InMux
    port map (
            O => \N__23234\,
            I => \N__23193\
        );

    \I__3145\ : InMux
    port map (
            O => \N__23233\,
            I => \N__23190\
        );

    \I__3144\ : InMux
    port map (
            O => \N__23232\,
            I => \N__23168\
        );

    \I__3143\ : InMux
    port map (
            O => \N__23231\,
            I => \N__23168\
        );

    \I__3142\ : InMux
    port map (
            O => \N__23230\,
            I => \N__23168\
        );

    \I__3141\ : InMux
    port map (
            O => \N__23229\,
            I => \N__23168\
        );

    \I__3140\ : InMux
    port map (
            O => \N__23228\,
            I => \N__23168\
        );

    \I__3139\ : InMux
    port map (
            O => \N__23227\,
            I => \N__23168\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__23224\,
            I => \N__23165\
        );

    \I__3137\ : InMux
    port map (
            O => \N__23223\,
            I => \N__23160\
        );

    \I__3136\ : InMux
    port map (
            O => \N__23222\,
            I => \N__23160\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__23217\,
            I => \N__23156\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__23212\,
            I => \N__23149\
        );

    \I__3133\ : Span4Mux_h
    port map (
            O => \N__23207\,
            I => \N__23149\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__23204\,
            I => \N__23149\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__23193\,
            I => \N__23144\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__23190\,
            I => \N__23144\
        );

    \I__3129\ : InMux
    port map (
            O => \N__23189\,
            I => \N__23141\
        );

    \I__3128\ : InMux
    port map (
            O => \N__23188\,
            I => \N__23128\
        );

    \I__3127\ : InMux
    port map (
            O => \N__23187\,
            I => \N__23128\
        );

    \I__3126\ : InMux
    port map (
            O => \N__23186\,
            I => \N__23128\
        );

    \I__3125\ : InMux
    port map (
            O => \N__23185\,
            I => \N__23128\
        );

    \I__3124\ : InMux
    port map (
            O => \N__23184\,
            I => \N__23128\
        );

    \I__3123\ : InMux
    port map (
            O => \N__23183\,
            I => \N__23128\
        );

    \I__3122\ : InMux
    port map (
            O => \N__23182\,
            I => \N__23123\
        );

    \I__3121\ : InMux
    port map (
            O => \N__23181\,
            I => \N__23123\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__23168\,
            I => \N__23120\
        );

    \I__3119\ : Span4Mux_v
    port map (
            O => \N__23165\,
            I => \N__23117\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__23160\,
            I => \N__23114\
        );

    \I__3117\ : InMux
    port map (
            O => \N__23159\,
            I => \N__23111\
        );

    \I__3116\ : Span4Mux_v
    port map (
            O => \N__23156\,
            I => \N__23106\
        );

    \I__3115\ : Span4Mux_v
    port map (
            O => \N__23149\,
            I => \N__23106\
        );

    \I__3114\ : Span4Mux_h
    port map (
            O => \N__23144\,
            I => \N__23103\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__23141\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__23128\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__23123\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3110\ : Odrv4
    port map (
            O => \N__23120\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3109\ : Odrv4
    port map (
            O => \N__23117\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3108\ : Odrv12
    port map (
            O => \N__23114\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__23111\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3106\ : Odrv4
    port map (
            O => \N__23106\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3105\ : Odrv4
    port map (
            O => \N__23103\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3104\ : CascadeMux
    port map (
            O => \N__23084\,
            I => \N__23078\
        );

    \I__3103\ : InMux
    port map (
            O => \N__23083\,
            I => \N__23068\
        );

    \I__3102\ : InMux
    port map (
            O => \N__23082\,
            I => \N__23068\
        );

    \I__3101\ : InMux
    port map (
            O => \N__23081\,
            I => \N__23065\
        );

    \I__3100\ : InMux
    port map (
            O => \N__23078\,
            I => \N__23058\
        );

    \I__3099\ : InMux
    port map (
            O => \N__23077\,
            I => \N__23058\
        );

    \I__3098\ : InMux
    port map (
            O => \N__23076\,
            I => \N__23055\
        );

    \I__3097\ : InMux
    port map (
            O => \N__23075\,
            I => \N__23030\
        );

    \I__3096\ : InMux
    port map (
            O => \N__23074\,
            I => \N__23030\
        );

    \I__3095\ : InMux
    port map (
            O => \N__23073\,
            I => \N__23027\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__23068\,
            I => \N__23024\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__23065\,
            I => \N__23021\
        );

    \I__3092\ : InMux
    port map (
            O => \N__23064\,
            I => \N__23016\
        );

    \I__3091\ : InMux
    port map (
            O => \N__23063\,
            I => \N__23016\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__23058\,
            I => \N__23011\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__23055\,
            I => \N__23011\
        );

    \I__3088\ : InMux
    port map (
            O => \N__23054\,
            I => \N__23002\
        );

    \I__3087\ : InMux
    port map (
            O => \N__23053\,
            I => \N__23002\
        );

    \I__3086\ : InMux
    port map (
            O => \N__23052\,
            I => \N__23002\
        );

    \I__3085\ : InMux
    port map (
            O => \N__23051\,
            I => \N__23002\
        );

    \I__3084\ : InMux
    port map (
            O => \N__23050\,
            I => \N__22997\
        );

    \I__3083\ : InMux
    port map (
            O => \N__23049\,
            I => \N__22997\
        );

    \I__3082\ : InMux
    port map (
            O => \N__23048\,
            I => \N__22990\
        );

    \I__3081\ : InMux
    port map (
            O => \N__23047\,
            I => \N__22990\
        );

    \I__3080\ : InMux
    port map (
            O => \N__23046\,
            I => \N__22990\
        );

    \I__3079\ : InMux
    port map (
            O => \N__23045\,
            I => \N__22977\
        );

    \I__3078\ : InMux
    port map (
            O => \N__23044\,
            I => \N__22977\
        );

    \I__3077\ : InMux
    port map (
            O => \N__23043\,
            I => \N__22977\
        );

    \I__3076\ : InMux
    port map (
            O => \N__23042\,
            I => \N__22977\
        );

    \I__3075\ : InMux
    port map (
            O => \N__23041\,
            I => \N__22977\
        );

    \I__3074\ : InMux
    port map (
            O => \N__23040\,
            I => \N__22977\
        );

    \I__3073\ : InMux
    port map (
            O => \N__23039\,
            I => \N__22966\
        );

    \I__3072\ : InMux
    port map (
            O => \N__23038\,
            I => \N__22966\
        );

    \I__3071\ : InMux
    port map (
            O => \N__23037\,
            I => \N__22966\
        );

    \I__3070\ : InMux
    port map (
            O => \N__23036\,
            I => \N__22966\
        );

    \I__3069\ : InMux
    port map (
            O => \N__23035\,
            I => \N__22966\
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__23030\,
            I => \N__22963\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__23027\,
            I => \N__22960\
        );

    \I__3066\ : Span4Mux_v
    port map (
            O => \N__23024\,
            I => \N__22955\
        );

    \I__3065\ : Span4Mux_v
    port map (
            O => \N__23021\,
            I => \N__22955\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__23016\,
            I => \N__22950\
        );

    \I__3063\ : Span4Mux_v
    port map (
            O => \N__23011\,
            I => \N__22950\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__23002\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__22997\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__22990\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__22977\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__22966\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__3057\ : Odrv4
    port map (
            O => \N__22963\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__3056\ : Odrv12
    port map (
            O => \N__22960\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__3055\ : Odrv4
    port map (
            O => \N__22955\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__3054\ : Odrv4
    port map (
            O => \N__22950\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__3053\ : CascadeMux
    port map (
            O => \N__22931\,
            I => \N__22928\
        );

    \I__3052\ : InMux
    port map (
            O => \N__22928\,
            I => \N__22925\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__22925\,
            I => \N__22922\
        );

    \I__3050\ : Span4Mux_h
    port map (
            O => \N__22922\,
            I => \N__22919\
        );

    \I__3049\ : Odrv4
    port map (
            O => \N__22919\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\
        );

    \I__3048\ : CascadeMux
    port map (
            O => \N__22916\,
            I => \N__22913\
        );

    \I__3047\ : InMux
    port map (
            O => \N__22913\,
            I => \N__22909\
        );

    \I__3046\ : InMux
    port map (
            O => \N__22912\,
            I => \N__22905\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__22909\,
            I => \N__22901\
        );

    \I__3044\ : CascadeMux
    port map (
            O => \N__22908\,
            I => \N__22898\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__22905\,
            I => \N__22895\
        );

    \I__3042\ : InMux
    port map (
            O => \N__22904\,
            I => \N__22892\
        );

    \I__3041\ : Span4Mux_h
    port map (
            O => \N__22901\,
            I => \N__22889\
        );

    \I__3040\ : InMux
    port map (
            O => \N__22898\,
            I => \N__22886\
        );

    \I__3039\ : Span4Mux_h
    port map (
            O => \N__22895\,
            I => \N__22883\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__22892\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__3037\ : Odrv4
    port map (
            O => \N__22889\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__22886\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__3035\ : Odrv4
    port map (
            O => \N__22883\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__3034\ : CascadeMux
    port map (
            O => \N__22874\,
            I => \N__22870\
        );

    \I__3033\ : InMux
    port map (
            O => \N__22873\,
            I => \N__22866\
        );

    \I__3032\ : InMux
    port map (
            O => \N__22870\,
            I => \N__22863\
        );

    \I__3031\ : InMux
    port map (
            O => \N__22869\,
            I => \N__22859\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__22866\,
            I => \N__22854\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__22863\,
            I => \N__22854\
        );

    \I__3028\ : InMux
    port map (
            O => \N__22862\,
            I => \N__22851\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__22859\,
            I => \N__22848\
        );

    \I__3026\ : Span4Mux_v
    port map (
            O => \N__22854\,
            I => \N__22843\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__22851\,
            I => \N__22843\
        );

    \I__3024\ : Span4Mux_v
    port map (
            O => \N__22848\,
            I => \N__22840\
        );

    \I__3023\ : Span4Mux_h
    port map (
            O => \N__22843\,
            I => \N__22837\
        );

    \I__3022\ : Odrv4
    port map (
            O => \N__22840\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__3021\ : Odrv4
    port map (
            O => \N__22837\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__3020\ : InMux
    port map (
            O => \N__22832\,
            I => \N__22827\
        );

    \I__3019\ : InMux
    port map (
            O => \N__22831\,
            I => \N__22824\
        );

    \I__3018\ : InMux
    port map (
            O => \N__22830\,
            I => \N__22821\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__22827\,
            I => \N__22817\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__22824\,
            I => \N__22814\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__22821\,
            I => \N__22811\
        );

    \I__3014\ : InMux
    port map (
            O => \N__22820\,
            I => \N__22808\
        );

    \I__3013\ : Span4Mux_h
    port map (
            O => \N__22817\,
            I => \N__22805\
        );

    \I__3012\ : Span4Mux_v
    port map (
            O => \N__22814\,
            I => \N__22800\
        );

    \I__3011\ : Span4Mux_h
    port map (
            O => \N__22811\,
            I => \N__22800\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__22808\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__3009\ : Odrv4
    port map (
            O => \N__22805\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__3008\ : Odrv4
    port map (
            O => \N__22800\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__3007\ : CascadeMux
    port map (
            O => \N__22793\,
            I => \N__22788\
        );

    \I__3006\ : CascadeMux
    port map (
            O => \N__22792\,
            I => \N__22785\
        );

    \I__3005\ : InMux
    port map (
            O => \N__22791\,
            I => \N__22782\
        );

    \I__3004\ : InMux
    port map (
            O => \N__22788\,
            I => \N__22779\
        );

    \I__3003\ : InMux
    port map (
            O => \N__22785\,
            I => \N__22776\
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__22782\,
            I => \N__22773\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__22779\,
            I => \N__22770\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__22776\,
            I => \N__22767\
        );

    \I__2999\ : Span4Mux_h
    port map (
            O => \N__22773\,
            I => \N__22763\
        );

    \I__2998\ : Span4Mux_h
    port map (
            O => \N__22770\,
            I => \N__22758\
        );

    \I__2997\ : Span4Mux_v
    port map (
            O => \N__22767\,
            I => \N__22758\
        );

    \I__2996\ : InMux
    port map (
            O => \N__22766\,
            I => \N__22755\
        );

    \I__2995\ : Odrv4
    port map (
            O => \N__22763\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__2994\ : Odrv4
    port map (
            O => \N__22758\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__22755\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__2992\ : InMux
    port map (
            O => \N__22748\,
            I => \N__22745\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__22745\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3\
        );

    \I__2990\ : CascadeMux
    port map (
            O => \N__22742\,
            I => \N__22739\
        );

    \I__2989\ : InMux
    port map (
            O => \N__22739\,
            I => \N__22736\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__22736\,
            I => \N__22733\
        );

    \I__2987\ : Span4Mux_h
    port map (
            O => \N__22733\,
            I => \N__22728\
        );

    \I__2986\ : InMux
    port map (
            O => \N__22732\,
            I => \N__22724\
        );

    \I__2985\ : InMux
    port map (
            O => \N__22731\,
            I => \N__22721\
        );

    \I__2984\ : Span4Mux_v
    port map (
            O => \N__22728\,
            I => \N__22718\
        );

    \I__2983\ : InMux
    port map (
            O => \N__22727\,
            I => \N__22715\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__22724\,
            I => \N__22710\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__22721\,
            I => \N__22710\
        );

    \I__2980\ : Odrv4
    port map (
            O => \N__22718\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__22715\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__2978\ : Odrv12
    port map (
            O => \N__22710\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__2977\ : CascadeMux
    port map (
            O => \N__22703\,
            I => \N__22700\
        );

    \I__2976\ : InMux
    port map (
            O => \N__22700\,
            I => \N__22696\
        );

    \I__2975\ : InMux
    port map (
            O => \N__22699\,
            I => \N__22691\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__22696\,
            I => \N__22688\
        );

    \I__2973\ : InMux
    port map (
            O => \N__22695\,
            I => \N__22685\
        );

    \I__2972\ : InMux
    port map (
            O => \N__22694\,
            I => \N__22682\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__22691\,
            I => \N__22679\
        );

    \I__2970\ : Odrv12
    port map (
            O => \N__22688\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__22685\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__22682\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__2967\ : Odrv4
    port map (
            O => \N__22679\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__2966\ : CascadeMux
    port map (
            O => \N__22670\,
            I => \current_shift_inst.PI_CTRL.N_44_cascade_\
        );

    \I__2965\ : InMux
    port map (
            O => \N__22667\,
            I => \N__22664\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__22664\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\
        );

    \I__2963\ : InMux
    port map (
            O => \N__22661\,
            I => \N__22658\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__22658\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\
        );

    \I__2961\ : InMux
    port map (
            O => \N__22655\,
            I => \N__22652\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__22652\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\
        );

    \I__2959\ : CascadeMux
    port map (
            O => \N__22649\,
            I => \N__22646\
        );

    \I__2958\ : InMux
    port map (
            O => \N__22646\,
            I => \N__22643\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__22643\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\
        );

    \I__2956\ : InMux
    port map (
            O => \N__22640\,
            I => \N__22637\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__22637\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\
        );

    \I__2954\ : CascadeMux
    port map (
            O => \N__22634\,
            I => \N__22621\
        );

    \I__2953\ : CascadeMux
    port map (
            O => \N__22633\,
            I => \N__22618\
        );

    \I__2952\ : CascadeMux
    port map (
            O => \N__22632\,
            I => \N__22603\
        );

    \I__2951\ : CascadeMux
    port map (
            O => \N__22631\,
            I => \N__22599\
        );

    \I__2950\ : InMux
    port map (
            O => \N__22630\,
            I => \N__22582\
        );

    \I__2949\ : InMux
    port map (
            O => \N__22629\,
            I => \N__22582\
        );

    \I__2948\ : InMux
    port map (
            O => \N__22628\,
            I => \N__22582\
        );

    \I__2947\ : InMux
    port map (
            O => \N__22627\,
            I => \N__22582\
        );

    \I__2946\ : InMux
    port map (
            O => \N__22626\,
            I => \N__22582\
        );

    \I__2945\ : InMux
    port map (
            O => \N__22625\,
            I => \N__22582\
        );

    \I__2944\ : InMux
    port map (
            O => \N__22624\,
            I => \N__22582\
        );

    \I__2943\ : InMux
    port map (
            O => \N__22621\,
            I => \N__22577\
        );

    \I__2942\ : InMux
    port map (
            O => \N__22618\,
            I => \N__22577\
        );

    \I__2941\ : InMux
    port map (
            O => \N__22617\,
            I => \N__22566\
        );

    \I__2940\ : InMux
    port map (
            O => \N__22616\,
            I => \N__22566\
        );

    \I__2939\ : InMux
    port map (
            O => \N__22615\,
            I => \N__22566\
        );

    \I__2938\ : InMux
    port map (
            O => \N__22614\,
            I => \N__22566\
        );

    \I__2937\ : InMux
    port map (
            O => \N__22613\,
            I => \N__22566\
        );

    \I__2936\ : InMux
    port map (
            O => \N__22612\,
            I => \N__22561\
        );

    \I__2935\ : InMux
    port map (
            O => \N__22611\,
            I => \N__22556\
        );

    \I__2934\ : InMux
    port map (
            O => \N__22610\,
            I => \N__22556\
        );

    \I__2933\ : InMux
    port map (
            O => \N__22609\,
            I => \N__22553\
        );

    \I__2932\ : CascadeMux
    port map (
            O => \N__22608\,
            I => \N__22548\
        );

    \I__2931\ : CascadeMux
    port map (
            O => \N__22607\,
            I => \N__22545\
        );

    \I__2930\ : CascadeMux
    port map (
            O => \N__22606\,
            I => \N__22542\
        );

    \I__2929\ : InMux
    port map (
            O => \N__22603\,
            I => \N__22538\
        );

    \I__2928\ : InMux
    port map (
            O => \N__22602\,
            I => \N__22533\
        );

    \I__2927\ : InMux
    port map (
            O => \N__22599\,
            I => \N__22533\
        );

    \I__2926\ : InMux
    port map (
            O => \N__22598\,
            I => \N__22528\
        );

    \I__2925\ : InMux
    port map (
            O => \N__22597\,
            I => \N__22528\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__22582\,
            I => \N__22525\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__22577\,
            I => \N__22520\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__22566\,
            I => \N__22520\
        );

    \I__2921\ : InMux
    port map (
            O => \N__22565\,
            I => \N__22515\
        );

    \I__2920\ : InMux
    port map (
            O => \N__22564\,
            I => \N__22515\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__22561\,
            I => \N__22510\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__22556\,
            I => \N__22510\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__22553\,
            I => \N__22507\
        );

    \I__2916\ : InMux
    port map (
            O => \N__22552\,
            I => \N__22494\
        );

    \I__2915\ : InMux
    port map (
            O => \N__22551\,
            I => \N__22494\
        );

    \I__2914\ : InMux
    port map (
            O => \N__22548\,
            I => \N__22494\
        );

    \I__2913\ : InMux
    port map (
            O => \N__22545\,
            I => \N__22494\
        );

    \I__2912\ : InMux
    port map (
            O => \N__22542\,
            I => \N__22494\
        );

    \I__2911\ : InMux
    port map (
            O => \N__22541\,
            I => \N__22494\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__22538\,
            I => \N__22491\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__22533\,
            I => \N__22488\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__22528\,
            I => \N__22485\
        );

    \I__2907\ : Span4Mux_h
    port map (
            O => \N__22525\,
            I => \N__22482\
        );

    \I__2906\ : Span4Mux_h
    port map (
            O => \N__22520\,
            I => \N__22479\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__22515\,
            I => \N__22472\
        );

    \I__2904\ : Span4Mux_v
    port map (
            O => \N__22510\,
            I => \N__22472\
        );

    \I__2903\ : Span4Mux_h
    port map (
            O => \N__22507\,
            I => \N__22472\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__22494\,
            I => \N__22465\
        );

    \I__2901\ : Span12Mux_v
    port map (
            O => \N__22491\,
            I => \N__22465\
        );

    \I__2900\ : Span12Mux_v
    port map (
            O => \N__22488\,
            I => \N__22465\
        );

    \I__2899\ : Odrv12
    port map (
            O => \N__22485\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__2898\ : Odrv4
    port map (
            O => \N__22482\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__2897\ : Odrv4
    port map (
            O => \N__22479\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__2896\ : Odrv4
    port map (
            O => \N__22472\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__2895\ : Odrv12
    port map (
            O => \N__22465\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__2894\ : InMux
    port map (
            O => \N__22454\,
            I => \N__22451\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__22451\,
            I => \N__22448\
        );

    \I__2892\ : Odrv12
    port map (
            O => \N__22448\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\
        );

    \I__2891\ : InMux
    port map (
            O => \N__22445\,
            I => \N__22442\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__22442\,
            I => \N__22439\
        );

    \I__2889\ : Odrv4
    port map (
            O => \N__22439\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\
        );

    \I__2888\ : InMux
    port map (
            O => \N__22436\,
            I => \N__22430\
        );

    \I__2887\ : InMux
    port map (
            O => \N__22435\,
            I => \N__22430\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__22430\,
            I => \N__22427\
        );

    \I__2885\ : Odrv4
    port map (
            O => \N__22427\,
            I => \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\
        );

    \I__2884\ : CascadeMux
    port map (
            O => \N__22424\,
            I => \pwm_generator_inst.un15_threshold_1_axb_16_cascade_\
        );

    \I__2883\ : InMux
    port map (
            O => \N__22421\,
            I => \N__22417\
        );

    \I__2882\ : InMux
    port map (
            O => \N__22420\,
            I => \N__22414\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__22417\,
            I => \N__22411\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__22414\,
            I => \N__22408\
        );

    \I__2879\ : Span4Mux_v
    port map (
            O => \N__22411\,
            I => \N__22405\
        );

    \I__2878\ : Odrv4
    port map (
            O => \N__22408\,
            I => \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\
        );

    \I__2877\ : Odrv4
    port map (
            O => \N__22405\,
            I => \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\
        );

    \I__2876\ : InMux
    port map (
            O => \N__22400\,
            I => \N__22396\
        );

    \I__2875\ : InMux
    port map (
            O => \N__22399\,
            I => \N__22393\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__22396\,
            I => \N__22390\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__22393\,
            I => \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\
        );

    \I__2872\ : Odrv4
    port map (
            O => \N__22390\,
            I => \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\
        );

    \I__2871\ : CascadeMux
    port map (
            O => \N__22385\,
            I => \N__22381\
        );

    \I__2870\ : InMux
    port map (
            O => \N__22384\,
            I => \N__22378\
        );

    \I__2869\ : InMux
    port map (
            O => \N__22381\,
            I => \N__22375\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__22378\,
            I => \N__22372\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__22375\,
            I => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\
        );

    \I__2866\ : Odrv4
    port map (
            O => \N__22372\,
            I => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\
        );

    \I__2865\ : CascadeMux
    port map (
            O => \N__22367\,
            I => \N__22364\
        );

    \I__2864\ : InMux
    port map (
            O => \N__22364\,
            I => \N__22360\
        );

    \I__2863\ : InMux
    port map (
            O => \N__22363\,
            I => \N__22357\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__22360\,
            I => \phase_controller_inst1.stoper_hc.runningZ0\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__22357\,
            I => \phase_controller_inst1.stoper_hc.runningZ0\
        );

    \I__2860\ : CascadeMux
    port map (
            O => \N__22352\,
            I => \N__22349\
        );

    \I__2859\ : InMux
    port map (
            O => \N__22349\,
            I => \N__22346\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__22346\,
            I => \N__22343\
        );

    \I__2857\ : Span12Mux_h
    port map (
            O => \N__22343\,
            I => \N__22340\
        );

    \I__2856\ : Odrv12
    port map (
            O => \N__22340\,
            I => \pwm_generator_inst.un2_threshold_2_14\
        );

    \I__2855\ : InMux
    port map (
            O => \N__22337\,
            I => \N__22334\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__22334\,
            I => \N__22331\
        );

    \I__2853\ : Odrv4
    port map (
            O => \N__22331\,
            I => \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0\
        );

    \I__2852\ : InMux
    port map (
            O => \N__22328\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_13\
        );

    \I__2851\ : CascadeMux
    port map (
            O => \N__22325\,
            I => \N__22322\
        );

    \I__2850\ : InMux
    port map (
            O => \N__22322\,
            I => \N__22319\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__22319\,
            I => \N__22316\
        );

    \I__2848\ : Odrv4
    port map (
            O => \N__22316\,
            I => \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0\
        );

    \I__2847\ : InMux
    port map (
            O => \N__22313\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_14\
        );

    \I__2846\ : InMux
    port map (
            O => \N__22310\,
            I => \N__22307\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__22307\,
            I => \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\
        );

    \I__2844\ : InMux
    port map (
            O => \N__22304\,
            I => \bfn_4_25_0_\
        );

    \I__2843\ : CascadeMux
    port map (
            O => \N__22301\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81_cascade_\
        );

    \I__2842\ : CascadeMux
    port map (
            O => \N__22298\,
            I => \N__22295\
        );

    \I__2841\ : InMux
    port map (
            O => \N__22295\,
            I => \N__22292\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__22292\,
            I => \N__22288\
        );

    \I__2839\ : InMux
    port map (
            O => \N__22291\,
            I => \N__22285\
        );

    \I__2838\ : Span4Mux_v
    port map (
            O => \N__22288\,
            I => \N__22280\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__22285\,
            I => \N__22280\
        );

    \I__2836\ : Span4Mux_h
    port map (
            O => \N__22280\,
            I => \N__22277\
        );

    \I__2835\ : Odrv4
    port map (
            O => \N__22277\,
            I => \pwm_generator_inst.O_10\
        );

    \I__2834\ : InMux
    port map (
            O => \N__22274\,
            I => \N__22271\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__22271\,
            I => \N__22268\
        );

    \I__2832\ : Span4Mux_h
    port map (
            O => \N__22268\,
            I => \N__22265\
        );

    \I__2831\ : Odrv4
    port map (
            O => \N__22265\,
            I => \pwm_generator_inst.un2_threshold_1_22\
        );

    \I__2830\ : CascadeMux
    port map (
            O => \N__22262\,
            I => \N__22259\
        );

    \I__2829\ : InMux
    port map (
            O => \N__22259\,
            I => \N__22256\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__22256\,
            I => \N__22253\
        );

    \I__2827\ : Span12Mux_h
    port map (
            O => \N__22253\,
            I => \N__22250\
        );

    \I__2826\ : Odrv12
    port map (
            O => \N__22250\,
            I => \pwm_generator_inst.un2_threshold_2_7\
        );

    \I__2825\ : CascadeMux
    port map (
            O => \N__22247\,
            I => \N__22244\
        );

    \I__2824\ : InMux
    port map (
            O => \N__22244\,
            I => \N__22241\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__22241\,
            I => \N__22238\
        );

    \I__2822\ : Odrv4
    port map (
            O => \N__22238\,
            I => \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0\
        );

    \I__2821\ : InMux
    port map (
            O => \N__22235\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_6\
        );

    \I__2820\ : InMux
    port map (
            O => \N__22232\,
            I => \N__22229\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__22229\,
            I => \N__22226\
        );

    \I__2818\ : Span12Mux_s9_h
    port map (
            O => \N__22226\,
            I => \N__22223\
        );

    \I__2817\ : Span12Mux_h
    port map (
            O => \N__22223\,
            I => \N__22220\
        );

    \I__2816\ : Odrv12
    port map (
            O => \N__22220\,
            I => \pwm_generator_inst.un2_threshold_2_8\
        );

    \I__2815\ : CascadeMux
    port map (
            O => \N__22217\,
            I => \N__22214\
        );

    \I__2814\ : InMux
    port map (
            O => \N__22214\,
            I => \N__22211\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__22211\,
            I => \N__22208\
        );

    \I__2812\ : Span4Mux_h
    port map (
            O => \N__22208\,
            I => \N__22205\
        );

    \I__2811\ : Odrv4
    port map (
            O => \N__22205\,
            I => \pwm_generator_inst.un2_threshold_1_23\
        );

    \I__2810\ : InMux
    port map (
            O => \N__22202\,
            I => \N__22199\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__22199\,
            I => \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0\
        );

    \I__2808\ : InMux
    port map (
            O => \N__22196\,
            I => \bfn_4_24_0_\
        );

    \I__2807\ : InMux
    port map (
            O => \N__22193\,
            I => \N__22190\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__22190\,
            I => \N__22187\
        );

    \I__2805\ : Span4Mux_h
    port map (
            O => \N__22187\,
            I => \N__22184\
        );

    \I__2804\ : Sp12to4
    port map (
            O => \N__22184\,
            I => \N__22181\
        );

    \I__2803\ : Span12Mux_h
    port map (
            O => \N__22181\,
            I => \N__22178\
        );

    \I__2802\ : Odrv12
    port map (
            O => \N__22178\,
            I => \pwm_generator_inst.un2_threshold_2_9\
        );

    \I__2801\ : CascadeMux
    port map (
            O => \N__22175\,
            I => \N__22172\
        );

    \I__2800\ : InMux
    port map (
            O => \N__22172\,
            I => \N__22169\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__22169\,
            I => \N__22166\
        );

    \I__2798\ : Span4Mux_v
    port map (
            O => \N__22166\,
            I => \N__22163\
        );

    \I__2797\ : Odrv4
    port map (
            O => \N__22163\,
            I => \pwm_generator_inst.un2_threshold_1_24\
        );

    \I__2796\ : InMux
    port map (
            O => \N__22160\,
            I => \N__22157\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__22157\,
            I => \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0\
        );

    \I__2794\ : InMux
    port map (
            O => \N__22154\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_8\
        );

    \I__2793\ : InMux
    port map (
            O => \N__22151\,
            I => \N__22148\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__22148\,
            I => \N__22145\
        );

    \I__2791\ : Span12Mux_s7_h
    port map (
            O => \N__22145\,
            I => \N__22142\
        );

    \I__2790\ : Span12Mux_h
    port map (
            O => \N__22142\,
            I => \N__22139\
        );

    \I__2789\ : Odrv12
    port map (
            O => \N__22139\,
            I => \pwm_generator_inst.un2_threshold_2_10\
        );

    \I__2788\ : InMux
    port map (
            O => \N__22136\,
            I => \N__22133\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__22133\,
            I => \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0\
        );

    \I__2786\ : InMux
    port map (
            O => \N__22130\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_9\
        );

    \I__2785\ : InMux
    port map (
            O => \N__22127\,
            I => \N__22124\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__22124\,
            I => \N__22121\
        );

    \I__2783\ : Span12Mux_s6_h
    port map (
            O => \N__22121\,
            I => \N__22118\
        );

    \I__2782\ : Span12Mux_h
    port map (
            O => \N__22118\,
            I => \N__22115\
        );

    \I__2781\ : Odrv12
    port map (
            O => \N__22115\,
            I => \pwm_generator_inst.un2_threshold_2_11\
        );

    \I__2780\ : InMux
    port map (
            O => \N__22112\,
            I => \N__22109\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__22109\,
            I => \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0\
        );

    \I__2778\ : InMux
    port map (
            O => \N__22106\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_10\
        );

    \I__2777\ : InMux
    port map (
            O => \N__22103\,
            I => \N__22100\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__22100\,
            I => \N__22097\
        );

    \I__2775\ : Sp12to4
    port map (
            O => \N__22097\,
            I => \N__22094\
        );

    \I__2774\ : Span12Mux_h
    port map (
            O => \N__22094\,
            I => \N__22091\
        );

    \I__2773\ : Odrv12
    port map (
            O => \N__22091\,
            I => \pwm_generator_inst.un2_threshold_2_12\
        );

    \I__2772\ : InMux
    port map (
            O => \N__22088\,
            I => \N__22085\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__22085\,
            I => \N__22082\
        );

    \I__2770\ : Odrv4
    port map (
            O => \N__22082\,
            I => \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0\
        );

    \I__2769\ : InMux
    port map (
            O => \N__22079\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_11\
        );

    \I__2768\ : InMux
    port map (
            O => \N__22076\,
            I => \N__22073\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__22073\,
            I => \N__22070\
        );

    \I__2766\ : Span12Mux_h
    port map (
            O => \N__22070\,
            I => \N__22067\
        );

    \I__2765\ : Odrv12
    port map (
            O => \N__22067\,
            I => \pwm_generator_inst.un2_threshold_2_13\
        );

    \I__2764\ : CascadeMux
    port map (
            O => \N__22064\,
            I => \N__22061\
        );

    \I__2763\ : InMux
    port map (
            O => \N__22061\,
            I => \N__22058\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__22058\,
            I => \N__22055\
        );

    \I__2761\ : Odrv4
    port map (
            O => \N__22055\,
            I => \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0\
        );

    \I__2760\ : InMux
    port map (
            O => \N__22052\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_12\
        );

    \I__2759\ : CascadeMux
    port map (
            O => \N__22049\,
            I => \N__22038\
        );

    \I__2758\ : CascadeMux
    port map (
            O => \N__22048\,
            I => \N__22034\
        );

    \I__2757\ : CascadeMux
    port map (
            O => \N__22047\,
            I => \N__22030\
        );

    \I__2756\ : CascadeMux
    port map (
            O => \N__22046\,
            I => \N__22026\
        );

    \I__2755\ : CascadeMux
    port map (
            O => \N__22045\,
            I => \N__22022\
        );

    \I__2754\ : CascadeMux
    port map (
            O => \N__22044\,
            I => \N__22018\
        );

    \I__2753\ : CascadeMux
    port map (
            O => \N__22043\,
            I => \N__22014\
        );

    \I__2752\ : CascadeMux
    port map (
            O => \N__22042\,
            I => \N__22009\
        );

    \I__2751\ : InMux
    port map (
            O => \N__22041\,
            I => \N__21993\
        );

    \I__2750\ : InMux
    port map (
            O => \N__22038\,
            I => \N__21993\
        );

    \I__2749\ : InMux
    port map (
            O => \N__22037\,
            I => \N__21993\
        );

    \I__2748\ : InMux
    port map (
            O => \N__22034\,
            I => \N__21993\
        );

    \I__2747\ : InMux
    port map (
            O => \N__22033\,
            I => \N__21993\
        );

    \I__2746\ : InMux
    port map (
            O => \N__22030\,
            I => \N__21993\
        );

    \I__2745\ : InMux
    port map (
            O => \N__22029\,
            I => \N__21993\
        );

    \I__2744\ : InMux
    port map (
            O => \N__22026\,
            I => \N__21976\
        );

    \I__2743\ : InMux
    port map (
            O => \N__22025\,
            I => \N__21976\
        );

    \I__2742\ : InMux
    port map (
            O => \N__22022\,
            I => \N__21976\
        );

    \I__2741\ : InMux
    port map (
            O => \N__22021\,
            I => \N__21976\
        );

    \I__2740\ : InMux
    port map (
            O => \N__22018\,
            I => \N__21976\
        );

    \I__2739\ : InMux
    port map (
            O => \N__22017\,
            I => \N__21976\
        );

    \I__2738\ : InMux
    port map (
            O => \N__22014\,
            I => \N__21976\
        );

    \I__2737\ : InMux
    port map (
            O => \N__22013\,
            I => \N__21976\
        );

    \I__2736\ : InMux
    port map (
            O => \N__22012\,
            I => \N__21969\
        );

    \I__2735\ : InMux
    port map (
            O => \N__22009\,
            I => \N__21969\
        );

    \I__2734\ : InMux
    port map (
            O => \N__22008\,
            I => \N__21969\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__21993\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__21976\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__21969\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\
        );

    \I__2730\ : InMux
    port map (
            O => \N__21962\,
            I => \N__21959\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__21959\,
            I => \N__21956\
        );

    \I__2728\ : Span12Mux_s9_h
    port map (
            O => \N__21956\,
            I => \N__21953\
        );

    \I__2727\ : Span12Mux_h
    port map (
            O => \N__21953\,
            I => \N__21950\
        );

    \I__2726\ : Odrv12
    port map (
            O => \N__21950\,
            I => \pwm_generator_inst.un2_threshold_2_0\
        );

    \I__2725\ : CascadeMux
    port map (
            O => \N__21947\,
            I => \N__21944\
        );

    \I__2724\ : InMux
    port map (
            O => \N__21944\,
            I => \N__21941\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__21941\,
            I => \N__21938\
        );

    \I__2722\ : Span4Mux_h
    port map (
            O => \N__21938\,
            I => \N__21935\
        );

    \I__2721\ : Odrv4
    port map (
            O => \N__21935\,
            I => \pwm_generator_inst.un2_threshold_1_15\
        );

    \I__2720\ : InMux
    port map (
            O => \N__21932\,
            I => \N__21929\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__21929\,
            I => \pwm_generator_inst.un3_threshold_axbZ0Z_4\
        );

    \I__2718\ : InMux
    port map (
            O => \N__21926\,
            I => \N__21923\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__21923\,
            I => \N__21920\
        );

    \I__2716\ : Span4Mux_h
    port map (
            O => \N__21920\,
            I => \N__21917\
        );

    \I__2715\ : Sp12to4
    port map (
            O => \N__21917\,
            I => \N__21914\
        );

    \I__2714\ : Span12Mux_h
    port map (
            O => \N__21914\,
            I => \N__21911\
        );

    \I__2713\ : Odrv12
    port map (
            O => \N__21911\,
            I => \pwm_generator_inst.un2_threshold_2_1\
        );

    \I__2712\ : CascadeMux
    port map (
            O => \N__21908\,
            I => \N__21905\
        );

    \I__2711\ : InMux
    port map (
            O => \N__21905\,
            I => \N__21902\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__21902\,
            I => \N__21899\
        );

    \I__2709\ : Span4Mux_h
    port map (
            O => \N__21899\,
            I => \N__21896\
        );

    \I__2708\ : Odrv4
    port map (
            O => \N__21896\,
            I => \pwm_generator_inst.un2_threshold_1_16\
        );

    \I__2707\ : CascadeMux
    port map (
            O => \N__21893\,
            I => \N__21890\
        );

    \I__2706\ : InMux
    port map (
            O => \N__21890\,
            I => \N__21887\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__21887\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701\
        );

    \I__2704\ : InMux
    port map (
            O => \N__21884\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_0\
        );

    \I__2703\ : InMux
    port map (
            O => \N__21881\,
            I => \N__21878\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__21878\,
            I => \N__21875\
        );

    \I__2701\ : Span12Mux_s7_h
    port map (
            O => \N__21875\,
            I => \N__21872\
        );

    \I__2700\ : Span12Mux_h
    port map (
            O => \N__21872\,
            I => \N__21869\
        );

    \I__2699\ : Odrv12
    port map (
            O => \N__21869\,
            I => \pwm_generator_inst.un2_threshold_2_2\
        );

    \I__2698\ : CascadeMux
    port map (
            O => \N__21866\,
            I => \N__21863\
        );

    \I__2697\ : InMux
    port map (
            O => \N__21863\,
            I => \N__21860\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__21860\,
            I => \N__21857\
        );

    \I__2695\ : Span4Mux_h
    port map (
            O => \N__21857\,
            I => \N__21854\
        );

    \I__2694\ : Odrv4
    port map (
            O => \N__21854\,
            I => \pwm_generator_inst.un2_threshold_1_17\
        );

    \I__2693\ : InMux
    port map (
            O => \N__21851\,
            I => \N__21848\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__21848\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801\
        );

    \I__2691\ : InMux
    port map (
            O => \N__21845\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_1\
        );

    \I__2690\ : InMux
    port map (
            O => \N__21842\,
            I => \N__21839\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__21839\,
            I => \N__21836\
        );

    \I__2688\ : Span12Mux_s6_h
    port map (
            O => \N__21836\,
            I => \N__21833\
        );

    \I__2687\ : Span12Mux_h
    port map (
            O => \N__21833\,
            I => \N__21830\
        );

    \I__2686\ : Odrv12
    port map (
            O => \N__21830\,
            I => \pwm_generator_inst.un2_threshold_2_3\
        );

    \I__2685\ : CascadeMux
    port map (
            O => \N__21827\,
            I => \N__21824\
        );

    \I__2684\ : InMux
    port map (
            O => \N__21824\,
            I => \N__21821\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__21821\,
            I => \N__21818\
        );

    \I__2682\ : Span4Mux_v
    port map (
            O => \N__21818\,
            I => \N__21815\
        );

    \I__2681\ : Odrv4
    port map (
            O => \N__21815\,
            I => \pwm_generator_inst.un2_threshold_1_18\
        );

    \I__2680\ : CascadeMux
    port map (
            O => \N__21812\,
            I => \N__21809\
        );

    \I__2679\ : InMux
    port map (
            O => \N__21809\,
            I => \N__21806\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__21806\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901\
        );

    \I__2677\ : InMux
    port map (
            O => \N__21803\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_2\
        );

    \I__2676\ : InMux
    port map (
            O => \N__21800\,
            I => \N__21797\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__21797\,
            I => \N__21794\
        );

    \I__2674\ : Span4Mux_v
    port map (
            O => \N__21794\,
            I => \N__21791\
        );

    \I__2673\ : Odrv4
    port map (
            O => \N__21791\,
            I => \pwm_generator_inst.un2_threshold_1_19\
        );

    \I__2672\ : CascadeMux
    port map (
            O => \N__21788\,
            I => \N__21785\
        );

    \I__2671\ : InMux
    port map (
            O => \N__21785\,
            I => \N__21782\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__21782\,
            I => \N__21779\
        );

    \I__2669\ : Span12Mux_s5_h
    port map (
            O => \N__21779\,
            I => \N__21776\
        );

    \I__2668\ : Span12Mux_h
    port map (
            O => \N__21776\,
            I => \N__21773\
        );

    \I__2667\ : Odrv12
    port map (
            O => \N__21773\,
            I => \pwm_generator_inst.un2_threshold_2_4\
        );

    \I__2666\ : InMux
    port map (
            O => \N__21770\,
            I => \N__21767\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__21767\,
            I => \N__21764\
        );

    \I__2664\ : Odrv4
    port map (
            O => \N__21764\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01\
        );

    \I__2663\ : InMux
    port map (
            O => \N__21761\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_3\
        );

    \I__2662\ : InMux
    port map (
            O => \N__21758\,
            I => \N__21755\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__21755\,
            I => \N__21752\
        );

    \I__2660\ : Span4Mux_h
    port map (
            O => \N__21752\,
            I => \N__21749\
        );

    \I__2659\ : Odrv4
    port map (
            O => \N__21749\,
            I => \pwm_generator_inst.un2_threshold_1_20\
        );

    \I__2658\ : CascadeMux
    port map (
            O => \N__21746\,
            I => \N__21743\
        );

    \I__2657\ : InMux
    port map (
            O => \N__21743\,
            I => \N__21740\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__21740\,
            I => \N__21737\
        );

    \I__2655\ : Span12Mux_h
    port map (
            O => \N__21737\,
            I => \N__21734\
        );

    \I__2654\ : Odrv12
    port map (
            O => \N__21734\,
            I => \pwm_generator_inst.un2_threshold_2_5\
        );

    \I__2653\ : CascadeMux
    port map (
            O => \N__21731\,
            I => \N__21728\
        );

    \I__2652\ : InMux
    port map (
            O => \N__21728\,
            I => \N__21725\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__21725\,
            I => \N__21722\
        );

    \I__2650\ : Odrv4
    port map (
            O => \N__21722\,
            I => \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0\
        );

    \I__2649\ : InMux
    port map (
            O => \N__21719\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_4\
        );

    \I__2648\ : InMux
    port map (
            O => \N__21716\,
            I => \N__21713\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__21713\,
            I => \N__21710\
        );

    \I__2646\ : Span4Mux_h
    port map (
            O => \N__21710\,
            I => \N__21707\
        );

    \I__2645\ : Odrv4
    port map (
            O => \N__21707\,
            I => \pwm_generator_inst.un2_threshold_1_21\
        );

    \I__2644\ : CascadeMux
    port map (
            O => \N__21704\,
            I => \N__21701\
        );

    \I__2643\ : InMux
    port map (
            O => \N__21701\,
            I => \N__21698\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__21698\,
            I => \N__21695\
        );

    \I__2641\ : Span12Mux_h
    port map (
            O => \N__21695\,
            I => \N__21692\
        );

    \I__2640\ : Odrv12
    port map (
            O => \N__21692\,
            I => \pwm_generator_inst.un2_threshold_2_6\
        );

    \I__2639\ : InMux
    port map (
            O => \N__21689\,
            I => \N__21686\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__21686\,
            I => \N__21683\
        );

    \I__2637\ : Odrv4
    port map (
            O => \N__21683\,
            I => \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0\
        );

    \I__2636\ : InMux
    port map (
            O => \N__21680\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_5\
        );

    \I__2635\ : CascadeMux
    port map (
            O => \N__21677\,
            I => \N__21674\
        );

    \I__2634\ : InMux
    port map (
            O => \N__21674\,
            I => \N__21671\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__21671\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\
        );

    \I__2632\ : InMux
    port map (
            O => \N__21668\,
            I => \N__21665\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__21665\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\
        );

    \I__2630\ : InMux
    port map (
            O => \N__21662\,
            I => \N__21659\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__21659\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\
        );

    \I__2628\ : InMux
    port map (
            O => \N__21656\,
            I => \N__21653\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__21653\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\
        );

    \I__2626\ : InMux
    port map (
            O => \N__21650\,
            I => \N__21647\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__21647\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\
        );

    \I__2624\ : InMux
    port map (
            O => \N__21644\,
            I => \N__21641\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__21641\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\
        );

    \I__2622\ : InMux
    port map (
            O => \N__21638\,
            I => \N__21634\
        );

    \I__2621\ : InMux
    port map (
            O => \N__21637\,
            I => \N__21631\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__21634\,
            I => \N__21628\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__21631\,
            I => \N__21625\
        );

    \I__2618\ : Span4Mux_h
    port map (
            O => \N__21628\,
            I => \N__21622\
        );

    \I__2617\ : Odrv4
    port map (
            O => \N__21625\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__2616\ : Odrv4
    port map (
            O => \N__21622\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__2615\ : InMux
    port map (
            O => \N__21617\,
            I => \N__21614\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__21614\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\
        );

    \I__2613\ : InMux
    port map (
            O => \N__21611\,
            I => \N__21608\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__21608\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\
        );

    \I__2611\ : InMux
    port map (
            O => \N__21605\,
            I => \N__21602\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__21602\,
            I => \N__21599\
        );

    \I__2609\ : Span4Mux_v
    port map (
            O => \N__21599\,
            I => \N__21593\
        );

    \I__2608\ : InMux
    port map (
            O => \N__21598\,
            I => \N__21590\
        );

    \I__2607\ : InMux
    port map (
            O => \N__21597\,
            I => \N__21587\
        );

    \I__2606\ : InMux
    port map (
            O => \N__21596\,
            I => \N__21584\
        );

    \I__2605\ : Odrv4
    port map (
            O => \N__21593\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__21590\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__21587\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__21584\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__2601\ : InMux
    port map (
            O => \N__21575\,
            I => \N__21571\
        );

    \I__2600\ : CascadeMux
    port map (
            O => \N__21574\,
            I => \N__21567\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__21571\,
            I => \N__21563\
        );

    \I__2598\ : InMux
    port map (
            O => \N__21570\,
            I => \N__21560\
        );

    \I__2597\ : InMux
    port map (
            O => \N__21567\,
            I => \N__21557\
        );

    \I__2596\ : InMux
    port map (
            O => \N__21566\,
            I => \N__21554\
        );

    \I__2595\ : Odrv12
    port map (
            O => \N__21563\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__21560\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__21557\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__21554\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__2591\ : CascadeMux
    port map (
            O => \N__21545\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_\
        );

    \I__2590\ : InMux
    port map (
            O => \N__21542\,
            I => \N__21539\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__21539\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\
        );

    \I__2588\ : CascadeMux
    port map (
            O => \N__21536\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_\
        );

    \I__2587\ : InMux
    port map (
            O => \N__21533\,
            I => \N__21530\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__21530\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\
        );

    \I__2585\ : InMux
    port map (
            O => \N__21527\,
            I => \N__21524\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__21524\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\
        );

    \I__2583\ : InMux
    port map (
            O => \N__21521\,
            I => \N__21518\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__21518\,
            I => \N__21512\
        );

    \I__2581\ : InMux
    port map (
            O => \N__21517\,
            I => \N__21509\
        );

    \I__2580\ : InMux
    port map (
            O => \N__21516\,
            I => \N__21504\
        );

    \I__2579\ : InMux
    port map (
            O => \N__21515\,
            I => \N__21504\
        );

    \I__2578\ : Odrv12
    port map (
            O => \N__21512\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__21509\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__21504\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__2575\ : InMux
    port map (
            O => \N__21497\,
            I => \N__21494\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__21494\,
            I => \N__21488\
        );

    \I__2573\ : InMux
    port map (
            O => \N__21493\,
            I => \N__21485\
        );

    \I__2572\ : InMux
    port map (
            O => \N__21492\,
            I => \N__21480\
        );

    \I__2571\ : InMux
    port map (
            O => \N__21491\,
            I => \N__21480\
        );

    \I__2570\ : Odrv12
    port map (
            O => \N__21488\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__21485\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__21480\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__2567\ : CascadeMux
    port map (
            O => \N__21473\,
            I => \N__21470\
        );

    \I__2566\ : InMux
    port map (
            O => \N__21470\,
            I => \N__21467\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__21467\,
            I => \N__21463\
        );

    \I__2564\ : CascadeMux
    port map (
            O => \N__21466\,
            I => \N__21459\
        );

    \I__2563\ : Span4Mux_v
    port map (
            O => \N__21463\,
            I => \N__21455\
        );

    \I__2562\ : InMux
    port map (
            O => \N__21462\,
            I => \N__21452\
        );

    \I__2561\ : InMux
    port map (
            O => \N__21459\,
            I => \N__21447\
        );

    \I__2560\ : InMux
    port map (
            O => \N__21458\,
            I => \N__21447\
        );

    \I__2559\ : Odrv4
    port map (
            O => \N__21455\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__21452\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__21447\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__2556\ : CascadeMux
    port map (
            O => \N__21440\,
            I => \N__21436\
        );

    \I__2555\ : CascadeMux
    port map (
            O => \N__21439\,
            I => \N__21432\
        );

    \I__2554\ : InMux
    port map (
            O => \N__21436\,
            I => \N__21429\
        );

    \I__2553\ : InMux
    port map (
            O => \N__21435\,
            I => \N__21424\
        );

    \I__2552\ : InMux
    port map (
            O => \N__21432\,
            I => \N__21424\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__21429\,
            I => \N__21420\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__21424\,
            I => \N__21417\
        );

    \I__2549\ : InMux
    port map (
            O => \N__21423\,
            I => \N__21414\
        );

    \I__2548\ : Span4Mux_v
    port map (
            O => \N__21420\,
            I => \N__21409\
        );

    \I__2547\ : Span4Mux_h
    port map (
            O => \N__21417\,
            I => \N__21409\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__21414\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__2545\ : Odrv4
    port map (
            O => \N__21409\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__2544\ : CascadeMux
    port map (
            O => \N__21404\,
            I => \N__21401\
        );

    \I__2543\ : InMux
    port map (
            O => \N__21401\,
            I => \N__21398\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__21398\,
            I => \N__21393\
        );

    \I__2541\ : InMux
    port map (
            O => \N__21397\,
            I => \N__21390\
        );

    \I__2540\ : InMux
    port map (
            O => \N__21396\,
            I => \N__21386\
        );

    \I__2539\ : Span4Mux_v
    port map (
            O => \N__21393\,
            I => \N__21381\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__21390\,
            I => \N__21381\
        );

    \I__2537\ : InMux
    port map (
            O => \N__21389\,
            I => \N__21378\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__21386\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__2535\ : Odrv4
    port map (
            O => \N__21381\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__21378\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__2533\ : CascadeMux
    port map (
            O => \N__21371\,
            I => \N__21368\
        );

    \I__2532\ : InMux
    port map (
            O => \N__21368\,
            I => \N__21365\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__21365\,
            I => \N__21360\
        );

    \I__2530\ : InMux
    port map (
            O => \N__21364\,
            I => \N__21357\
        );

    \I__2529\ : InMux
    port map (
            O => \N__21363\,
            I => \N__21353\
        );

    \I__2528\ : Span4Mux_v
    port map (
            O => \N__21360\,
            I => \N__21348\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__21357\,
            I => \N__21348\
        );

    \I__2526\ : InMux
    port map (
            O => \N__21356\,
            I => \N__21345\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__21353\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__2524\ : Odrv4
    port map (
            O => \N__21348\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__21345\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__2522\ : InMux
    port map (
            O => \N__21338\,
            I => \N__21335\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__21335\,
            I => \N__21329\
        );

    \I__2520\ : InMux
    port map (
            O => \N__21334\,
            I => \N__21326\
        );

    \I__2519\ : InMux
    port map (
            O => \N__21333\,
            I => \N__21321\
        );

    \I__2518\ : InMux
    port map (
            O => \N__21332\,
            I => \N__21321\
        );

    \I__2517\ : Odrv12
    port map (
            O => \N__21329\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__21326\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__21321\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__2514\ : CascadeMux
    port map (
            O => \N__21314\,
            I => \N__21310\
        );

    \I__2513\ : CascadeMux
    port map (
            O => \N__21313\,
            I => \N__21306\
        );

    \I__2512\ : InMux
    port map (
            O => \N__21310\,
            I => \N__21303\
        );

    \I__2511\ : InMux
    port map (
            O => \N__21309\,
            I => \N__21300\
        );

    \I__2510\ : InMux
    port map (
            O => \N__21306\,
            I => \N__21297\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__21303\,
            I => \N__21293\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__21300\,
            I => \N__21288\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__21297\,
            I => \N__21288\
        );

    \I__2506\ : InMux
    port map (
            O => \N__21296\,
            I => \N__21285\
        );

    \I__2505\ : Span4Mux_v
    port map (
            O => \N__21293\,
            I => \N__21280\
        );

    \I__2504\ : Span4Mux_v
    port map (
            O => \N__21288\,
            I => \N__21280\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__21285\,
            I => \N__21277\
        );

    \I__2502\ : Odrv4
    port map (
            O => \N__21280\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__2501\ : Odrv4
    port map (
            O => \N__21277\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__2500\ : CascadeMux
    port map (
            O => \N__21272\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_\
        );

    \I__2499\ : InMux
    port map (
            O => \N__21269\,
            I => \N__21266\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__21266\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15\
        );

    \I__2497\ : InMux
    port map (
            O => \N__21263\,
            I => \N__21260\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__21260\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\
        );

    \I__2495\ : InMux
    port map (
            O => \N__21257\,
            I => \N__21254\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__21254\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\
        );

    \I__2493\ : CascadeMux
    port map (
            O => \N__21251\,
            I => \N__21248\
        );

    \I__2492\ : InMux
    port map (
            O => \N__21248\,
            I => \N__21245\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__21245\,
            I => \N__21241\
        );

    \I__2490\ : InMux
    port map (
            O => \N__21244\,
            I => \N__21236\
        );

    \I__2489\ : Span4Mux_v
    port map (
            O => \N__21241\,
            I => \N__21233\
        );

    \I__2488\ : InMux
    port map (
            O => \N__21240\,
            I => \N__21228\
        );

    \I__2487\ : InMux
    port map (
            O => \N__21239\,
            I => \N__21228\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__21236\,
            I => \N__21225\
        );

    \I__2485\ : Odrv4
    port map (
            O => \N__21233\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__21228\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__2483\ : Odrv4
    port map (
            O => \N__21225\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__2482\ : InMux
    port map (
            O => \N__21218\,
            I => \N__21215\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__21215\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_2\
        );

    \I__2480\ : InMux
    port map (
            O => \N__21212\,
            I => \N__21209\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__21209\,
            I => \N__21206\
        );

    \I__2478\ : Odrv12
    port map (
            O => \N__21206\,
            I => \current_shift_inst.PI_CTRL.N_43\
        );

    \I__2477\ : InMux
    port map (
            O => \N__21203\,
            I => \N__21200\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__21200\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\
        );

    \I__2475\ : CascadeMux
    port map (
            O => \N__21197\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15_cascade_\
        );

    \I__2474\ : InMux
    port map (
            O => \N__21194\,
            I => \N__21191\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__21191\,
            I => \N__21188\
        );

    \I__2472\ : Span4Mux_v
    port map (
            O => \N__21188\,
            I => \N__21182\
        );

    \I__2471\ : InMux
    port map (
            O => \N__21187\,
            I => \N__21179\
        );

    \I__2470\ : InMux
    port map (
            O => \N__21186\,
            I => \N__21174\
        );

    \I__2469\ : InMux
    port map (
            O => \N__21185\,
            I => \N__21174\
        );

    \I__2468\ : Odrv4
    port map (
            O => \N__21182\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__21179\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__21174\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__2465\ : CascadeMux
    port map (
            O => \N__21167\,
            I => \N__21164\
        );

    \I__2464\ : InMux
    port map (
            O => \N__21164\,
            I => \N__21161\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__21161\,
            I => \N__21158\
        );

    \I__2462\ : Span4Mux_v
    port map (
            O => \N__21158\,
            I => \N__21152\
        );

    \I__2461\ : InMux
    port map (
            O => \N__21157\,
            I => \N__21149\
        );

    \I__2460\ : InMux
    port map (
            O => \N__21156\,
            I => \N__21144\
        );

    \I__2459\ : InMux
    port map (
            O => \N__21155\,
            I => \N__21144\
        );

    \I__2458\ : Odrv4
    port map (
            O => \N__21152\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__21149\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__21144\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__2455\ : CascadeMux
    port map (
            O => \N__21137\,
            I => \N__21134\
        );

    \I__2454\ : InMux
    port map (
            O => \N__21134\,
            I => \N__21131\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__21131\,
            I => \N__21126\
        );

    \I__2452\ : CascadeMux
    port map (
            O => \N__21130\,
            I => \N__21123\
        );

    \I__2451\ : CascadeMux
    port map (
            O => \N__21129\,
            I => \N__21120\
        );

    \I__2450\ : Span4Mux_v
    port map (
            O => \N__21126\,
            I => \N__21116\
        );

    \I__2449\ : InMux
    port map (
            O => \N__21123\,
            I => \N__21111\
        );

    \I__2448\ : InMux
    port map (
            O => \N__21120\,
            I => \N__21111\
        );

    \I__2447\ : InMux
    port map (
            O => \N__21119\,
            I => \N__21108\
        );

    \I__2446\ : Odrv4
    port map (
            O => \N__21116\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__21111\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__21108\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__2443\ : CascadeMux
    port map (
            O => \N__21101\,
            I => \N__21098\
        );

    \I__2442\ : InMux
    port map (
            O => \N__21098\,
            I => \N__21095\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__21095\,
            I => \N__21092\
        );

    \I__2440\ : Span4Mux_v
    port map (
            O => \N__21092\,
            I => \N__21086\
        );

    \I__2439\ : InMux
    port map (
            O => \N__21091\,
            I => \N__21083\
        );

    \I__2438\ : InMux
    port map (
            O => \N__21090\,
            I => \N__21080\
        );

    \I__2437\ : InMux
    port map (
            O => \N__21089\,
            I => \N__21077\
        );

    \I__2436\ : Odrv4
    port map (
            O => \N__21086\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__21083\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__21080\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__21077\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__2432\ : CascadeMux
    port map (
            O => \N__21068\,
            I => \N__21065\
        );

    \I__2431\ : InMux
    port map (
            O => \N__21065\,
            I => \N__21062\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__21062\,
            I => \N__21056\
        );

    \I__2429\ : InMux
    port map (
            O => \N__21061\,
            I => \N__21053\
        );

    \I__2428\ : InMux
    port map (
            O => \N__21060\,
            I => \N__21048\
        );

    \I__2427\ : InMux
    port map (
            O => \N__21059\,
            I => \N__21048\
        );

    \I__2426\ : Odrv12
    port map (
            O => \N__21056\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__21053\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__21048\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__2423\ : InMux
    port map (
            O => \N__21041\,
            I => \N__21038\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__21038\,
            I => \N__21033\
        );

    \I__2421\ : InMux
    port map (
            O => \N__21037\,
            I => \N__21027\
        );

    \I__2420\ : InMux
    port map (
            O => \N__21036\,
            I => \N__21027\
        );

    \I__2419\ : Span12Mux_h
    port map (
            O => \N__21033\,
            I => \N__21024\
        );

    \I__2418\ : InMux
    port map (
            O => \N__21032\,
            I => \N__21021\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__21027\,
            I => \N__21018\
        );

    \I__2416\ : Odrv12
    port map (
            O => \N__21024\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__21021\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__2414\ : Odrv4
    port map (
            O => \N__21018\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__2413\ : InMux
    port map (
            O => \N__21011\,
            I => \N__21006\
        );

    \I__2412\ : CascadeMux
    port map (
            O => \N__21010\,
            I => \N__21002\
        );

    \I__2411\ : CascadeMux
    port map (
            O => \N__21009\,
            I => \N__20999\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__21006\,
            I => \N__20996\
        );

    \I__2409\ : InMux
    port map (
            O => \N__21005\,
            I => \N__20993\
        );

    \I__2408\ : InMux
    port map (
            O => \N__21002\,
            I => \N__20988\
        );

    \I__2407\ : InMux
    port map (
            O => \N__20999\,
            I => \N__20988\
        );

    \I__2406\ : Odrv12
    port map (
            O => \N__20996\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__20993\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__20988\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__2403\ : CascadeMux
    port map (
            O => \N__20981\,
            I => \N__20978\
        );

    \I__2402\ : InMux
    port map (
            O => \N__20978\,
            I => \N__20975\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__20975\,
            I => \N__20969\
        );

    \I__2400\ : InMux
    port map (
            O => \N__20974\,
            I => \N__20966\
        );

    \I__2399\ : InMux
    port map (
            O => \N__20973\,
            I => \N__20961\
        );

    \I__2398\ : InMux
    port map (
            O => \N__20972\,
            I => \N__20961\
        );

    \I__2397\ : Odrv12
    port map (
            O => \N__20969\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__20966\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__20961\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__2394\ : CascadeMux
    port map (
            O => \N__20954\,
            I => \N__20951\
        );

    \I__2393\ : InMux
    port map (
            O => \N__20951\,
            I => \N__20948\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__20948\,
            I => \N__20942\
        );

    \I__2391\ : InMux
    port map (
            O => \N__20947\,
            I => \N__20939\
        );

    \I__2390\ : InMux
    port map (
            O => \N__20946\,
            I => \N__20936\
        );

    \I__2389\ : InMux
    port map (
            O => \N__20945\,
            I => \N__20933\
        );

    \I__2388\ : Odrv4
    port map (
            O => \N__20942\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__20939\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__20936\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__20933\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__2384\ : InMux
    port map (
            O => \N__20924\,
            I => \pwm_generator_inst.un3_threshold_cry_19\
        );

    \I__2383\ : InMux
    port map (
            O => \N__20921\,
            I => \N__20918\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__20918\,
            I => \N__20915\
        );

    \I__2381\ : Span12Mux_h
    port map (
            O => \N__20915\,
            I => \N__20912\
        );

    \I__2380\ : Odrv12
    port map (
            O => \N__20912\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\
        );

    \I__2379\ : CascadeMux
    port map (
            O => \N__20909\,
            I => \N__20906\
        );

    \I__2378\ : InMux
    port map (
            O => \N__20906\,
            I => \N__20903\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__20903\,
            I => \N__20900\
        );

    \I__2376\ : Odrv4
    port map (
            O => \N__20900\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\
        );

    \I__2375\ : CascadeMux
    port map (
            O => \N__20897\,
            I => \N__20894\
        );

    \I__2374\ : InMux
    port map (
            O => \N__20894\,
            I => \N__20891\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__20891\,
            I => \N__20888\
        );

    \I__2372\ : Odrv12
    port map (
            O => \N__20888\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\
        );

    \I__2371\ : CascadeMux
    port map (
            O => \N__20885\,
            I => \N__20881\
        );

    \I__2370\ : InMux
    port map (
            O => \N__20884\,
            I => \N__20877\
        );

    \I__2369\ : InMux
    port map (
            O => \N__20881\,
            I => \N__20874\
        );

    \I__2368\ : InMux
    port map (
            O => \N__20880\,
            I => \N__20871\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__20877\,
            I => \N__20868\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__20874\,
            I => \N__20865\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__20871\,
            I => \N__20862\
        );

    \I__2364\ : Span4Mux_h
    port map (
            O => \N__20868\,
            I => \N__20859\
        );

    \I__2363\ : Span4Mux_h
    port map (
            O => \N__20865\,
            I => \N__20856\
        );

    \I__2362\ : Span4Mux_v
    port map (
            O => \N__20862\,
            I => \N__20853\
        );

    \I__2361\ : Odrv4
    port map (
            O => \N__20859\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__2360\ : Odrv4
    port map (
            O => \N__20856\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__2359\ : Odrv4
    port map (
            O => \N__20853\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__2358\ : CascadeMux
    port map (
            O => \N__20846\,
            I => \N__20842\
        );

    \I__2357\ : InMux
    port map (
            O => \N__20845\,
            I => \N__20839\
        );

    \I__2356\ : InMux
    port map (
            O => \N__20842\,
            I => \N__20835\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__20839\,
            I => \N__20831\
        );

    \I__2354\ : CascadeMux
    port map (
            O => \N__20838\,
            I => \N__20828\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__20835\,
            I => \N__20825\
        );

    \I__2352\ : InMux
    port map (
            O => \N__20834\,
            I => \N__20821\
        );

    \I__2351\ : Span4Mux_v
    port map (
            O => \N__20831\,
            I => \N__20818\
        );

    \I__2350\ : InMux
    port map (
            O => \N__20828\,
            I => \N__20815\
        );

    \I__2349\ : Span4Mux_h
    port map (
            O => \N__20825\,
            I => \N__20812\
        );

    \I__2348\ : InMux
    port map (
            O => \N__20824\,
            I => \N__20809\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__20821\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__2346\ : Odrv4
    port map (
            O => \N__20818\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__20815\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__2344\ : Odrv4
    port map (
            O => \N__20812\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__20809\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__2342\ : CascadeMux
    port map (
            O => \N__20798\,
            I => \current_shift_inst.PI_CTRL.N_77_cascade_\
        );

    \I__2341\ : CascadeMux
    port map (
            O => \N__20795\,
            I => \N__20792\
        );

    \I__2340\ : InMux
    port map (
            O => \N__20792\,
            I => \N__20788\
        );

    \I__2339\ : InMux
    port map (
            O => \N__20791\,
            I => \N__20784\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__20788\,
            I => \N__20781\
        );

    \I__2337\ : InMux
    port map (
            O => \N__20787\,
            I => \N__20777\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__20784\,
            I => \N__20774\
        );

    \I__2335\ : Span4Mux_v
    port map (
            O => \N__20781\,
            I => \N__20771\
        );

    \I__2334\ : InMux
    port map (
            O => \N__20780\,
            I => \N__20768\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__20777\,
            I => \N__20765\
        );

    \I__2332\ : Odrv4
    port map (
            O => \N__20774\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__2331\ : Odrv4
    port map (
            O => \N__20771\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__20768\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__2329\ : Odrv4
    port map (
            O => \N__20765\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__2328\ : InMux
    port map (
            O => \N__20756\,
            I => \N__20753\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__20753\,
            I => \N__20750\
        );

    \I__2326\ : Odrv4
    port map (
            O => \N__20750\,
            I => \pwm_generator_inst.O_12\
        );

    \I__2325\ : InMux
    port map (
            O => \N__20747\,
            I => \pwm_generator_inst.un3_threshold_cry_0\
        );

    \I__2324\ : InMux
    port map (
            O => \N__20744\,
            I => \N__20741\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__20741\,
            I => \N__20738\
        );

    \I__2322\ : Odrv4
    port map (
            O => \N__20738\,
            I => \pwm_generator_inst.O_13\
        );

    \I__2321\ : InMux
    port map (
            O => \N__20735\,
            I => \pwm_generator_inst.un3_threshold_cry_1\
        );

    \I__2320\ : InMux
    port map (
            O => \N__20732\,
            I => \N__20729\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__20729\,
            I => \N__20726\
        );

    \I__2318\ : Odrv12
    port map (
            O => \N__20726\,
            I => \pwm_generator_inst.O_14\
        );

    \I__2317\ : InMux
    port map (
            O => \N__20723\,
            I => \pwm_generator_inst.un3_threshold_cry_2\
        );

    \I__2316\ : InMux
    port map (
            O => \N__20720\,
            I => \pwm_generator_inst.un3_threshold_cry_3\
        );

    \I__2315\ : InMux
    port map (
            O => \N__20717\,
            I => \pwm_generator_inst.un3_threshold_cry_4\
        );

    \I__2314\ : InMux
    port map (
            O => \N__20714\,
            I => \pwm_generator_inst.un3_threshold_cry_5\
        );

    \I__2313\ : InMux
    port map (
            O => \N__20711\,
            I => \pwm_generator_inst.un3_threshold_cry_6\
        );

    \I__2312\ : InMux
    port map (
            O => \N__20708\,
            I => \bfn_3_25_0_\
        );

    \I__2311\ : CascadeMux
    port map (
            O => \N__20705\,
            I => \N__20701\
        );

    \I__2310\ : InMux
    port map (
            O => \N__20704\,
            I => \N__20696\
        );

    \I__2309\ : InMux
    port map (
            O => \N__20701\,
            I => \N__20696\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__20696\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__2307\ : InMux
    port map (
            O => \N__20693\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\
        );

    \I__2306\ : InMux
    port map (
            O => \N__20690\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\
        );

    \I__2305\ : InMux
    port map (
            O => \N__20687\,
            I => \N__20683\
        );

    \I__2304\ : CascadeMux
    port map (
            O => \N__20686\,
            I => \N__20680\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__20683\,
            I => \N__20676\
        );

    \I__2302\ : InMux
    port map (
            O => \N__20680\,
            I => \N__20673\
        );

    \I__2301\ : InMux
    port map (
            O => \N__20679\,
            I => \N__20670\
        );

    \I__2300\ : Span4Mux_v
    port map (
            O => \N__20676\,
            I => \N__20664\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__20673\,
            I => \N__20664\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__20670\,
            I => \N__20661\
        );

    \I__2297\ : InMux
    port map (
            O => \N__20669\,
            I => \N__20658\
        );

    \I__2296\ : Span4Mux_v
    port map (
            O => \N__20664\,
            I => \N__20655\
        );

    \I__2295\ : Sp12to4
    port map (
            O => \N__20661\,
            I => \N__20650\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__20658\,
            I => \N__20650\
        );

    \I__2293\ : Odrv4
    port map (
            O => \N__20655\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2292\ : Odrv12
    port map (
            O => \N__20650\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2291\ : InMux
    port map (
            O => \N__20645\,
            I => \N__20642\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__20642\,
            I => \N__20638\
        );

    \I__2289\ : InMux
    port map (
            O => \N__20641\,
            I => \N__20635\
        );

    \I__2288\ : Span4Mux_s3_h
    port map (
            O => \N__20638\,
            I => \N__20631\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__20635\,
            I => \N__20628\
        );

    \I__2286\ : InMux
    port map (
            O => \N__20634\,
            I => \N__20625\
        );

    \I__2285\ : Span4Mux_v
    port map (
            O => \N__20631\,
            I => \N__20622\
        );

    \I__2284\ : Sp12to4
    port map (
            O => \N__20628\,
            I => \N__20617\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__20625\,
            I => \N__20617\
        );

    \I__2282\ : Odrv4
    port map (
            O => \N__20622\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__2281\ : Odrv12
    port map (
            O => \N__20617\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__2280\ : InMux
    port map (
            O => \N__20612\,
            I => \N__20609\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__20609\,
            I => \current_shift_inst.PI_CTRL.N_98\
        );

    \I__2278\ : CascadeMux
    port map (
            O => \N__20606\,
            I => \N__20603\
        );

    \I__2277\ : InMux
    port map (
            O => \N__20603\,
            I => \N__20600\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__20600\,
            I => \N__20596\
        );

    \I__2275\ : InMux
    port map (
            O => \N__20599\,
            I => \N__20593\
        );

    \I__2274\ : Span4Mux_v
    port map (
            O => \N__20596\,
            I => \N__20590\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__20593\,
            I => \N__20587\
        );

    \I__2272\ : Odrv4
    port map (
            O => \N__20590\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__2271\ : Odrv4
    port map (
            O => \N__20587\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__2270\ : InMux
    port map (
            O => \N__20582\,
            I => \N__20578\
        );

    \I__2269\ : InMux
    port map (
            O => \N__20581\,
            I => \N__20575\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__20578\,
            I => \N__20572\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__20575\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__2266\ : Odrv4
    port map (
            O => \N__20572\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__2265\ : CascadeMux
    port map (
            O => \N__20567\,
            I => \N__20564\
        );

    \I__2264\ : InMux
    port map (
            O => \N__20564\,
            I => \N__20560\
        );

    \I__2263\ : InMux
    port map (
            O => \N__20563\,
            I => \N__20557\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__20560\,
            I => \N__20552\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__20557\,
            I => \N__20552\
        );

    \I__2260\ : Odrv4
    port map (
            O => \N__20552\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__2259\ : CascadeMux
    port map (
            O => \N__20549\,
            I => \N__20545\
        );

    \I__2258\ : InMux
    port map (
            O => \N__20548\,
            I => \N__20542\
        );

    \I__2257\ : InMux
    port map (
            O => \N__20545\,
            I => \N__20539\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__20542\,
            I => \N__20536\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__20539\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__2254\ : Odrv4
    port map (
            O => \N__20536\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__2253\ : InMux
    port map (
            O => \N__20531\,
            I => \N__20528\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__20528\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\
        );

    \I__2251\ : InMux
    port map (
            O => \N__20525\,
            I => \N__20521\
        );

    \I__2250\ : InMux
    port map (
            O => \N__20524\,
            I => \N__20517\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__20521\,
            I => \N__20514\
        );

    \I__2248\ : InMux
    port map (
            O => \N__20520\,
            I => \N__20511\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__20517\,
            I => \N__20508\
        );

    \I__2246\ : Span12Mux_s3_h
    port map (
            O => \N__20514\,
            I => \N__20503\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__20511\,
            I => \N__20503\
        );

    \I__2244\ : Odrv4
    port map (
            O => \N__20508\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2243\ : Odrv12
    port map (
            O => \N__20503\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2242\ : CascadeMux
    port map (
            O => \N__20498\,
            I => \N__20495\
        );

    \I__2241\ : InMux
    port map (
            O => \N__20495\,
            I => \N__20492\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__20492\,
            I => \N__20488\
        );

    \I__2239\ : InMux
    port map (
            O => \N__20491\,
            I => \N__20485\
        );

    \I__2238\ : Span4Mux_s3_h
    port map (
            O => \N__20488\,
            I => \N__20481\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__20485\,
            I => \N__20478\
        );

    \I__2236\ : InMux
    port map (
            O => \N__20484\,
            I => \N__20475\
        );

    \I__2235\ : Span4Mux_v
    port map (
            O => \N__20481\,
            I => \N__20472\
        );

    \I__2234\ : Span4Mux_v
    port map (
            O => \N__20478\,
            I => \N__20467\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__20475\,
            I => \N__20467\
        );

    \I__2232\ : Odrv4
    port map (
            O => \N__20472\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__2231\ : Odrv4
    port map (
            O => \N__20467\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__2230\ : InMux
    port map (
            O => \N__20462\,
            I => \N__20458\
        );

    \I__2229\ : CascadeMux
    port map (
            O => \N__20461\,
            I => \N__20454\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__20458\,
            I => \N__20451\
        );

    \I__2227\ : InMux
    port map (
            O => \N__20457\,
            I => \N__20448\
        );

    \I__2226\ : InMux
    port map (
            O => \N__20454\,
            I => \N__20445\
        );

    \I__2225\ : Span12Mux_v
    port map (
            O => \N__20451\,
            I => \N__20442\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__20448\,
            I => \N__20439\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__20445\,
            I => \N__20436\
        );

    \I__2222\ : Odrv12
    port map (
            O => \N__20442\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2221\ : Odrv12
    port map (
            O => \N__20439\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2220\ : Odrv4
    port map (
            O => \N__20436\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2219\ : InMux
    port map (
            O => \N__20429\,
            I => \N__20426\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__20426\,
            I => \N__20422\
        );

    \I__2217\ : InMux
    port map (
            O => \N__20425\,
            I => \N__20419\
        );

    \I__2216\ : Span4Mux_h
    port map (
            O => \N__20422\,
            I => \N__20415\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__20419\,
            I => \N__20412\
        );

    \I__2214\ : InMux
    port map (
            O => \N__20418\,
            I => \N__20409\
        );

    \I__2213\ : Span4Mux_v
    port map (
            O => \N__20415\,
            I => \N__20406\
        );

    \I__2212\ : Span4Mux_v
    port map (
            O => \N__20412\,
            I => \N__20401\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__20409\,
            I => \N__20401\
        );

    \I__2210\ : Odrv4
    port map (
            O => \N__20406\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__2209\ : Odrv4
    port map (
            O => \N__20401\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__2208\ : CascadeMux
    port map (
            O => \N__20396\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_\
        );

    \I__2207\ : InMux
    port map (
            O => \N__20393\,
            I => \N__20390\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__20390\,
            I => \N__20387\
        );

    \I__2205\ : Span4Mux_s3_h
    port map (
            O => \N__20387\,
            I => \N__20383\
        );

    \I__2204\ : InMux
    port map (
            O => \N__20386\,
            I => \N__20380\
        );

    \I__2203\ : Span4Mux_v
    port map (
            O => \N__20383\,
            I => \N__20376\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__20380\,
            I => \N__20373\
        );

    \I__2201\ : InMux
    port map (
            O => \N__20379\,
            I => \N__20370\
        );

    \I__2200\ : Odrv4
    port map (
            O => \N__20376\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2199\ : Odrv12
    port map (
            O => \N__20373\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__20370\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2197\ : CascadeMux
    port map (
            O => \N__20363\,
            I => \N__20360\
        );

    \I__2196\ : InMux
    port map (
            O => \N__20360\,
            I => \N__20357\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__20357\,
            I => \N__20353\
        );

    \I__2194\ : CascadeMux
    port map (
            O => \N__20356\,
            I => \N__20350\
        );

    \I__2193\ : Span4Mux_v
    port map (
            O => \N__20353\,
            I => \N__20347\
        );

    \I__2192\ : InMux
    port map (
            O => \N__20350\,
            I => \N__20344\
        );

    \I__2191\ : Odrv4
    port map (
            O => \N__20347\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__20344\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__2189\ : InMux
    port map (
            O => \N__20339\,
            I => \N__20335\
        );

    \I__2188\ : InMux
    port map (
            O => \N__20338\,
            I => \N__20332\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__20335\,
            I => \N__20329\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__20332\,
            I => \N__20325\
        );

    \I__2185\ : Span4Mux_h
    port map (
            O => \N__20329\,
            I => \N__20322\
        );

    \I__2184\ : InMux
    port map (
            O => \N__20328\,
            I => \N__20319\
        );

    \I__2183\ : Span4Mux_s1_h
    port map (
            O => \N__20325\,
            I => \N__20316\
        );

    \I__2182\ : Odrv4
    port map (
            O => \N__20322\,
            I => pwm_duty_input_3
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__20319\,
            I => pwm_duty_input_3
        );

    \I__2180\ : Odrv4
    port map (
            O => \N__20316\,
            I => pwm_duty_input_3
        );

    \I__2179\ : InMux
    port map (
            O => \N__20309\,
            I => \N__20305\
        );

    \I__2178\ : InMux
    port map (
            O => \N__20308\,
            I => \N__20301\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__20305\,
            I => \N__20298\
        );

    \I__2176\ : InMux
    port map (
            O => \N__20304\,
            I => \N__20295\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__20301\,
            I => \N__20290\
        );

    \I__2174\ : Span4Mux_v
    port map (
            O => \N__20298\,
            I => \N__20290\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__20295\,
            I => pwm_duty_input_4
        );

    \I__2172\ : Odrv4
    port map (
            O => \N__20290\,
            I => pwm_duty_input_4
        );

    \I__2171\ : CascadeMux
    port map (
            O => \N__20285\,
            I => \N__20282\
        );

    \I__2170\ : InMux
    port map (
            O => \N__20282\,
            I => \N__20278\
        );

    \I__2169\ : InMux
    port map (
            O => \N__20281\,
            I => \N__20274\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__20278\,
            I => \N__20271\
        );

    \I__2167\ : InMux
    port map (
            O => \N__20277\,
            I => \N__20268\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__20274\,
            I => \N__20265\
        );

    \I__2165\ : Odrv4
    port map (
            O => \N__20271\,
            I => pwm_duty_input_5
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__20268\,
            I => pwm_duty_input_5
        );

    \I__2163\ : Odrv4
    port map (
            O => \N__20265\,
            I => pwm_duty_input_5
        );

    \I__2162\ : InMux
    port map (
            O => \N__20258\,
            I => \N__20255\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__20255\,
            I => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\
        );

    \I__2160\ : InMux
    port map (
            O => \N__20252\,
            I => \N__20248\
        );

    \I__2159\ : InMux
    port map (
            O => \N__20251\,
            I => \N__20245\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__20248\,
            I => \N__20242\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__20245\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__2156\ : Odrv4
    port map (
            O => \N__20242\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__2155\ : InMux
    port map (
            O => \N__20237\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\
        );

    \I__2154\ : CascadeMux
    port map (
            O => \N__20234\,
            I => \N__20230\
        );

    \I__2153\ : InMux
    port map (
            O => \N__20233\,
            I => \N__20225\
        );

    \I__2152\ : InMux
    port map (
            O => \N__20230\,
            I => \N__20225\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__20225\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__2150\ : InMux
    port map (
            O => \N__20222\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\
        );

    \I__2149\ : InMux
    port map (
            O => \N__20219\,
            I => \N__20213\
        );

    \I__2148\ : InMux
    port map (
            O => \N__20218\,
            I => \N__20213\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__20213\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__2146\ : InMux
    port map (
            O => \N__20210\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\
        );

    \I__2145\ : InMux
    port map (
            O => \N__20207\,
            I => \N__20201\
        );

    \I__2144\ : InMux
    port map (
            O => \N__20206\,
            I => \N__20201\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__20201\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__2142\ : InMux
    port map (
            O => \N__20198\,
            I => \bfn_3_20_0_\
        );

    \I__2141\ : InMux
    port map (
            O => \N__20195\,
            I => \N__20189\
        );

    \I__2140\ : InMux
    port map (
            O => \N__20194\,
            I => \N__20189\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__20189\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__2138\ : InMux
    port map (
            O => \N__20186\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\
        );

    \I__2137\ : InMux
    port map (
            O => \N__20183\,
            I => \N__20177\
        );

    \I__2136\ : InMux
    port map (
            O => \N__20182\,
            I => \N__20177\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__20177\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__2134\ : InMux
    port map (
            O => \N__20174\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\
        );

    \I__2133\ : InMux
    port map (
            O => \N__20171\,
            I => \N__20167\
        );

    \I__2132\ : InMux
    port map (
            O => \N__20170\,
            I => \N__20164\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__20167\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__20164\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__2129\ : InMux
    port map (
            O => \N__20159\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\
        );

    \I__2128\ : InMux
    port map (
            O => \N__20156\,
            I => \N__20150\
        );

    \I__2127\ : InMux
    port map (
            O => \N__20155\,
            I => \N__20150\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__20150\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__2125\ : InMux
    port map (
            O => \N__20147\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\
        );

    \I__2124\ : InMux
    port map (
            O => \N__20144\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\
        );

    \I__2123\ : InMux
    port map (
            O => \N__20141\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\
        );

    \I__2122\ : InMux
    port map (
            O => \N__20138\,
            I => \N__20134\
        );

    \I__2121\ : InMux
    port map (
            O => \N__20137\,
            I => \N__20131\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__20134\,
            I => \N__20128\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__20131\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__2118\ : Odrv4
    port map (
            O => \N__20128\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__2117\ : InMux
    port map (
            O => \N__20123\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\
        );

    \I__2116\ : CascadeMux
    port map (
            O => \N__20120\,
            I => \N__20117\
        );

    \I__2115\ : InMux
    port map (
            O => \N__20117\,
            I => \N__20113\
        );

    \I__2114\ : CascadeMux
    port map (
            O => \N__20116\,
            I => \N__20110\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__20113\,
            I => \N__20107\
        );

    \I__2112\ : InMux
    port map (
            O => \N__20110\,
            I => \N__20104\
        );

    \I__2111\ : Odrv4
    port map (
            O => \N__20107\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__20104\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__2109\ : InMux
    port map (
            O => \N__20099\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\
        );

    \I__2108\ : InMux
    port map (
            O => \N__20096\,
            I => \N__20090\
        );

    \I__2107\ : InMux
    port map (
            O => \N__20095\,
            I => \N__20090\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__20090\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__2105\ : InMux
    port map (
            O => \N__20087\,
            I => \bfn_3_19_0_\
        );

    \I__2104\ : InMux
    port map (
            O => \N__20084\,
            I => \N__20078\
        );

    \I__2103\ : InMux
    port map (
            O => \N__20083\,
            I => \N__20078\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__20078\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__2101\ : InMux
    port map (
            O => \N__20075\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\
        );

    \I__2100\ : InMux
    port map (
            O => \N__20072\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\
        );

    \I__2099\ : InMux
    port map (
            O => \N__20069\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\
        );

    \I__2098\ : InMux
    port map (
            O => \N__20066\,
            I => \N__20062\
        );

    \I__2097\ : InMux
    port map (
            O => \N__20065\,
            I => \N__20059\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__20062\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__20059\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__2094\ : InMux
    port map (
            O => \N__20054\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\
        );

    \I__2093\ : InMux
    port map (
            O => \N__20051\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\
        );

    \I__2092\ : InMux
    port map (
            O => \N__20048\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\
        );

    \I__2091\ : InMux
    port map (
            O => \N__20045\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\
        );

    \I__2090\ : InMux
    port map (
            O => \N__20042\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\
        );

    \I__2089\ : InMux
    port map (
            O => \N__20039\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\
        );

    \I__2088\ : InMux
    port map (
            O => \N__20036\,
            I => \bfn_3_18_0_\
        );

    \I__2087\ : InMux
    port map (
            O => \N__20033\,
            I => \N__20027\
        );

    \I__2086\ : InMux
    port map (
            O => \N__20032\,
            I => \N__20027\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__20027\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__2084\ : InMux
    port map (
            O => \N__20024\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\
        );

    \I__2083\ : InMux
    port map (
            O => \N__20021\,
            I => \N__20018\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__20018\,
            I => \N__20014\
        );

    \I__2081\ : InMux
    port map (
            O => \N__20017\,
            I => \N__20011\
        );

    \I__2080\ : Odrv4
    port map (
            O => \N__20014\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__20011\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__2078\ : InMux
    port map (
            O => \N__20006\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\
        );

    \I__2077\ : CascadeMux
    port map (
            O => \N__20003\,
            I => \N__20000\
        );

    \I__2076\ : InMux
    port map (
            O => \N__20000\,
            I => \N__19997\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__19997\,
            I => \N__19993\
        );

    \I__2074\ : InMux
    port map (
            O => \N__19996\,
            I => \N__19990\
        );

    \I__2073\ : Odrv4
    port map (
            O => \N__19993\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__19990\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__2071\ : InMux
    port map (
            O => \N__19985\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\
        );

    \I__2070\ : InMux
    port map (
            O => \N__19982\,
            I => \N__19979\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__19979\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\
        );

    \I__2068\ : CascadeMux
    port map (
            O => \N__19976\,
            I => \N__19973\
        );

    \I__2067\ : InMux
    port map (
            O => \N__19973\,
            I => \N__19970\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__19970\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\
        );

    \I__2065\ : InMux
    port map (
            O => \N__19967\,
            I => \N__19964\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__19964\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\
        );

    \I__2063\ : InMux
    port map (
            O => \N__19961\,
            I => \N__19958\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__19958\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\
        );

    \I__2061\ : CascadeMux
    port map (
            O => \N__19955\,
            I => \N__19952\
        );

    \I__2060\ : InMux
    port map (
            O => \N__19952\,
            I => \N__19949\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__19949\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\
        );

    \I__2058\ : CascadeMux
    port map (
            O => \N__19946\,
            I => \N__19943\
        );

    \I__2057\ : InMux
    port map (
            O => \N__19943\,
            I => \N__19940\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__19940\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\
        );

    \I__2055\ : InMux
    port map (
            O => \N__19937\,
            I => \N__19934\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__19934\,
            I => \N__19931\
        );

    \I__2053\ : Span4Mux_s3_h
    port map (
            O => \N__19931\,
            I => \N__19928\
        );

    \I__2052\ : Span4Mux_v
    port map (
            O => \N__19928\,
            I => \N__19925\
        );

    \I__2051\ : Odrv4
    port map (
            O => \N__19925\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\
        );

    \I__2050\ : InMux
    port map (
            O => \N__19922\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\
        );

    \I__2049\ : InMux
    port map (
            O => \N__19919\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\
        );

    \I__2048\ : CascadeMux
    port map (
            O => \N__19916\,
            I => \N__19913\
        );

    \I__2047\ : InMux
    port map (
            O => \N__19913\,
            I => \N__19910\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__19910\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\
        );

    \I__2045\ : CascadeMux
    port map (
            O => \N__19907\,
            I => \N__19904\
        );

    \I__2044\ : InMux
    port map (
            O => \N__19904\,
            I => \N__19901\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__19901\,
            I => \N__19897\
        );

    \I__2042\ : CascadeMux
    port map (
            O => \N__19900\,
            I => \N__19894\
        );

    \I__2041\ : Span4Mux_v
    port map (
            O => \N__19897\,
            I => \N__19891\
        );

    \I__2040\ : InMux
    port map (
            O => \N__19894\,
            I => \N__19888\
        );

    \I__2039\ : Sp12to4
    port map (
            O => \N__19891\,
            I => \N__19883\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__19888\,
            I => \N__19883\
        );

    \I__2037\ : Span12Mux_h
    port map (
            O => \N__19883\,
            I => \N__19880\
        );

    \I__2036\ : Odrv12
    port map (
            O => \N__19880\,
            I => \current_shift_inst.PI_CTRL.un1_integrator\
        );

    \I__2035\ : CascadeMux
    port map (
            O => \N__19877\,
            I => \N__19874\
        );

    \I__2034\ : InMux
    port map (
            O => \N__19874\,
            I => \N__19871\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__19871\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\
        );

    \I__2032\ : CascadeMux
    port map (
            O => \N__19868\,
            I => \N__19865\
        );

    \I__2031\ : InMux
    port map (
            O => \N__19865\,
            I => \N__19862\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__19862\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\
        );

    \I__2029\ : InMux
    port map (
            O => \N__19859\,
            I => \N__19856\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__19856\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\
        );

    \I__2027\ : CascadeMux
    port map (
            O => \N__19853\,
            I => \N__19850\
        );

    \I__2026\ : InMux
    port map (
            O => \N__19850\,
            I => \N__19847\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__19847\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\
        );

    \I__2024\ : InMux
    port map (
            O => \N__19844\,
            I => \N__19841\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__19841\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\
        );

    \I__2022\ : CascadeMux
    port map (
            O => \N__19838\,
            I => \N__19835\
        );

    \I__2021\ : InMux
    port map (
            O => \N__19835\,
            I => \N__19832\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__19832\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\
        );

    \I__2019\ : InMux
    port map (
            O => \N__19829\,
            I => \N__19826\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__19826\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\
        );

    \I__2017\ : CascadeMux
    port map (
            O => \N__19823\,
            I => \N__19819\
        );

    \I__2016\ : CascadeMux
    port map (
            O => \N__19822\,
            I => \N__19815\
        );

    \I__2015\ : InMux
    port map (
            O => \N__19819\,
            I => \N__19810\
        );

    \I__2014\ : InMux
    port map (
            O => \N__19818\,
            I => \N__19810\
        );

    \I__2013\ : InMux
    port map (
            O => \N__19815\,
            I => \N__19804\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__19810\,
            I => \N__19800\
        );

    \I__2011\ : InMux
    port map (
            O => \N__19809\,
            I => \N__19791\
        );

    \I__2010\ : InMux
    port map (
            O => \N__19808\,
            I => \N__19791\
        );

    \I__2009\ : InMux
    port map (
            O => \N__19807\,
            I => \N__19791\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__19804\,
            I => \N__19788\
        );

    \I__2007\ : InMux
    port map (
            O => \N__19803\,
            I => \N__19785\
        );

    \I__2006\ : Span4Mux_v
    port map (
            O => \N__19800\,
            I => \N__19782\
        );

    \I__2005\ : InMux
    port map (
            O => \N__19799\,
            I => \N__19779\
        );

    \I__2004\ : InMux
    port map (
            O => \N__19798\,
            I => \N__19776\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__19791\,
            I => \N__19769\
        );

    \I__2002\ : Span4Mux_v
    port map (
            O => \N__19788\,
            I => \N__19769\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__19785\,
            I => \N__19769\
        );

    \I__2000\ : Odrv4
    port map (
            O => \N__19782\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__19779\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__19776\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\
        );

    \I__1997\ : Odrv4
    port map (
            O => \N__19769\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\
        );

    \I__1996\ : CascadeMux
    port map (
            O => \N__19760\,
            I => \current_shift_inst.PI_CTRL.N_96_cascade_\
        );

    \I__1995\ : InMux
    port map (
            O => \N__19757\,
            I => \N__19753\
        );

    \I__1994\ : InMux
    port map (
            O => \N__19756\,
            I => \N__19750\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__19753\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__19750\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\
        );

    \I__1991\ : CascadeMux
    port map (
            O => \N__19745\,
            I => \N__19741\
        );

    \I__1990\ : CascadeMux
    port map (
            O => \N__19744\,
            I => \N__19738\
        );

    \I__1989\ : InMux
    port map (
            O => \N__19741\,
            I => \N__19732\
        );

    \I__1988\ : InMux
    port map (
            O => \N__19738\,
            I => \N__19732\
        );

    \I__1987\ : CascadeMux
    port map (
            O => \N__19737\,
            I => \N__19729\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__19732\,
            I => \N__19726\
        );

    \I__1985\ : InMux
    port map (
            O => \N__19729\,
            I => \N__19723\
        );

    \I__1984\ : Odrv4
    port map (
            O => \N__19726\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_3\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__19723\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_3\
        );

    \I__1982\ : InMux
    port map (
            O => \N__19718\,
            I => \N__19715\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__19715\,
            I => \N__19711\
        );

    \I__1980\ : InMux
    port map (
            O => \N__19714\,
            I => \N__19708\
        );

    \I__1979\ : Span4Mux_s1_h
    port map (
            O => \N__19711\,
            I => \N__19705\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__19708\,
            I => pwm_duty_input_0
        );

    \I__1977\ : Odrv4
    port map (
            O => \N__19705\,
            I => pwm_duty_input_0
        );

    \I__1976\ : InMux
    port map (
            O => \N__19700\,
            I => \N__19696\
        );

    \I__1975\ : InMux
    port map (
            O => \N__19699\,
            I => \N__19693\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__19696\,
            I => \N__19690\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__19693\,
            I => pwm_duty_input_1
        );

    \I__1972\ : Odrv4
    port map (
            O => \N__19690\,
            I => pwm_duty_input_1
        );

    \I__1971\ : InMux
    port map (
            O => \N__19685\,
            I => \N__19682\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__19682\,
            I => \N__19678\
        );

    \I__1969\ : InMux
    port map (
            O => \N__19681\,
            I => \N__19675\
        );

    \I__1968\ : Span4Mux_s1_h
    port map (
            O => \N__19678\,
            I => \N__19672\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__19675\,
            I => pwm_duty_input_2
        );

    \I__1966\ : Odrv4
    port map (
            O => \N__19672\,
            I => pwm_duty_input_2
        );

    \I__1965\ : CascadeMux
    port map (
            O => \N__19667\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\
        );

    \I__1964\ : InMux
    port map (
            O => \N__19664\,
            I => \N__19661\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__19661\,
            I => \pwm_generator_inst.un1_duty_inputlt3\
        );

    \I__1962\ : CascadeMux
    port map (
            O => \N__19658\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_\
        );

    \I__1961\ : InMux
    port map (
            O => \N__19655\,
            I => \N__19650\
        );

    \I__1960\ : InMux
    port map (
            O => \N__19654\,
            I => \N__19645\
        );

    \I__1959\ : InMux
    port map (
            O => \N__19653\,
            I => \N__19645\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__19650\,
            I => \N__19642\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__19645\,
            I => pwm_duty_input_9
        );

    \I__1956\ : Odrv4
    port map (
            O => \N__19642\,
            I => pwm_duty_input_9
        );

    \I__1955\ : InMux
    port map (
            O => \N__19637\,
            I => \N__19632\
        );

    \I__1954\ : InMux
    port map (
            O => \N__19636\,
            I => \N__19627\
        );

    \I__1953\ : InMux
    port map (
            O => \N__19635\,
            I => \N__19627\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__19632\,
            I => \N__19624\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__19627\,
            I => pwm_duty_input_7
        );

    \I__1950\ : Odrv4
    port map (
            O => \N__19624\,
            I => pwm_duty_input_7
        );

    \I__1949\ : CascadeMux
    port map (
            O => \N__19619\,
            I => \N__19614\
        );

    \I__1948\ : InMux
    port map (
            O => \N__19618\,
            I => \N__19611\
        );

    \I__1947\ : InMux
    port map (
            O => \N__19617\,
            I => \N__19608\
        );

    \I__1946\ : InMux
    port map (
            O => \N__19614\,
            I => \N__19605\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__19611\,
            I => \N__19602\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__19608\,
            I => pwm_duty_input_6
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__19605\,
            I => pwm_duty_input_6
        );

    \I__1942\ : Odrv4
    port map (
            O => \N__19602\,
            I => pwm_duty_input_6
        );

    \I__1941\ : InMux
    port map (
            O => \N__19595\,
            I => \N__19590\
        );

    \I__1940\ : InMux
    port map (
            O => \N__19594\,
            I => \N__19587\
        );

    \I__1939\ : InMux
    port map (
            O => \N__19593\,
            I => \N__19584\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__19590\,
            I => pwm_duty_input_8
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__19587\,
            I => pwm_duty_input_8
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__19584\,
            I => pwm_duty_input_8
        );

    \I__1935\ : CascadeMux
    port map (
            O => \N__19577\,
            I => \N__19574\
        );

    \I__1934\ : InMux
    port map (
            O => \N__19574\,
            I => \N__19571\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__19571\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\
        );

    \I__1932\ : CascadeMux
    port map (
            O => \N__19568\,
            I => \N__19565\
        );

    \I__1931\ : InMux
    port map (
            O => \N__19565\,
            I => \N__19562\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__19562\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\
        );

    \I__1929\ : CascadeMux
    port map (
            O => \N__19559\,
            I => \N__19556\
        );

    \I__1928\ : InMux
    port map (
            O => \N__19556\,
            I => \N__19553\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__19553\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\
        );

    \I__1926\ : InMux
    port map (
            O => \N__19550\,
            I => \N__19547\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__19547\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\
        );

    \I__1924\ : InMux
    port map (
            O => \N__19544\,
            I => \N__19541\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__19541\,
            I => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0\
        );

    \I__1922\ : CascadeMux
    port map (
            O => \N__19538\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\
        );

    \I__1921\ : InMux
    port map (
            O => \N__19535\,
            I => \N__19532\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__19532\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\
        );

    \I__1919\ : CascadeMux
    port map (
            O => \N__19529\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_\
        );

    \I__1918\ : InMux
    port map (
            O => \N__19526\,
            I => \N__19523\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__19523\,
            I => \N__19520\
        );

    \I__1916\ : Odrv4
    port map (
            O => \N__19520\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\
        );

    \I__1915\ : InMux
    port map (
            O => \N__19517\,
            I => \N__19514\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__19514\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\
        );

    \I__1913\ : InMux
    port map (
            O => \N__19511\,
            I => \N__19504\
        );

    \I__1912\ : InMux
    port map (
            O => \N__19510\,
            I => \N__19504\
        );

    \I__1911\ : InMux
    port map (
            O => \N__19509\,
            I => \N__19501\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__19504\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__19501\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__1908\ : CascadeMux
    port map (
            O => \N__19496\,
            I => \N__19491\
        );

    \I__1907\ : InMux
    port map (
            O => \N__19495\,
            I => \N__19485\
        );

    \I__1906\ : InMux
    port map (
            O => \N__19494\,
            I => \N__19482\
        );

    \I__1905\ : InMux
    port map (
            O => \N__19491\,
            I => \N__19475\
        );

    \I__1904\ : InMux
    port map (
            O => \N__19490\,
            I => \N__19475\
        );

    \I__1903\ : InMux
    port map (
            O => \N__19489\,
            I => \N__19475\
        );

    \I__1902\ : CascadeMux
    port map (
            O => \N__19488\,
            I => \N__19472\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__19485\,
            I => \N__19465\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__19482\,
            I => \N__19465\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__19475\,
            I => \N__19465\
        );

    \I__1898\ : InMux
    port map (
            O => \N__19472\,
            I => \N__19461\
        );

    \I__1897\ : Span4Mux_v
    port map (
            O => \N__19465\,
            I => \N__19458\
        );

    \I__1896\ : InMux
    port map (
            O => \N__19464\,
            I => \N__19455\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__19461\,
            I => \current_shift_inst.PI_CTRL.N_159\
        );

    \I__1894\ : Odrv4
    port map (
            O => \N__19458\,
            I => \current_shift_inst.PI_CTRL.N_159\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__19455\,
            I => \current_shift_inst.PI_CTRL.N_159\
        );

    \I__1892\ : InMux
    port map (
            O => \N__19448\,
            I => \N__19436\
        );

    \I__1891\ : InMux
    port map (
            O => \N__19447\,
            I => \N__19436\
        );

    \I__1890\ : InMux
    port map (
            O => \N__19446\,
            I => \N__19436\
        );

    \I__1889\ : InMux
    port map (
            O => \N__19445\,
            I => \N__19436\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__19436\,
            I => \current_shift_inst.PI_CTRL.N_96\
        );

    \I__1887\ : CascadeMux
    port map (
            O => \N__19433\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\
        );

    \I__1886\ : InMux
    port map (
            O => \N__19430\,
            I => \N__19427\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__19427\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\
        );

    \I__1884\ : InMux
    port map (
            O => \N__19424\,
            I => \N__19421\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__19421\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\
        );

    \I__1882\ : CascadeMux
    port map (
            O => \N__19418\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_\
        );

    \I__1881\ : InMux
    port map (
            O => \N__19415\,
            I => \N__19412\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__19412\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\
        );

    \I__1879\ : CascadeMux
    port map (
            O => \N__19409\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_\
        );

    \I__1878\ : InMux
    port map (
            O => \N__19406\,
            I => \N__19403\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__19403\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\
        );

    \I__1876\ : CascadeMux
    port map (
            O => \N__19400\,
            I => \N__19397\
        );

    \I__1875\ : InMux
    port map (
            O => \N__19397\,
            I => \N__19394\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__19394\,
            I => \N__19391\
        );

    \I__1873\ : Span4Mux_v
    port map (
            O => \N__19391\,
            I => \N__19388\
        );

    \I__1872\ : Odrv4
    port map (
            O => \N__19388\,
            I => \current_shift_inst.PI_CTRL.integrator_1_26\
        );

    \I__1871\ : InMux
    port map (
            O => \N__19385\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\
        );

    \I__1870\ : CascadeMux
    port map (
            O => \N__19382\,
            I => \N__19379\
        );

    \I__1869\ : InMux
    port map (
            O => \N__19379\,
            I => \N__19376\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__19376\,
            I => \N__19373\
        );

    \I__1867\ : Span4Mux_v
    port map (
            O => \N__19373\,
            I => \N__19370\
        );

    \I__1866\ : Odrv4
    port map (
            O => \N__19370\,
            I => \current_shift_inst.PI_CTRL.integrator_1_27\
        );

    \I__1865\ : InMux
    port map (
            O => \N__19367\,
            I => \N__19364\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__19364\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\
        );

    \I__1863\ : InMux
    port map (
            O => \N__19361\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\
        );

    \I__1862\ : CascadeMux
    port map (
            O => \N__19358\,
            I => \N__19355\
        );

    \I__1861\ : InMux
    port map (
            O => \N__19355\,
            I => \N__19352\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__19352\,
            I => \N__19349\
        );

    \I__1859\ : Span4Mux_h
    port map (
            O => \N__19349\,
            I => \N__19346\
        );

    \I__1858\ : Odrv4
    port map (
            O => \N__19346\,
            I => \current_shift_inst.PI_CTRL.integrator_1_28\
        );

    \I__1857\ : InMux
    port map (
            O => \N__19343\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\
        );

    \I__1856\ : CascadeMux
    port map (
            O => \N__19340\,
            I => \N__19337\
        );

    \I__1855\ : InMux
    port map (
            O => \N__19337\,
            I => \N__19334\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__19334\,
            I => \N__19331\
        );

    \I__1853\ : Odrv4
    port map (
            O => \N__19331\,
            I => \current_shift_inst.PI_CTRL.integrator_1_29\
        );

    \I__1852\ : InMux
    port map (
            O => \N__19328\,
            I => \N__19325\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__19325\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\
        );

    \I__1850\ : InMux
    port map (
            O => \N__19322\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\
        );

    \I__1849\ : CascadeMux
    port map (
            O => \N__19319\,
            I => \N__19316\
        );

    \I__1848\ : InMux
    port map (
            O => \N__19316\,
            I => \N__19313\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__19313\,
            I => \N__19310\
        );

    \I__1846\ : Odrv4
    port map (
            O => \N__19310\,
            I => \current_shift_inst.PI_CTRL.integrator_1_30\
        );

    \I__1845\ : InMux
    port map (
            O => \N__19307\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\
        );

    \I__1844\ : InMux
    port map (
            O => \N__19304\,
            I => \N__19301\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__19301\,
            I => \N__19298\
        );

    \I__1842\ : Odrv4
    port map (
            O => \N__19298\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\
        );

    \I__1841\ : CascadeMux
    port map (
            O => \N__19295\,
            I => \N__19292\
        );

    \I__1840\ : InMux
    port map (
            O => \N__19292\,
            I => \N__19289\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__19289\,
            I => \N__19286\
        );

    \I__1838\ : Span4Mux_v
    port map (
            O => \N__19286\,
            I => \N__19283\
        );

    \I__1837\ : Odrv4
    port map (
            O => \N__19283\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30\
        );

    \I__1836\ : InMux
    port map (
            O => \N__19280\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\
        );

    \I__1835\ : InMux
    port map (
            O => \N__19277\,
            I => \N__19274\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__19274\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\
        );

    \I__1833\ : InMux
    port map (
            O => \N__19271\,
            I => \N__19268\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__19268\,
            I => \N__19265\
        );

    \I__1831\ : Span4Mux_v
    port map (
            O => \N__19265\,
            I => \N__19262\
        );

    \I__1830\ : Odrv4
    port map (
            O => \N__19262\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\
        );

    \I__1829\ : CascadeMux
    port map (
            O => \N__19259\,
            I => \N__19256\
        );

    \I__1828\ : InMux
    port map (
            O => \N__19256\,
            I => \N__19253\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__19253\,
            I => \N__19250\
        );

    \I__1826\ : Odrv4
    port map (
            O => \N__19250\,
            I => \current_shift_inst.PI_CTRL.integrator_1_18\
        );

    \I__1825\ : InMux
    port map (
            O => \N__19247\,
            I => \N__19244\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__19244\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\
        );

    \I__1823\ : InMux
    port map (
            O => \N__19241\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\
        );

    \I__1822\ : CascadeMux
    port map (
            O => \N__19238\,
            I => \N__19235\
        );

    \I__1821\ : InMux
    port map (
            O => \N__19235\,
            I => \N__19232\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__19232\,
            I => \N__19229\
        );

    \I__1819\ : Odrv4
    port map (
            O => \N__19229\,
            I => \current_shift_inst.PI_CTRL.integrator_1_19\
        );

    \I__1818\ : InMux
    port map (
            O => \N__19226\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\
        );

    \I__1817\ : CascadeMux
    port map (
            O => \N__19223\,
            I => \N__19220\
        );

    \I__1816\ : InMux
    port map (
            O => \N__19220\,
            I => \N__19217\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__19217\,
            I => \N__19214\
        );

    \I__1814\ : Odrv4
    port map (
            O => \N__19214\,
            I => \current_shift_inst.PI_CTRL.integrator_1_20\
        );

    \I__1813\ : InMux
    port map (
            O => \N__19211\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\
        );

    \I__1812\ : CascadeMux
    port map (
            O => \N__19208\,
            I => \N__19205\
        );

    \I__1811\ : InMux
    port map (
            O => \N__19205\,
            I => \N__19202\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__19202\,
            I => \N__19199\
        );

    \I__1809\ : Span4Mux_v
    port map (
            O => \N__19199\,
            I => \N__19196\
        );

    \I__1808\ : Odrv4
    port map (
            O => \N__19196\,
            I => \current_shift_inst.PI_CTRL.integrator_1_21\
        );

    \I__1807\ : InMux
    port map (
            O => \N__19193\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\
        );

    \I__1806\ : CascadeMux
    port map (
            O => \N__19190\,
            I => \N__19187\
        );

    \I__1805\ : InMux
    port map (
            O => \N__19187\,
            I => \N__19184\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__19184\,
            I => \N__19181\
        );

    \I__1803\ : Span4Mux_v
    port map (
            O => \N__19181\,
            I => \N__19178\
        );

    \I__1802\ : Odrv4
    port map (
            O => \N__19178\,
            I => \current_shift_inst.PI_CTRL.integrator_1_22\
        );

    \I__1801\ : InMux
    port map (
            O => \N__19175\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\
        );

    \I__1800\ : CascadeMux
    port map (
            O => \N__19172\,
            I => \N__19169\
        );

    \I__1799\ : InMux
    port map (
            O => \N__19169\,
            I => \N__19166\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__19166\,
            I => \N__19163\
        );

    \I__1797\ : Span4Mux_h
    port map (
            O => \N__19163\,
            I => \N__19160\
        );

    \I__1796\ : Odrv4
    port map (
            O => \N__19160\,
            I => \current_shift_inst.PI_CTRL.integrator_1_23\
        );

    \I__1795\ : InMux
    port map (
            O => \N__19157\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\
        );

    \I__1794\ : CascadeMux
    port map (
            O => \N__19154\,
            I => \N__19151\
        );

    \I__1793\ : InMux
    port map (
            O => \N__19151\,
            I => \N__19148\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__19148\,
            I => \current_shift_inst.PI_CTRL.integrator_1_24\
        );

    \I__1791\ : InMux
    port map (
            O => \N__19145\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\
        );

    \I__1790\ : CascadeMux
    port map (
            O => \N__19142\,
            I => \N__19139\
        );

    \I__1789\ : InMux
    port map (
            O => \N__19139\,
            I => \N__19136\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__19136\,
            I => \N__19133\
        );

    \I__1787\ : Span4Mux_h
    port map (
            O => \N__19133\,
            I => \N__19130\
        );

    \I__1786\ : Odrv4
    port map (
            O => \N__19130\,
            I => \current_shift_inst.PI_CTRL.integrator_1_25\
        );

    \I__1785\ : InMux
    port map (
            O => \N__19127\,
            I => \bfn_2_16_0_\
        );

    \I__1784\ : CascadeMux
    port map (
            O => \N__19124\,
            I => \N__19121\
        );

    \I__1783\ : InMux
    port map (
            O => \N__19121\,
            I => \N__19118\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__19118\,
            I => \N__19115\
        );

    \I__1781\ : Span4Mux_v
    port map (
            O => \N__19115\,
            I => \N__19112\
        );

    \I__1780\ : Span4Mux_v
    port map (
            O => \N__19112\,
            I => \N__19109\
        );

    \I__1779\ : Odrv4
    port map (
            O => \N__19109\,
            I => \current_shift_inst.PI_CTRL.integrator_1_10\
        );

    \I__1778\ : InMux
    port map (
            O => \N__19106\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\
        );

    \I__1777\ : CascadeMux
    port map (
            O => \N__19103\,
            I => \N__19100\
        );

    \I__1776\ : InMux
    port map (
            O => \N__19100\,
            I => \N__19097\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__19097\,
            I => \N__19094\
        );

    \I__1774\ : Span4Mux_v
    port map (
            O => \N__19094\,
            I => \N__19091\
        );

    \I__1773\ : Span4Mux_v
    port map (
            O => \N__19091\,
            I => \N__19088\
        );

    \I__1772\ : Odrv4
    port map (
            O => \N__19088\,
            I => \current_shift_inst.PI_CTRL.integrator_1_11\
        );

    \I__1771\ : InMux
    port map (
            O => \N__19085\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\
        );

    \I__1770\ : CascadeMux
    port map (
            O => \N__19082\,
            I => \N__19079\
        );

    \I__1769\ : InMux
    port map (
            O => \N__19079\,
            I => \N__19076\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__19076\,
            I => \N__19073\
        );

    \I__1767\ : Span4Mux_v
    port map (
            O => \N__19073\,
            I => \N__19070\
        );

    \I__1766\ : Span4Mux_v
    port map (
            O => \N__19070\,
            I => \N__19067\
        );

    \I__1765\ : Odrv4
    port map (
            O => \N__19067\,
            I => \current_shift_inst.PI_CTRL.integrator_1_12\
        );

    \I__1764\ : CascadeMux
    port map (
            O => \N__19064\,
            I => \N__19061\
        );

    \I__1763\ : InMux
    port map (
            O => \N__19061\,
            I => \N__19058\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__19058\,
            I => \N__19055\
        );

    \I__1761\ : Span4Mux_v
    port map (
            O => \N__19055\,
            I => \N__19052\
        );

    \I__1760\ : Odrv4
    port map (
            O => \N__19052\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\
        );

    \I__1759\ : InMux
    port map (
            O => \N__19049\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\
        );

    \I__1758\ : CascadeMux
    port map (
            O => \N__19046\,
            I => \N__19043\
        );

    \I__1757\ : InMux
    port map (
            O => \N__19043\,
            I => \N__19040\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__19040\,
            I => \N__19037\
        );

    \I__1755\ : Span4Mux_v
    port map (
            O => \N__19037\,
            I => \N__19034\
        );

    \I__1754\ : Span4Mux_v
    port map (
            O => \N__19034\,
            I => \N__19031\
        );

    \I__1753\ : Odrv4
    port map (
            O => \N__19031\,
            I => \current_shift_inst.PI_CTRL.integrator_1_13\
        );

    \I__1752\ : InMux
    port map (
            O => \N__19028\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\
        );

    \I__1751\ : CascadeMux
    port map (
            O => \N__19025\,
            I => \N__19022\
        );

    \I__1750\ : InMux
    port map (
            O => \N__19022\,
            I => \N__19019\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__19019\,
            I => \N__19016\
        );

    \I__1748\ : Span4Mux_v
    port map (
            O => \N__19016\,
            I => \N__19013\
        );

    \I__1747\ : Span4Mux_v
    port map (
            O => \N__19013\,
            I => \N__19010\
        );

    \I__1746\ : Odrv4
    port map (
            O => \N__19010\,
            I => \current_shift_inst.PI_CTRL.integrator_1_14\
        );

    \I__1745\ : InMux
    port map (
            O => \N__19007\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\
        );

    \I__1744\ : CascadeMux
    port map (
            O => \N__19004\,
            I => \N__19001\
        );

    \I__1743\ : InMux
    port map (
            O => \N__19001\,
            I => \N__18998\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__18998\,
            I => \N__18995\
        );

    \I__1741\ : Span4Mux_v
    port map (
            O => \N__18995\,
            I => \N__18992\
        );

    \I__1740\ : Span4Mux_v
    port map (
            O => \N__18992\,
            I => \N__18989\
        );

    \I__1739\ : Odrv4
    port map (
            O => \N__18989\,
            I => \current_shift_inst.PI_CTRL.integrator_1_15\
        );

    \I__1738\ : InMux
    port map (
            O => \N__18986\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\
        );

    \I__1737\ : CascadeMux
    port map (
            O => \N__18983\,
            I => \N__18980\
        );

    \I__1736\ : InMux
    port map (
            O => \N__18980\,
            I => \N__18977\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__18977\,
            I => \current_shift_inst.PI_CTRL.integrator_1_16\
        );

    \I__1734\ : InMux
    port map (
            O => \N__18974\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\
        );

    \I__1733\ : CascadeMux
    port map (
            O => \N__18971\,
            I => \N__18968\
        );

    \I__1732\ : InMux
    port map (
            O => \N__18968\,
            I => \N__18965\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__18965\,
            I => \N__18962\
        );

    \I__1730\ : Span4Mux_h
    port map (
            O => \N__18962\,
            I => \N__18959\
        );

    \I__1729\ : Odrv4
    port map (
            O => \N__18959\,
            I => \current_shift_inst.PI_CTRL.integrator_1_17\
        );

    \I__1728\ : InMux
    port map (
            O => \N__18956\,
            I => \bfn_2_15_0_\
        );

    \I__1727\ : CascadeMux
    port map (
            O => \N__18953\,
            I => \N__18950\
        );

    \I__1726\ : InMux
    port map (
            O => \N__18950\,
            I => \N__18947\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__18947\,
            I => \N__18944\
        );

    \I__1724\ : Span4Mux_v
    port map (
            O => \N__18944\,
            I => \N__18941\
        );

    \I__1723\ : Span4Mux_v
    port map (
            O => \N__18941\,
            I => \N__18938\
        );

    \I__1722\ : Odrv4
    port map (
            O => \N__18938\,
            I => \current_shift_inst.PI_CTRL.integrator_1_2\
        );

    \I__1721\ : InMux
    port map (
            O => \N__18935\,
            I => \N__18932\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__18932\,
            I => \N__18929\
        );

    \I__1719\ : Span4Mux_v
    port map (
            O => \N__18929\,
            I => \N__18926\
        );

    \I__1718\ : Odrv4
    port map (
            O => \N__18926\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\
        );

    \I__1717\ : InMux
    port map (
            O => \N__18923\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\
        );

    \I__1716\ : CascadeMux
    port map (
            O => \N__18920\,
            I => \N__18917\
        );

    \I__1715\ : InMux
    port map (
            O => \N__18917\,
            I => \N__18914\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__18914\,
            I => \N__18911\
        );

    \I__1713\ : Span4Mux_s3_h
    port map (
            O => \N__18911\,
            I => \N__18908\
        );

    \I__1712\ : Span4Mux_v
    port map (
            O => \N__18908\,
            I => \N__18905\
        );

    \I__1711\ : Span4Mux_v
    port map (
            O => \N__18905\,
            I => \N__18902\
        );

    \I__1710\ : Odrv4
    port map (
            O => \N__18902\,
            I => \current_shift_inst.PI_CTRL.integrator_1_3\
        );

    \I__1709\ : InMux
    port map (
            O => \N__18899\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\
        );

    \I__1708\ : CascadeMux
    port map (
            O => \N__18896\,
            I => \N__18893\
        );

    \I__1707\ : InMux
    port map (
            O => \N__18893\,
            I => \N__18890\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__18890\,
            I => \N__18887\
        );

    \I__1705\ : Span4Mux_v
    port map (
            O => \N__18887\,
            I => \N__18884\
        );

    \I__1704\ : Span4Mux_v
    port map (
            O => \N__18884\,
            I => \N__18881\
        );

    \I__1703\ : Odrv4
    port map (
            O => \N__18881\,
            I => \current_shift_inst.PI_CTRL.integrator_1_4\
        );

    \I__1702\ : CascadeMux
    port map (
            O => \N__18878\,
            I => \N__18875\
        );

    \I__1701\ : InMux
    port map (
            O => \N__18875\,
            I => \N__18872\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__18872\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\
        );

    \I__1699\ : InMux
    port map (
            O => \N__18869\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\
        );

    \I__1698\ : CascadeMux
    port map (
            O => \N__18866\,
            I => \N__18863\
        );

    \I__1697\ : InMux
    port map (
            O => \N__18863\,
            I => \N__18860\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__18860\,
            I => \N__18857\
        );

    \I__1695\ : Span4Mux_v
    port map (
            O => \N__18857\,
            I => \N__18854\
        );

    \I__1694\ : Span4Mux_v
    port map (
            O => \N__18854\,
            I => \N__18851\
        );

    \I__1693\ : Odrv4
    port map (
            O => \N__18851\,
            I => \current_shift_inst.PI_CTRL.integrator_1_5\
        );

    \I__1692\ : InMux
    port map (
            O => \N__18848\,
            I => \N__18845\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__18845\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\
        );

    \I__1690\ : InMux
    port map (
            O => \N__18842\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\
        );

    \I__1689\ : CascadeMux
    port map (
            O => \N__18839\,
            I => \N__18836\
        );

    \I__1688\ : InMux
    port map (
            O => \N__18836\,
            I => \N__18833\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__18833\,
            I => \N__18830\
        );

    \I__1686\ : Span4Mux_v
    port map (
            O => \N__18830\,
            I => \N__18827\
        );

    \I__1685\ : Span4Mux_v
    port map (
            O => \N__18827\,
            I => \N__18824\
        );

    \I__1684\ : Odrv4
    port map (
            O => \N__18824\,
            I => \current_shift_inst.PI_CTRL.integrator_1_6\
        );

    \I__1683\ : InMux
    port map (
            O => \N__18821\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\
        );

    \I__1682\ : CascadeMux
    port map (
            O => \N__18818\,
            I => \N__18815\
        );

    \I__1681\ : InMux
    port map (
            O => \N__18815\,
            I => \N__18812\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__18812\,
            I => \N__18809\
        );

    \I__1679\ : Span12Mux_v
    port map (
            O => \N__18809\,
            I => \N__18806\
        );

    \I__1678\ : Odrv12
    port map (
            O => \N__18806\,
            I => \current_shift_inst.PI_CTRL.integrator_1_7\
        );

    \I__1677\ : InMux
    port map (
            O => \N__18803\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\
        );

    \I__1676\ : CascadeMux
    port map (
            O => \N__18800\,
            I => \N__18797\
        );

    \I__1675\ : InMux
    port map (
            O => \N__18797\,
            I => \N__18794\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__18794\,
            I => \N__18791\
        );

    \I__1673\ : Span4Mux_v
    port map (
            O => \N__18791\,
            I => \N__18788\
        );

    \I__1672\ : Span4Mux_v
    port map (
            O => \N__18788\,
            I => \N__18785\
        );

    \I__1671\ : Odrv4
    port map (
            O => \N__18785\,
            I => \current_shift_inst.PI_CTRL.integrator_1_8\
        );

    \I__1670\ : InMux
    port map (
            O => \N__18782\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\
        );

    \I__1669\ : CascadeMux
    port map (
            O => \N__18779\,
            I => \N__18776\
        );

    \I__1668\ : InMux
    port map (
            O => \N__18776\,
            I => \N__18773\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__18773\,
            I => \N__18770\
        );

    \I__1666\ : Span12Mux_h
    port map (
            O => \N__18770\,
            I => \N__18767\
        );

    \I__1665\ : Odrv12
    port map (
            O => \N__18767\,
            I => \current_shift_inst.PI_CTRL.integrator_1_9\
        );

    \I__1664\ : InMux
    port map (
            O => \N__18764\,
            I => \bfn_2_14_0_\
        );

    \I__1663\ : InMux
    port map (
            O => \N__18761\,
            I => \N__18758\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__18758\,
            I => \N__18755\
        );

    \I__1661\ : Odrv4
    port map (
            O => \N__18755\,
            I => \current_shift_inst.PI_CTRL.N_91\
        );

    \I__1660\ : InMux
    port map (
            O => \N__18752\,
            I => \N__18749\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__18749\,
            I => \N_42_i_i\
        );

    \I__1658\ : InMux
    port map (
            O => \N__18746\,
            I => \N__18743\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__18743\,
            I => un7_start_stop_0_a2
        );

    \I__1656\ : InMux
    port map (
            O => \N__18740\,
            I => \N__18737\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__18737\,
            I => \N__18734\
        );

    \I__1654\ : Odrv4
    port map (
            O => \N__18734\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\
        );

    \I__1653\ : InMux
    port map (
            O => \N__18731\,
            I => \N__18722\
        );

    \I__1652\ : InMux
    port map (
            O => \N__18730\,
            I => \N__18722\
        );

    \I__1651\ : InMux
    port map (
            O => \N__18729\,
            I => \N__18722\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__18722\,
            I => \current_shift_inst.PI_CTRL.N_97\
        );

    \I__1649\ : InMux
    port map (
            O => \N__18719\,
            I => \N__18716\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__18716\,
            I => \N__18713\
        );

    \I__1647\ : Odrv4
    port map (
            O => \N__18713\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\
        );

    \I__1646\ : InMux
    port map (
            O => \N__18710\,
            I => \N__18707\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__18707\,
            I => \N__18704\
        );

    \I__1644\ : Odrv4
    port map (
            O => \N__18704\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_11\
        );

    \I__1643\ : InMux
    port map (
            O => \N__18701\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\
        );

    \I__1642\ : InMux
    port map (
            O => \N__18698\,
            I => \N__18695\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__18695\,
            I => \N__18692\
        );

    \I__1640\ : Odrv4
    port map (
            O => \N__18692\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_12\
        );

    \I__1639\ : InMux
    port map (
            O => \N__18689\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\
        );

    \I__1638\ : InMux
    port map (
            O => \N__18686\,
            I => \N__18683\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__18683\,
            I => \N__18680\
        );

    \I__1636\ : Odrv4
    port map (
            O => \N__18680\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_13\
        );

    \I__1635\ : InMux
    port map (
            O => \N__18677\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\
        );

    \I__1634\ : InMux
    port map (
            O => \N__18674\,
            I => \N__18671\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__18671\,
            I => \N__18668\
        );

    \I__1632\ : Span4Mux_h
    port map (
            O => \N__18668\,
            I => \N__18665\
        );

    \I__1631\ : Odrv4
    port map (
            O => \N__18665\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_14\
        );

    \I__1630\ : CascadeMux
    port map (
            O => \N__18662\,
            I => \N__18649\
        );

    \I__1629\ : CascadeMux
    port map (
            O => \N__18661\,
            I => \N__18646\
        );

    \I__1628\ : CascadeMux
    port map (
            O => \N__18660\,
            I => \N__18643\
        );

    \I__1627\ : CascadeMux
    port map (
            O => \N__18659\,
            I => \N__18640\
        );

    \I__1626\ : CascadeMux
    port map (
            O => \N__18658\,
            I => \N__18637\
        );

    \I__1625\ : CascadeMux
    port map (
            O => \N__18657\,
            I => \N__18634\
        );

    \I__1624\ : CascadeMux
    port map (
            O => \N__18656\,
            I => \N__18631\
        );

    \I__1623\ : CascadeMux
    port map (
            O => \N__18655\,
            I => \N__18628\
        );

    \I__1622\ : CascadeMux
    port map (
            O => \N__18654\,
            I => \N__18625\
        );

    \I__1621\ : CascadeMux
    port map (
            O => \N__18653\,
            I => \N__18622\
        );

    \I__1620\ : InMux
    port map (
            O => \N__18652\,
            I => \N__18618\
        );

    \I__1619\ : InMux
    port map (
            O => \N__18649\,
            I => \N__18609\
        );

    \I__1618\ : InMux
    port map (
            O => \N__18646\,
            I => \N__18609\
        );

    \I__1617\ : InMux
    port map (
            O => \N__18643\,
            I => \N__18609\
        );

    \I__1616\ : InMux
    port map (
            O => \N__18640\,
            I => \N__18609\
        );

    \I__1615\ : InMux
    port map (
            O => \N__18637\,
            I => \N__18606\
        );

    \I__1614\ : InMux
    port map (
            O => \N__18634\,
            I => \N__18599\
        );

    \I__1613\ : InMux
    port map (
            O => \N__18631\,
            I => \N__18599\
        );

    \I__1612\ : InMux
    port map (
            O => \N__18628\,
            I => \N__18599\
        );

    \I__1611\ : InMux
    port map (
            O => \N__18625\,
            I => \N__18592\
        );

    \I__1610\ : InMux
    port map (
            O => \N__18622\,
            I => \N__18592\
        );

    \I__1609\ : InMux
    port map (
            O => \N__18621\,
            I => \N__18592\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__18618\,
            I => \N__18585\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__18609\,
            I => \N__18585\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__18606\,
            I => \N__18585\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__18599\,
            I => \N__18580\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__18592\,
            I => \N__18580\
        );

    \I__1603\ : Span4Mux_v
    port map (
            O => \N__18585\,
            I => \N__18575\
        );

    \I__1602\ : Span4Mux_v
    port map (
            O => \N__18580\,
            I => \N__18575\
        );

    \I__1601\ : Odrv4
    port map (
            O => \N__18575\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_19\
        );

    \I__1600\ : InMux
    port map (
            O => \N__18572\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\
        );

    \I__1599\ : InMux
    port map (
            O => \N__18569\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\
        );

    \I__1598\ : InMux
    port map (
            O => \N__18566\,
            I => \N__18563\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__18563\,
            I => \N__18560\
        );

    \I__1596\ : Span4Mux_v
    port map (
            O => \N__18560\,
            I => \N__18557\
        );

    \I__1595\ : Odrv4
    port map (
            O => \N__18557\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_3\
        );

    \I__1594\ : CascadeMux
    port map (
            O => \N__18554\,
            I => \N__18551\
        );

    \I__1593\ : InMux
    port map (
            O => \N__18551\,
            I => \N__18548\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__18548\,
            I => \N__18545\
        );

    \I__1591\ : Span4Mux_v
    port map (
            O => \N__18545\,
            I => \N__18542\
        );

    \I__1590\ : Span4Mux_v
    port map (
            O => \N__18542\,
            I => \N__18539\
        );

    \I__1589\ : Odrv4
    port map (
            O => \N__18539\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_18\
        );

    \I__1588\ : InMux
    port map (
            O => \N__18536\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\
        );

    \I__1587\ : CascadeMux
    port map (
            O => \N__18533\,
            I => \N__18530\
        );

    \I__1586\ : InMux
    port map (
            O => \N__18530\,
            I => \N__18527\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__18527\,
            I => \N__18524\
        );

    \I__1584\ : Odrv4
    port map (
            O => \N__18524\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_4\
        );

    \I__1583\ : InMux
    port map (
            O => \N__18521\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\
        );

    \I__1582\ : InMux
    port map (
            O => \N__18518\,
            I => \N__18515\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__18515\,
            I => \N__18512\
        );

    \I__1580\ : Odrv4
    port map (
            O => \N__18512\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_5\
        );

    \I__1579\ : InMux
    port map (
            O => \N__18509\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\
        );

    \I__1578\ : InMux
    port map (
            O => \N__18506\,
            I => \N__18503\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__18503\,
            I => \N__18500\
        );

    \I__1576\ : Odrv4
    port map (
            O => \N__18500\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_6\
        );

    \I__1575\ : InMux
    port map (
            O => \N__18497\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\
        );

    \I__1574\ : InMux
    port map (
            O => \N__18494\,
            I => \N__18491\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__18491\,
            I => \N__18488\
        );

    \I__1572\ : Odrv4
    port map (
            O => \N__18488\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_7\
        );

    \I__1571\ : InMux
    port map (
            O => \N__18485\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\
        );

    \I__1570\ : InMux
    port map (
            O => \N__18482\,
            I => \N__18479\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__18479\,
            I => \N__18476\
        );

    \I__1568\ : Span4Mux_v
    port map (
            O => \N__18476\,
            I => \N__18473\
        );

    \I__1567\ : Odrv4
    port map (
            O => \N__18473\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_8\
        );

    \I__1566\ : InMux
    port map (
            O => \N__18470\,
            I => \bfn_1_14_0_\
        );

    \I__1565\ : InMux
    port map (
            O => \N__18467\,
            I => \N__18464\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__18464\,
            I => \N__18461\
        );

    \I__1563\ : Span4Mux_v
    port map (
            O => \N__18461\,
            I => \N__18458\
        );

    \I__1562\ : Odrv4
    port map (
            O => \N__18458\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_9\
        );

    \I__1561\ : InMux
    port map (
            O => \N__18455\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\
        );

    \I__1560\ : InMux
    port map (
            O => \N__18452\,
            I => \N__18449\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__18449\,
            I => \N__18446\
        );

    \I__1558\ : Odrv4
    port map (
            O => \N__18446\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_10\
        );

    \I__1557\ : InMux
    port map (
            O => \N__18443\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\
        );

    \I__1556\ : InMux
    port map (
            O => \N__18440\,
            I => \N__18437\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__18437\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_15\
        );

    \I__1554\ : InMux
    port map (
            O => \N__18434\,
            I => \N__18431\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__18431\,
            I => \N__18428\
        );

    \I__1552\ : Span4Mux_v
    port map (
            O => \N__18428\,
            I => \N__18425\
        );

    \I__1551\ : Odrv4
    port map (
            O => \N__18425\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_0\
        );

    \I__1550\ : CascadeMux
    port map (
            O => \N__18422\,
            I => \N__18419\
        );

    \I__1549\ : InMux
    port map (
            O => \N__18419\,
            I => \N__18416\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__18416\,
            I => \N__18413\
        );

    \I__1547\ : Span4Mux_v
    port map (
            O => \N__18413\,
            I => \N__18410\
        );

    \I__1546\ : Odrv4
    port map (
            O => \N__18410\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_15\
        );

    \I__1545\ : InMux
    port map (
            O => \N__18407\,
            I => \N__18404\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__18404\,
            I => \N__18401\
        );

    \I__1543\ : Span4Mux_v
    port map (
            O => \N__18401\,
            I => \N__18398\
        );

    \I__1542\ : Odrv4
    port map (
            O => \N__18398\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_1\
        );

    \I__1541\ : CascadeMux
    port map (
            O => \N__18395\,
            I => \N__18392\
        );

    \I__1540\ : InMux
    port map (
            O => \N__18392\,
            I => \N__18389\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__18389\,
            I => \N__18386\
        );

    \I__1538\ : Span4Mux_v
    port map (
            O => \N__18386\,
            I => \N__18383\
        );

    \I__1537\ : Odrv4
    port map (
            O => \N__18383\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_16\
        );

    \I__1536\ : InMux
    port map (
            O => \N__18380\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\
        );

    \I__1535\ : InMux
    port map (
            O => \N__18377\,
            I => \N__18374\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__18374\,
            I => \N__18371\
        );

    \I__1533\ : Span4Mux_h
    port map (
            O => \N__18371\,
            I => \N__18368\
        );

    \I__1532\ : Odrv4
    port map (
            O => \N__18368\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_2\
        );

    \I__1531\ : CascadeMux
    port map (
            O => \N__18365\,
            I => \N__18362\
        );

    \I__1530\ : InMux
    port map (
            O => \N__18362\,
            I => \N__18359\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__18359\,
            I => \N__18356\
        );

    \I__1528\ : Span4Mux_v
    port map (
            O => \N__18356\,
            I => \N__18353\
        );

    \I__1527\ : Odrv4
    port map (
            O => \N__18353\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_17\
        );

    \I__1526\ : InMux
    port map (
            O => \N__18350\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\
        );

    \I__1525\ : IoInMux
    port map (
            O => \N__18347\,
            I => \N__18344\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__18344\,
            I => \N__18341\
        );

    \I__1523\ : Span4Mux_s3_v
    port map (
            O => \N__18341\,
            I => \N__18338\
        );

    \I__1522\ : Span4Mux_h
    port map (
            O => \N__18338\,
            I => \N__18335\
        );

    \I__1521\ : Sp12to4
    port map (
            O => \N__18335\,
            I => \N__18332\
        );

    \I__1520\ : Span12Mux_v
    port map (
            O => \N__18332\,
            I => \N__18329\
        );

    \I__1519\ : Span12Mux_v
    port map (
            O => \N__18329\,
            I => \N__18326\
        );

    \I__1518\ : Odrv12
    port map (
            O => \N__18326\,
            I => delay_tr_input_ibuf_gb_io_gb_input
        );

    \I__1517\ : IoInMux
    port map (
            O => \N__18323\,
            I => \N__18320\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__18320\,
            I => \N__18317\
        );

    \I__1515\ : IoSpan4Mux
    port map (
            O => \N__18317\,
            I => \N__18314\
        );

    \I__1514\ : IoSpan4Mux
    port map (
            O => \N__18314\,
            I => \N__18311\
        );

    \I__1513\ : Odrv4
    port map (
            O => \N__18311\,
            I => delay_hc_input_ibuf_gb_io_gb_input
        );

    \IN_MUX_bfv_3_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_24_0_\
        );

    \IN_MUX_bfv_3_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_cry_7\,
            carryinitout => \bfn_3_25_0_\
        );

    \IN_MUX_bfv_3_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_cry_15\,
            carryinitout => \bfn_3_26_0_\
        );

    \IN_MUX_bfv_14_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_8_0_\
        );

    \IN_MUX_bfv_14_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_14_9_0_\
        );

    \IN_MUX_bfv_14_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_14_10_0_\
        );

    \IN_MUX_bfv_14_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_14_11_0_\
        );

    \IN_MUX_bfv_11_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_8_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_11_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_11_10_0_\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_11_11_0_\
        );

    \IN_MUX_bfv_17_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_10_0_\
        );

    \IN_MUX_bfv_17_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_17_11_0_\
        );

    \IN_MUX_bfv_17_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_17_12_0_\
        );

    \IN_MUX_bfv_17_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_17_13_0_\
        );

    \IN_MUX_bfv_8_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_5_0_\
        );

    \IN_MUX_bfv_8_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_8_6_0_\
        );

    \IN_MUX_bfv_8_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_8_7_0_\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_8_8_0_\
        );

    \IN_MUX_bfv_12_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_15_0_\
        );

    \IN_MUX_bfv_12_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s1\,
            carryinitout => \bfn_12_16_0_\
        );

    \IN_MUX_bfv_12_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s1\,
            carryinitout => \bfn_12_17_0_\
        );

    \IN_MUX_bfv_12_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s1\,
            carryinitout => \bfn_12_18_0_\
        );

    \IN_MUX_bfv_14_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_13_0_\
        );

    \IN_MUX_bfv_14_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s0\,
            carryinitout => \bfn_14_14_0_\
        );

    \IN_MUX_bfv_14_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s0\,
            carryinitout => \bfn_14_15_0_\
        );

    \IN_MUX_bfv_14_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s0\,
            carryinitout => \bfn_14_16_0_\
        );

    \IN_MUX_bfv_16_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_14_0_\
        );

    \IN_MUX_bfv_16_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_7\,
            carryinitout => \bfn_16_15_0_\
        );

    \IN_MUX_bfv_16_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_15\,
            carryinitout => \bfn_16_16_0_\
        );

    \IN_MUX_bfv_16_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_23\,
            carryinitout => \bfn_16_17_0_\
        );

    \IN_MUX_bfv_2_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_13_0_\
        );

    \IN_MUX_bfv_2_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            carryinitout => \bfn_2_14_0_\
        );

    \IN_MUX_bfv_2_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            carryinitout => \bfn_2_15_0_\
        );

    \IN_MUX_bfv_2_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            carryinitout => \bfn_2_16_0_\
        );

    \IN_MUX_bfv_3_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_17_0_\
        );

    \IN_MUX_bfv_3_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            carryinitout => \bfn_3_18_0_\
        );

    \IN_MUX_bfv_3_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            carryinitout => \bfn_3_19_0_\
        );

    \IN_MUX_bfv_3_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            carryinitout => \bfn_3_20_0_\
        );

    \IN_MUX_bfv_4_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_23_0_\
        );

    \IN_MUX_bfv_4_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_add_1_cry_7\,
            carryinitout => \bfn_4_24_0_\
        );

    \IN_MUX_bfv_4_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_add_1_cry_15\,
            carryinitout => \bfn_4_25_0_\
        );

    \IN_MUX_bfv_7_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_23_0_\
        );

    \IN_MUX_bfv_7_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un19_threshold_cry_7\,
            carryinitout => \bfn_7_24_0_\
        );

    \IN_MUX_bfv_5_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_25_0_\
        );

    \IN_MUX_bfv_5_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_1_cry_7\,
            carryinitout => \bfn_5_26_0_\
        );

    \IN_MUX_bfv_5_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_1_cry_15\,
            carryinitout => \bfn_5_27_0_\
        );

    \IN_MUX_bfv_9_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_24_0_\
        );

    \IN_MUX_bfv_9_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un14_counter_cry_7\,
            carryinitout => \bfn_9_25_0_\
        );

    \IN_MUX_bfv_10_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_24_0_\
        );

    \IN_MUX_bfv_10_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.counter_cry_7\,
            carryinitout => \bfn_10_25_0_\
        );

    \IN_MUX_bfv_15_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_7_0_\
        );

    \IN_MUX_bfv_15_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un4_running_cry_8\,
            carryinitout => \bfn_15_8_0_\
        );

    \IN_MUX_bfv_15_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un4_running_cry_16\,
            carryinitout => \bfn_15_9_0_\
        );

    \IN_MUX_bfv_10_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_7_0_\
        );

    \IN_MUX_bfv_10_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un4_running_cry_8\,
            carryinitout => \bfn_10_8_0_\
        );

    \IN_MUX_bfv_10_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un4_running_cry_16\,
            carryinitout => \bfn_10_9_0_\
        );

    \IN_MUX_bfv_16_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_11_0_\
        );

    \IN_MUX_bfv_16_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un4_running_cry_8\,
            carryinitout => \bfn_16_12_0_\
        );

    \IN_MUX_bfv_16_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un4_running_cry_16\,
            carryinitout => \bfn_16_13_0_\
        );

    \IN_MUX_bfv_8_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_9_0_\
        );

    \IN_MUX_bfv_8_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un4_running_cry_8\,
            carryinitout => \bfn_8_10_0_\
        );

    \IN_MUX_bfv_8_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un4_running_cry_16\,
            carryinitout => \bfn_8_11_0_\
        );

    \IN_MUX_bfv_15_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_10_0_\
        );

    \IN_MUX_bfv_15_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_15_11_0_\
        );

    \IN_MUX_bfv_15_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_15_12_0_\
        );

    \IN_MUX_bfv_15_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_15_13_0_\
        );

    \IN_MUX_bfv_13_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_10_0_\
        );

    \IN_MUX_bfv_13_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            carryinitout => \bfn_13_11_0_\
        );

    \IN_MUX_bfv_13_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            carryinitout => \bfn_13_12_0_\
        );

    \IN_MUX_bfv_13_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            carryinitout => \bfn_13_13_0_\
        );

    \IN_MUX_bfv_10_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_12_0_\
        );

    \IN_MUX_bfv_10_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_10_13_0_\
        );

    \IN_MUX_bfv_10_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_10_14_0_\
        );

    \IN_MUX_bfv_10_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_10_15_0_\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_15_0_\
        );

    \IN_MUX_bfv_9_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            carryinitout => \bfn_9_16_0_\
        );

    \IN_MUX_bfv_9_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            carryinitout => \bfn_9_17_0_\
        );

    \IN_MUX_bfv_9_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            carryinitout => \bfn_9_18_0_\
        );

    \IN_MUX_bfv_9_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_19_0_\
        );

    \IN_MUX_bfv_9_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_7\,
            carryinitout => \bfn_9_20_0_\
        );

    \IN_MUX_bfv_15_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_18_0_\
        );

    \IN_MUX_bfv_15_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_15_19_0_\
        );

    \IN_MUX_bfv_15_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_15_20_0_\
        );

    \IN_MUX_bfv_15_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_15_21_0_\
        );

    \IN_MUX_bfv_18_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_14_0_\
        );

    \IN_MUX_bfv_18_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_8\,
            carryinitout => \bfn_18_15_0_\
        );

    \IN_MUX_bfv_18_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_16\,
            carryinitout => \bfn_18_16_0_\
        );

    \IN_MUX_bfv_18_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_24\,
            carryinitout => \bfn_18_17_0_\
        );

    \IN_MUX_bfv_17_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_18_0_\
        );

    \IN_MUX_bfv_17_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_7\,
            carryinitout => \bfn_17_19_0_\
        );

    \IN_MUX_bfv_17_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_15\,
            carryinitout => \bfn_17_20_0_\
        );

    \IN_MUX_bfv_17_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_23\,
            carryinitout => \bfn_17_21_0_\
        );

    \IN_MUX_bfv_1_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_13_0_\
        );

    \IN_MUX_bfv_1_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\,
            carryinitout => \bfn_1_14_0_\
        );

    \IN_MUX_bfv_8_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_19_0_\
        );

    \IN_MUX_bfv_8_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            carryinitout => \bfn_8_20_0_\
        );

    \delay_tr_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__18347\,
            GLOBALBUFFEROUTPUT => delay_tr_input_c_g
        );

    \delay_hc_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__18323\,
            GLOBALBUFFEROUTPUT => delay_hc_input_c_g
        );

    \current_shift_inst.timer_s1.running_RNII51H_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__33686\,
            GLOBALBUFFEROUTPUT => \current_shift_inst.timer_s1.N_162_i_g\
        );

    \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__34180\,
            GLOBALBUFFEROUTPUT => \phase_controller_inst2.stoper_tr.un1_start_g\
        );

    \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__32198\,
            GLOBALBUFFEROUTPUT => \phase_controller_inst2.stoper_hc.un1_start_g\
        );

    \osc\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b10"
        )
    port map (
            CLKHFPU => \N__38001\,
            CLKHFEN => \N__38003\,
            CLKHF => clk_12mhz
        );

    \rgb_drv\ : SB_RGBA_DRV
    generic map (
            RGB2_CURRENT => "0b111111",
            CURRENT_MODE => "0b0",
            RGB0_CURRENT => "0b111111",
            RGB1_CURRENT => "0b111111"
        )
    port map (
            RGBLEDEN => \N__38002\,
            RGB2PWM => \N__18752\,
            RGB1 => rgb_g_wire,
            CURREN => \N__37975\,
            RGB2 => rgb_b_wire,
            RGB1PWM => \N__18746\,
            RGB0PWM => \N__46961\,
            RGB0 => rgb_r_wire
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18440\,
            in2 => \_gnd_net_\,
            in3 => \N__18652\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18434\,
            in2 => \N__18422\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_16\,
            ltout => OPEN,
            carryin => \bfn_1_13_0_\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18407\,
            in2 => \N__18395\,
            in3 => \N__18380\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18377\,
            in2 => \N__18365\,
            in3 => \N__18350\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18566\,
            in2 => \N__18554\,
            in3 => \N__18536\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18621\,
            in2 => \N__18533\,
            in3 => \N__18521\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18518\,
            in2 => \N__18653\,
            in3 => \N__18509\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18506\,
            in2 => \N__18658\,
            in3 => \N__18497\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18494\,
            in2 => \N__18654\,
            in3 => \N__18485\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18482\,
            in2 => \N__18659\,
            in3 => \N__18470\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_24\,
            ltout => OPEN,
            carryin => \bfn_1_14_0_\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18467\,
            in2 => \N__18655\,
            in3 => \N__18455\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18452\,
            in2 => \N__18660\,
            in3 => \N__18443\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18710\,
            in2 => \N__18656\,
            in3 => \N__18701\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18698\,
            in2 => \N__18661\,
            in3 => \N__18689\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18686\,
            in2 => \N__18657\,
            in3 => \N__18677\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18674\,
            in2 => \N__18662\,
            in3 => \N__18572\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18569\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_29_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001100"
        )
    port map (
            in0 => \N__23064\,
            in1 => \N__23255\,
            in2 => \N__22634\,
            in3 => \N__19328\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47673\,
            ce => 'H',
            sr => \N__46919\
        );

    \current_shift_inst.PI_CTRL.integrator_18_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001100"
        )
    port map (
            in0 => \N__23063\,
            in1 => \N__23254\,
            in2 => \N__22633\,
            in3 => \N__19247\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47673\,
            ce => 'H',
            sr => \N__46919\
        );

    \current_shift_inst.PI_CTRL.integrator_12_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101010"
        )
    port map (
            in0 => \N__23181\,
            in1 => \N__23077\,
            in2 => \N__19064\,
            in3 => \N__22598\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47662\,
            ce => 'H',
            sr => \N__46923\
        );

    \current_shift_inst.PI_CTRL.integrator_27_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111001000100"
        )
    port map (
            in0 => \N__22597\,
            in1 => \N__23182\,
            in2 => \N__23084\,
            in3 => \N__19367\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47662\,
            ce => 'H',
            sr => \N__46923\
        );

    \current_shift_inst.PI_CTRL.integrator_2_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__18935\,
            in1 => \N__23076\,
            in2 => \_gnd_net_\,
            in3 => \N__22609\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47652\,
            ce => 'H',
            sr => \N__46927\
        );

    \current_shift_inst.PI_CTRL.prop_term_0_LC_1_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24997\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47639\,
            ce => 'H',
            sr => \N__46931\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_0_LC_1_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18740\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47617\,
            ce => 'H',
            sr => \N__46936\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_1_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__19511\,
            in1 => \N__43843\,
            in2 => \_gnd_net_\,
            in3 => \N__19799\,
            lcout => \current_shift_inst.PI_CTRL.N_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_1_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101010101"
        )
    port map (
            in0 => \N__43844\,
            in1 => \N__19798\,
            in2 => \N__20686\,
            in3 => \N__19510\,
            lcout => \current_shift_inst.PI_CTRL.N_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_7_LC_1_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001100100010"
        )
    port map (
            in0 => \N__19818\,
            in1 => \N__43845\,
            in2 => \N__19488\,
            in3 => \N__20462\,
            lcout => pwm_duty_input_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47596\,
            ce => 'H',
            sr => \N__46937\
        );

    \current_shift_inst.PI_CTRL.control_out_2_LC_1_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__18731\,
            in1 => \N__19937\,
            in2 => \N__19745\,
            in3 => \N__19448\,
            lcout => pwm_duty_input_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47596\,
            ce => 'H',
            sr => \N__46937\
        );

    \current_shift_inst.PI_CTRL.control_out_1_LC_1_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__19445\,
            in1 => \N__19271\,
            in2 => \N__19737\,
            in3 => \N__18730\,
            lcout => pwm_duty_input_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47596\,
            ce => 'H',
            sr => \N__46937\
        );

    \current_shift_inst.PI_CTRL.control_out_0_LC_1_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__18729\,
            in1 => \N__18719\,
            in2 => \N__19744\,
            in3 => \N__19447\,
            lcout => pwm_duty_input_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47596\,
            ce => 'H',
            sr => \N__46937\
        );

    \current_shift_inst.PI_CTRL.control_out_3_LC_1_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110011011101"
        )
    port map (
            in0 => \N__19446\,
            in1 => \N__20645\,
            in2 => \N__19823\,
            in3 => \N__19757\,
            lcout => pwm_duty_input_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47596\,
            ce => 'H',
            sr => \N__46937\
        );

    \current_shift_inst.PI_CTRL.control_out_9_LC_1_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111100001010"
        )
    port map (
            in0 => \N__19807\,
            in1 => \N__19490\,
            in2 => \N__43855\,
            in3 => \N__20393\,
            lcout => pwm_duty_input_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47589\,
            ce => 'H',
            sr => \N__46939\
        );

    \current_shift_inst.PI_CTRL.control_out_5_LC_1_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011111100"
        )
    port map (
            in0 => \N__19489\,
            in1 => \N__19808\,
            in2 => \N__20498\,
            in3 => \N__43846\,
            lcout => pwm_duty_input_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47589\,
            ce => 'H',
            sr => \N__46939\
        );

    \current_shift_inst.PI_CTRL.control_out_4_LC_1_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001100110011"
        )
    port map (
            in0 => \N__20687\,
            in1 => \N__18761\,
            in2 => \N__20363\,
            in3 => \N__19495\,
            lcout => pwm_duty_input_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47589\,
            ce => 'H',
            sr => \N__46939\
        );

    \current_shift_inst.PI_CTRL.control_out_6_LC_1_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101110"
        )
    port map (
            in0 => \N__20429\,
            in1 => \N__19809\,
            in2 => \N__19496\,
            in3 => \N__43847\,
            lcout => pwm_duty_input_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47589\,
            ce => 'H',
            sr => \N__46939\
        );

    \current_shift_inst.PI_CTRL.control_out_8_LC_1_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011111010"
        )
    port map (
            in0 => \N__20525\,
            in1 => \N__19494\,
            in2 => \N__19822\,
            in3 => \N__43851\,
            lcout => pwm_duty_input_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47583\,
            ce => 'H',
            sr => \N__46940\
        );

    \phase_controller_inst1.N_42_i_i_LC_1_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__30826\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46959\,
            lcout => \N_42_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.un7_start_stop_0_a2_LC_1_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__46960\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30827\,
            lcout => un7_start_stop_0_a2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_4_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101100"
        )
    port map (
            in0 => \N__23082\,
            in1 => \N__23223\,
            in2 => \N__18878\,
            in3 => \N__22602\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47694\,
            ce => 'H',
            sr => \N__46903\
        );

    \current_shift_inst.PI_CTRL.integrator_5_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100010011000101"
        )
    port map (
            in0 => \N__23222\,
            in1 => \N__18848\,
            in2 => \N__22631\,
            in3 => \N__23083\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47694\,
            ce => 'H',
            sr => \N__46903\
        );

    \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20824\,
            in2 => \N__19900\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_13_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20880\,
            in2 => \N__18953\,
            in3 => \N__18923\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22862\,
            in2 => \N__18920\,
            in3 => \N__18899\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22766\,
            in2 => \N__18896\,
            in3 => \N__18869\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22820\,
            in2 => \N__18866\,
            in3 => \N__18842\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20787\,
            in2 => \N__18839\,
            in3 => \N__18821\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22912\,
            in2 => \N__18818\,
            in3 => \N__18803\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21244\,
            in2 => \N__18800\,
            in3 => \N__18782\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23287\,
            in2 => \N__18779\,
            in3 => \N__18764\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_2_14_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21119\,
            in2 => \N__19124\,
            in3 => \N__19106\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21356\,
            in2 => \N__19103\,
            in3 => \N__19085\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21296\,
            in2 => \N__19082\,
            in3 => \N__19049\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21157\,
            in2 => \N__19046\,
            in3 => \N__19028\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21389\,
            in2 => \N__19025\,
            in3 => \N__19007\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21187\,
            in2 => \N__19004\,
            in3 => \N__18986\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21090\,
            in2 => \N__18983\,
            in3 => \N__18974\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20974\,
            in2 => \N__18971\,
            in3 => \N__18956\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_2_15_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21032\,
            in2 => \N__19259\,
            in3 => \N__19241\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21061\,
            in2 => \N__19238\,
            in3 => \N__19226\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21570\,
            in2 => \N__19223\,
            in3 => \N__19211\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20947\,
            in2 => \N__19208\,
            in3 => \N__19193\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21005\,
            in2 => \N__19190\,
            in3 => \N__19175\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22695\,
            in2 => \N__19172\,
            in3 => \N__19157\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21597\,
            in2 => \N__19154\,
            in3 => \N__19145\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21462\,
            in2 => \N__19142\,
            in3 => \N__19127\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\,
            ltout => OPEN,
            carryin => \bfn_2_16_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21517\,
            in2 => \N__19400\,
            in3 => \N__19385\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_2_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21423\,
            in2 => \N__19382\,
            in3 => \N__19361\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21493\,
            in2 => \N__19358\,
            in3 => \N__19343\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22727\,
            in2 => \N__19340\,
            in3 => \N__19322\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21334\,
            in2 => \N__19319\,
            in3 => \N__19307\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19304\,
            in1 => \N__23159\,
            in2 => \N__19295\,
            in3 => \N__19280\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_31_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001100"
        )
    port map (
            in0 => \N__23081\,
            in1 => \N__23189\,
            in2 => \N__22632\,
            in3 => \N__19277\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47641\,
            ce => 'H',
            sr => \N__46924\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21637\,
            in2 => \_gnd_net_\,
            in3 => \N__20845\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47628\,
            ce => 'H',
            sr => \N__46928\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20379\,
            in2 => \_gnd_net_\,
            in3 => \N__20484\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_2_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20219\,
            in1 => \N__20581\,
            in2 => \N__20549\,
            in3 => \N__20233\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_2_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19996\,
            in2 => \_gnd_net_\,
            in3 => \N__20032\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_2_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20170\,
            in1 => \N__20017\,
            in2 => \N__19433\,
            in3 => \N__19430\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_2_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20033\,
            in1 => \N__20156\,
            in2 => \N__20116\,
            in3 => \N__20137\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_2_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20155\,
            in1 => \N__20218\,
            in2 => \N__20234\,
            in3 => \N__20065\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_2_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20021\,
            in1 => \N__19424\,
            in2 => \N__20003\,
            in3 => \N__19550\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_2_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20704\,
            in2 => \_gnd_net_\,
            in3 => \N__20183\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_2_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20171\,
            in1 => \N__20251\,
            in2 => \N__19418\,
            in3 => \N__20066\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_2_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19415\,
            in1 => \N__19517\,
            in2 => \N__19409\,
            in3 => \N__19406\,
            lcout => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_2_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20083\,
            in2 => \_gnd_net_\,
            in3 => \N__20095\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_2_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__20524\,
            in1 => \N__19544\,
            in2 => \N__20461\,
            in3 => \N__20418\,
            lcout => \current_shift_inst.PI_CTRL.N_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_2_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20182\,
            in1 => \N__20084\,
            in2 => \N__20705\,
            in3 => \N__20096\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_2_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__20138\,
            in1 => \_gnd_net_\,
            in2 => \N__20120\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_2_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20194\,
            in1 => \N__20206\,
            in2 => \N__19538\,
            in3 => \N__20252\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_2_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19535\,
            in1 => \N__20531\,
            in2 => \N__19529\,
            in3 => \N__19526\,
            lcout => \current_shift_inst.PI_CTRL.N_159\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_2_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20207\,
            in1 => \N__20563\,
            in2 => \N__20606\,
            in3 => \N__20195\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__20679\,
            in1 => \N__43804\,
            in2 => \_gnd_net_\,
            in3 => \N__19509\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__19464\,
            in1 => \N__20612\,
            in2 => \N__20356\,
            in3 => \N__43821\,
            lcout => \current_shift_inst.PI_CTRL.N_96\,
            ltout => \current_shift_inst.PI_CTRL.N_96_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101010000"
        )
    port map (
            in0 => \N__20641\,
            in1 => \N__19803\,
            in2 => \N__19760\,
            in3 => \N__19756\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un1_duty_inputlto2_LC_2_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__19714\,
            in1 => \N__19699\,
            in2 => \_gnd_net_\,
            in3 => \N__19681\,
            lcout => \pwm_generator_inst.un1_duty_inputlt3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19636\,
            in2 => \_gnd_net_\,
            in3 => \N__20277\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__19617\,
            in1 => \N__19595\,
            in2 => \N__19667\,
            in3 => \N__19654\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_LC_2_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111011"
        )
    port map (
            in0 => \N__19664\,
            in1 => \N__20328\,
            in2 => \N__19658\,
            in3 => \N__20304\,
            lcout => \pwm_generator_inst.N_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19653\,
            in1 => \N__19635\,
            in2 => \N__19619\,
            in3 => \N__19594\,
            lcout => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_14_LC_3_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101010"
        )
    port map (
            in0 => \N__23228\,
            in1 => \N__23047\,
            in2 => \N__19577\,
            in3 => \N__22629\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47663\,
            ce => 'H',
            sr => \N__46907\
        );

    \current_shift_inst.PI_CTRL.integrator_11_LC_3_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010011100100"
        )
    port map (
            in0 => \N__22624\,
            in1 => \N__23230\,
            in2 => \N__19568\,
            in3 => \N__23051\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47663\,
            ce => 'H',
            sr => \N__46907\
        );

    \current_shift_inst.PI_CTRL.integrator_16_LC_3_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010011100100"
        )
    port map (
            in0 => \N__22626\,
            in1 => \N__23232\,
            in2 => \N__19559\,
            in3 => \N__23053\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47663\,
            ce => 'H',
            sr => \N__46907\
        );

    \current_shift_inst.PI_CTRL.integrator_15_LC_3_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101010"
        )
    port map (
            in0 => \N__23229\,
            in1 => \N__23048\,
            in2 => \N__19916\,
            in3 => \N__22630\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47663\,
            ce => 'H',
            sr => \N__46907\
        );

    \current_shift_inst.PI_CTRL.integrator_1_LC_3_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000101000"
        )
    port map (
            in0 => \N__22627\,
            in1 => \N__20834\,
            in2 => \N__19907\,
            in3 => \N__23054\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47663\,
            ce => 'H',
            sr => \N__46907\
        );

    \current_shift_inst.PI_CTRL.integrator_10_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101010"
        )
    port map (
            in0 => \N__23227\,
            in1 => \N__23046\,
            in2 => \N__19877\,
            in3 => \N__22628\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47663\,
            ce => 'H',
            sr => \N__46907\
        );

    \current_shift_inst.PI_CTRL.integrator_13_LC_3_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010011100100"
        )
    port map (
            in0 => \N__22625\,
            in1 => \N__23231\,
            in2 => \N__19868\,
            in3 => \N__23052\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47663\,
            ce => 'H',
            sr => \N__46907\
        );

    \current_shift_inst.PI_CTRL.integrator_24_LC_3_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110011011000"
        )
    port map (
            in0 => \N__22615\,
            in1 => \N__19859\,
            in2 => \N__23259\,
            in3 => \N__23039\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47653\,
            ce => 'H',
            sr => \N__46911\
        );

    \current_shift_inst.PI_CTRL.integrator_19_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101100"
        )
    port map (
            in0 => \N__23035\,
            in1 => \N__23234\,
            in2 => \N__19853\,
            in3 => \N__22616\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47653\,
            ce => 'H',
            sr => \N__46911\
        );

    \current_shift_inst.PI_CTRL.integrator_22_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110011011000"
        )
    port map (
            in0 => \N__22614\,
            in1 => \N__19844\,
            in2 => \N__23258\,
            in3 => \N__23038\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47653\,
            ce => 'H',
            sr => \N__46911\
        );

    \current_shift_inst.PI_CTRL.integrator_23_LC_3_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101100"
        )
    port map (
            in0 => \N__23036\,
            in1 => \N__23235\,
            in2 => \N__19838\,
            in3 => \N__22617\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47653\,
            ce => 'H',
            sr => \N__46911\
        );

    \current_shift_inst.PI_CTRL.integrator_20_LC_3_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110011011000"
        )
    port map (
            in0 => \N__22613\,
            in1 => \N__19829\,
            in2 => \N__23257\,
            in3 => \N__23037\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47653\,
            ce => 'H',
            sr => \N__46911\
        );

    \current_shift_inst.PI_CTRL.integrator_30_LC_3_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001010"
        )
    port map (
            in0 => \N__23185\,
            in1 => \N__23045\,
            in2 => \N__22608\,
            in3 => \N__19982\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47642\,
            ce => 'H',
            sr => \N__46916\
        );

    \current_shift_inst.PI_CTRL.integrator_17_LC_3_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001111100000"
        )
    port map (
            in0 => \N__23040\,
            in1 => \N__22541\,
            in2 => \N__19976\,
            in3 => \N__23188\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47642\,
            ce => 'H',
            sr => \N__46916\
        );

    \current_shift_inst.PI_CTRL.integrator_21_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001010"
        )
    port map (
            in0 => \N__23183\,
            in1 => \N__23043\,
            in2 => \N__22606\,
            in3 => \N__19967\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47642\,
            ce => 'H',
            sr => \N__46916\
        );

    \current_shift_inst.PI_CTRL.integrator_25_LC_3_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001010"
        )
    port map (
            in0 => \N__23184\,
            in1 => \N__23044\,
            in2 => \N__22607\,
            in3 => \N__19961\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47642\,
            ce => 'H',
            sr => \N__46916\
        );

    \current_shift_inst.PI_CTRL.integrator_26_LC_3_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101100"
        )
    port map (
            in0 => \N__23041\,
            in1 => \N__23186\,
            in2 => \N__19955\,
            in3 => \N__22551\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47642\,
            ce => 'H',
            sr => \N__46916\
        );

    \current_shift_inst.PI_CTRL.integrator_28_LC_3_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101100"
        )
    port map (
            in0 => \N__23042\,
            in1 => \N__23187\,
            in2 => \N__19946\,
            in3 => \N__22552\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47642\,
            ce => 'H',
            sr => \N__46916\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21638\,
            in2 => \N__20846\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_17_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_2_LC_3_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22445\,
            in2 => \N__20885\,
            in3 => \N__19922\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            clk => \N__47629\,
            ce => 'H',
            sr => \N__46920\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_3_LC_3_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22454\,
            in2 => \N__22874\,
            in3 => \N__19919\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            clk => \N__47629\,
            ce => 'H',
            sr => \N__46920\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_4_LC_3_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21617\,
            in2 => \N__22792\,
            in3 => \N__20051\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            clk => \N__47629\,
            ce => 'H',
            sr => \N__46920\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_5_LC_3_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22831\,
            in2 => \N__21677\,
            in3 => \N__20048\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            clk => \N__47629\,
            ce => 'H',
            sr => \N__46920\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_6_LC_3_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21263\,
            in2 => \N__20795\,
            in3 => \N__20045\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            clk => \N__47629\,
            ce => 'H',
            sr => \N__46920\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_7_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21668\,
            in2 => \N__22916\,
            in3 => \N__20042\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            clk => \N__47629\,
            ce => 'H',
            sr => \N__46920\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_8_LC_3_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21257\,
            in2 => \N__21251\,
            in3 => \N__20039\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            clk => \N__47629\,
            ce => 'H',
            sr => \N__46920\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_9_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21650\,
            in2 => \N__23294\,
            in3 => \N__20036\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_3_18_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            clk => \N__47618\,
            ce => 'H',
            sr => \N__46925\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_10_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21611\,
            in2 => \N__21137\,
            in3 => \N__20024\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            clk => \N__47618\,
            ce => 'H',
            sr => \N__46925\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_11_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21656\,
            in2 => \N__21371\,
            in3 => \N__20006\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            clk => \N__47618\,
            ce => 'H',
            sr => \N__46925\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_12_LC_3_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21644\,
            in2 => \N__21314\,
            in3 => \N__19985\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            clk => \N__47618\,
            ce => 'H',
            sr => \N__46925\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_13_LC_3_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21662\,
            in2 => \N__21167\,
            in3 => \N__20144\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            clk => \N__47618\,
            ce => 'H',
            sr => \N__46925\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_14_LC_3_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22008\,
            in2 => \N__21404\,
            in3 => \N__20141\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            clk => \N__47618\,
            ce => 'H',
            sr => \N__46925\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_15_LC_3_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21194\,
            in2 => \N__22042\,
            in3 => \N__20123\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            clk => \N__47618\,
            ce => 'H',
            sr => \N__46925\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_16_LC_3_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22012\,
            in2 => \N__21101\,
            in3 => \N__20099\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            clk => \N__47618\,
            ce => 'H',
            sr => \N__46925\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_17_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22013\,
            in2 => \N__20981\,
            in3 => \N__20087\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_3_19_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            clk => \N__47606\,
            ce => 'H',
            sr => \N__46929\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_18_LC_3_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21041\,
            in2 => \N__22043\,
            in3 => \N__20075\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            clk => \N__47606\,
            ce => 'H',
            sr => \N__46929\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_19_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22017\,
            in2 => \N__21068\,
            in3 => \N__20072\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            clk => \N__47606\,
            ce => 'H',
            sr => \N__46929\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_20_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21575\,
            in2 => \N__22044\,
            in3 => \N__20069\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            clk => \N__47606\,
            ce => 'H',
            sr => \N__46929\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_21_LC_3_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22021\,
            in2 => \N__20954\,
            in3 => \N__20054\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            clk => \N__47606\,
            ce => 'H',
            sr => \N__46929\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_22_LC_3_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21011\,
            in2 => \N__22045\,
            in3 => \N__20237\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            clk => \N__47606\,
            ce => 'H',
            sr => \N__46929\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_23_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22025\,
            in2 => \N__22703\,
            in3 => \N__20222\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            clk => \N__47606\,
            ce => 'H',
            sr => \N__46929\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_24_LC_3_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21605\,
            in2 => \N__22046\,
            in3 => \N__20210\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            clk => \N__47606\,
            ce => 'H',
            sr => \N__46929\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_25_LC_3_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22029\,
            in2 => \N__21473\,
            in3 => \N__20198\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_3_20_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            clk => \N__47597\,
            ce => 'H',
            sr => \N__46932\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_26_LC_3_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21521\,
            in2 => \N__22047\,
            in3 => \N__20186\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            clk => \N__47597\,
            ce => 'H',
            sr => \N__46932\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_27_LC_3_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22033\,
            in2 => \N__21440\,
            in3 => \N__20174\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            clk => \N__47597\,
            ce => 'H',
            sr => \N__46932\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_28_LC_3_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21497\,
            in2 => \N__22048\,
            in3 => \N__20159\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            clk => \N__47597\,
            ce => 'H',
            sr => \N__46932\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_29_LC_3_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22037\,
            in2 => \N__22742\,
            in3 => \N__20147\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            clk => \N__47597\,
            ce => 'H',
            sr => \N__46932\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_30_LC_3_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21338\,
            in2 => \N__22049\,
            in3 => \N__20693\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\,
            clk => \N__47597\,
            ce => 'H',
            sr => \N__46932\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_31_LC_3_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23256\,
            in1 => \N__22041\,
            in2 => \_gnd_net_\,
            in3 => \N__20690\,
            lcout => \current_shift_inst.PI_CTRL.un8_enablelto31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47597\,
            ce => 'H',
            sr => \N__46932\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_3_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20669\,
            in2 => \_gnd_net_\,
            in3 => \N__20634\,
            lcout => \current_shift_inst.PI_CTRL.N_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_3_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20599\,
            in1 => \N__20582\,
            in2 => \N__20567\,
            in3 => \N__20548\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_3_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20520\,
            in2 => \_gnd_net_\,
            in3 => \N__20491\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_3_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20457\,
            in1 => \N__20425\,
            in2 => \N__20396\,
            in3 => \N__20386\,
            lcout => \current_shift_inst.PI_CTRL.N_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_LC_3_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__20339\,
            in1 => \N__20308\,
            in2 => \N__20285\,
            in3 => \N__20258\,
            lcout => \pwm_generator_inst.N_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_3_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__23565\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22291\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_0_c_LC_3_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23530\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_24_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_3_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20756\,
            in2 => \_gnd_net_\,
            in3 => \N__20747\,
            lcout => \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_0\,
            carryout => \pwm_generator_inst.un3_threshold_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_3_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20744\,
            in2 => \_gnd_net_\,
            in3 => \N__20735\,
            lcout => \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_1\,
            carryout => \pwm_generator_inst.un3_threshold_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_3_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20732\,
            in2 => \_gnd_net_\,
            in3 => \N__20723\,
            lcout => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_2\,
            carryout => \pwm_generator_inst.un3_threshold_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_3_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21932\,
            in2 => \_gnd_net_\,
            in3 => \N__20720\,
            lcout => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_3\,
            carryout => \pwm_generator_inst.un3_threshold_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_3_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37818\,
            in2 => \N__21893\,
            in3 => \N__20717\,
            lcout => \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_4\,
            carryout => \pwm_generator_inst.un3_threshold_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_3_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21851\,
            in2 => \N__37917\,
            in3 => \N__20714\,
            lcout => \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_5\,
            carryout => \pwm_generator_inst.un3_threshold_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_3_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37822\,
            in2 => \N__21812\,
            in3 => \N__20711\,
            lcout => \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_6\,
            carryout => \pwm_generator_inst.un3_threshold_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_3_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21770\,
            in2 => \_gnd_net_\,
            in3 => \N__20708\,
            lcout => \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11\,
            ltout => OPEN,
            carryin => \bfn_3_25_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_9_c_LC_3_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21731\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_8\,
            carryout => \pwm_generator_inst.un3_threshold_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_10_c_LC_3_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21689\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_9\,
            carryout => \pwm_generator_inst.un3_threshold_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_11_c_LC_3_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22247\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_10\,
            carryout => \pwm_generator_inst.un3_threshold_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_12_c_LC_3_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22202\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_11\,
            carryout => \pwm_generator_inst.un3_threshold_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_13_c_LC_3_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22160\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_12\,
            carryout => \pwm_generator_inst.un3_threshold_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_14_c_LC_3_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22136\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_13\,
            carryout => \pwm_generator_inst.un3_threshold_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_15_c_LC_3_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22112\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_14\,
            carryout => \pwm_generator_inst.un3_threshold_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_16_c_LC_3_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22088\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_26_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_17_c_LC_3_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22064\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_16\,
            carryout => \pwm_generator_inst.un3_threshold_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_18_c_LC_3_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22337\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_17\,
            carryout => \pwm_generator_inst.un3_threshold_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_c_LC_3_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22325\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_18\,
            carryout => \pwm_generator_inst.un3_threshold_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_3_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20924\,
            lcout => \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_3_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__20921\,
            in1 => \N__23073\,
            in2 => \_gnd_net_\,
            in3 => \N__22612\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47684\,
            ce => 'H',
            sr => \N__46888\
        );

    \current_shift_inst.PI_CTRL.integrator_8_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011000010110001"
        )
    port map (
            in0 => \N__22610\,
            in1 => \N__23261\,
            in2 => \N__20909\,
            in3 => \N__23075\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47664\,
            ce => 'H',
            sr => \N__46899\
        );

    \current_shift_inst.PI_CTRL.integrator_6_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100000011110001"
        )
    port map (
            in0 => \N__23074\,
            in1 => \N__22611\,
            in2 => \N__20897\,
            in3 => \N__23260\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47664\,
            ce => 'H',
            sr => \N__46899\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010111"
        )
    port map (
            in0 => \N__22873\,
            in1 => \N__20884\,
            in2 => \N__20838\,
            in3 => \N__22791\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_77_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__23283\,
            in1 => \N__20791\,
            in2 => \N__20798\,
            in3 => \N__21218\,
            lcout => \current_shift_inst.PI_CTRL.N_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21239\,
            in1 => \N__20780\,
            in2 => \N__22908\,
            in3 => \N__23282\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21363\,
            in1 => \N__21091\,
            in2 => \N__21313\,
            in3 => \N__21396\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__21240\,
            in1 => \N__22830\,
            in2 => \_gnd_net_\,
            in3 => \N__22904\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21060\,
            in1 => \N__21036\,
            in2 => \N__21010\,
            in3 => \N__20973\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21186\,
            in1 => \N__21156\,
            in2 => \N__21130\,
            in3 => \N__22732\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21212\,
            in1 => \N__21203\,
            in2 => \N__21197\,
            in3 => \N__21533\,
            lcout => \current_shift_inst.PI_CTRL.N_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21185\,
            in1 => \N__21155\,
            in2 => \N__21129\,
            in3 => \N__21089\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21059\,
            in1 => \N__21037\,
            in2 => \N__21009\,
            in3 => \N__20972\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23233\,
            in1 => \N__20946\,
            in2 => \N__21574\,
            in3 => \N__21598\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21515\,
            in2 => \_gnd_net_\,
            in3 => \N__20945\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__21596\,
            in1 => \N__21566\,
            in2 => \N__21545\,
            in3 => \N__21527\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__21542\,
            in1 => \N__23245\,
            in2 => \N__21536\,
            in3 => \N__22694\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21491\,
            in1 => \N__21458\,
            in2 => \N__21439\,
            in3 => \N__21332\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21516\,
            in1 => \N__21492\,
            in2 => \N__21466\,
            in3 => \N__21435\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21397\,
            in2 => \_gnd_net_\,
            in3 => \N__21364\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_4_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21333\,
            in1 => \N__21309\,
            in2 => \N__21272\,
            in3 => \N__21269\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_6_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25228\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47619\,
            ce => 'H',
            sr => \N__46917\
        );

    \current_shift_inst.PI_CTRL.prop_term_8_LC_4_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25159\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47619\,
            ce => 'H',
            sr => \N__46917\
        );

    \current_shift_inst.PI_CTRL.prop_term_5_LC_4_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25261\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47619\,
            ce => 'H',
            sr => \N__46917\
        );

    \current_shift_inst.PI_CTRL.prop_term_7_LC_4_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25195\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47619\,
            ce => 'H',
            sr => \N__46917\
        );

    \current_shift_inst.PI_CTRL.prop_term_13_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25531\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47607\,
            ce => 'H',
            sr => \N__46921\
        );

    \current_shift_inst.PI_CTRL.prop_term_11_LC_4_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25597\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47607\,
            ce => 'H',
            sr => \N__46921\
        );

    \current_shift_inst.PI_CTRL.prop_term_9_LC_4_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25132\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47607\,
            ce => 'H',
            sr => \N__46921\
        );

    \current_shift_inst.PI_CTRL.prop_term_12_LC_4_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25567\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47607\,
            ce => 'H',
            sr => \N__46921\
        );

    \current_shift_inst.PI_CTRL.prop_term_1_LC_4_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25385\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47607\,
            ce => 'H',
            sr => \N__46921\
        );

    \current_shift_inst.PI_CTRL.prop_term_4_LC_4_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25294\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47607\,
            ce => 'H',
            sr => \N__46921\
        );

    \current_shift_inst.PI_CTRL.prop_term_10_LC_4_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25627\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47598\,
            ce => 'H',
            sr => \N__46926\
        );

    \current_shift_inst.PI_CTRL.prop_term_14_LC_4_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25442\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47598\,
            ce => 'H',
            sr => \N__46926\
        );

    \pwm_generator_inst.un3_threshold_axb_4_LC_4_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21962\,
            in2 => \N__21947\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un3_threshold_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \bfn_4_23_0_\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_4_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21926\,
            in2 => \N__21908\,
            in3 => \N__21884\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_0\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_4_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21881\,
            in2 => \N__21866\,
            in3 => \N__21845\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_1\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_4_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21842\,
            in2 => \N__21827\,
            in3 => \N__21803\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_2\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_4_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21800\,
            in2 => \N__21788\,
            in3 => \N__21761\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_3\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_4_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21758\,
            in2 => \N__21746\,
            in3 => \N__21719\,
            lcout => \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_4\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_4_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21716\,
            in2 => \N__21704\,
            in3 => \N__21680\,
            lcout => \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_5\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_4_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22274\,
            in2 => \N__22262\,
            in3 => \N__22235\,
            lcout => \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_6\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_4_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22232\,
            in2 => \N__22217\,
            in3 => \N__22196\,
            lcout => \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \bfn_4_24_0_\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_4_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22193\,
            in2 => \N__22175\,
            in3 => \N__22154\,
            lcout => \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_8\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_4_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22151\,
            in2 => \N__46071\,
            in3 => \N__22130\,
            lcout => \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_9\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_4_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22127\,
            in2 => \N__46073\,
            in3 => \N__22106\,
            lcout => \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_10\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_4_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22103\,
            in2 => \N__46072\,
            in3 => \N__22079\,
            lcout => \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_11\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_4_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22076\,
            in2 => \N__46074\,
            in3 => \N__22052\,
            lcout => \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_12\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_4_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46064\,
            in2 => \N__22352\,
            in3 => \N__22328\,
            lcout => \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_13\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_4_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46057\,
            in2 => \N__46010\,
            in3 => \N__22313\,
            lcout => \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_14\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_4_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23456\,
            in1 => \N__22310\,
            in2 => \_gnd_net_\,
            in3 => \N__22304\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\,
            ltout => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_4_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110001011100"
        )
    port map (
            in0 => \N__23801\,
            in1 => \N__22420\,
            in2 => \N__22301\,
            in3 => \N__23818\,
            lcout => \pwm_generator_inst.un19_threshold_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_4_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__23741\,
            in1 => \N__23758\,
            in2 => \N__22385\,
            in3 => \N__24011\,
            lcout => \pwm_generator_inst.un19_threshold_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_4_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__23419\,
            in1 => \N__23768\,
            in2 => \N__23792\,
            in3 => \N__24010\,
            lcout => \pwm_generator_inst.un19_threshold_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_4_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110001011100"
        )
    port map (
            in0 => \N__23693\,
            in1 => \N__22399\,
            in2 => \N__24030\,
            in3 => \N__23710\,
            lcout => \pwm_generator_inst.un19_threshold_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_4_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__23543\,
            in1 => \N__23569\,
            in2 => \N__22298\,
            in3 => \N__24009\,
            lcout => \pwm_generator_inst.un19_threshold_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_4_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22435\,
            in2 => \_gnd_net_\,
            in3 => \N__23732\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_16\,
            ltout => \pwm_generator_inst.un15_threshold_1_axb_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_4_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__22436\,
            in1 => \N__24019\,
            in2 => \N__22424\,
            in3 => \N__23720\,
            lcout => \pwm_generator_inst.un19_threshold_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_4_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__23509\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23443\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_4_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22421\,
            in2 => \_gnd_net_\,
            in3 => \N__23819\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_4_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22400\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23711\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_4_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22384\,
            in2 => \_gnd_net_\,
            in3 => \N__23759\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_4_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24079\,
            in2 => \_gnd_net_\,
            in3 => \N__24100\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.running_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111110000"
        )
    port map (
            in0 => \N__23918\,
            in1 => \N__24913\,
            in2 => \N__22367\,
            in3 => \N__32368\,
            lcout => \phase_controller_inst1.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47685\,
            ce => 'H',
            sr => \N__46878\
        );

    \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__23915\,
            in1 => \N__22363\,
            in2 => \_gnd_net_\,
            in3 => \N__33763\,
            lcout => \phase_controller_inst1.stoper_hc.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__23916\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33764\,
            lcout => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101000001010"
        )
    port map (
            in0 => \N__34588\,
            in1 => \N__24914\,
            in2 => \N__32377\,
            in3 => \N__23917\,
            lcout => \phase_controller_inst1.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47665\,
            ce => 'H',
            sr => \N__46889\
        );

    \current_shift_inst.PI_CTRL.integrator_9_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000001010001"
        )
    port map (
            in0 => \N__23253\,
            in1 => \N__23050\,
            in2 => \N__23306\,
            in3 => \N__22565\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47643\,
            ce => 'H',
            sr => \N__46900\
        );

    \current_shift_inst.PI_CTRL.integrator_7_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000001010001"
        )
    port map (
            in0 => \N__23252\,
            in1 => \N__23049\,
            in2 => \N__22931\,
            in3 => \N__22564\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47643\,
            ce => 'H',
            sr => \N__46900\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__22869\,
            in1 => \N__22832\,
            in2 => \N__22793\,
            in3 => \N__22748\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_44_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22731\,
            in1 => \N__22699\,
            in2 => \N__22670\,
            in3 => \N__22667\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_5_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22661\,
            in1 => \N__22655\,
            in2 => \N__22649\,
            in3 => \N__22640\,
            lcout => \current_shift_inst.PI_CTRL.N_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_3_LC_5_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25324\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47608\,
            ce => 'H',
            sr => \N__46912\
        );

    \current_shift_inst.PI_CTRL.prop_term_2_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25354\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47608\,
            ce => 'H',
            sr => \N__46912\
        );

    \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_5_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__46283\,
            in1 => \N__23477\,
            in2 => \N__46208\,
            in3 => \N__46075\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_5_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__23489\,
            in1 => \N__23510\,
            in2 => \N__23444\,
            in3 => \N__24018\,
            lcout => \pwm_generator_inst.un19_threshold_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_5_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23420\,
            in2 => \_gnd_net_\,
            in3 => \N__23790\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_5_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23390\,
            in2 => \_gnd_net_\,
            in3 => \N__23405\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_5_25_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_5_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23369\,
            in2 => \_gnd_net_\,
            in3 => \N__23384\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_0\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_5_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23351\,
            in2 => \_gnd_net_\,
            in3 => \N__23363\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_1\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_5_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23333\,
            in2 => \_gnd_net_\,
            in3 => \N__23345\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_2\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_5_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23312\,
            in2 => \_gnd_net_\,
            in3 => \N__23327\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_3\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_5_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23660\,
            in2 => \_gnd_net_\,
            in3 => \N__23675\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_4\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_5_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23639\,
            in2 => \_gnd_net_\,
            in3 => \N__23654\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_5\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_5_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23618\,
            in2 => \_gnd_net_\,
            in3 => \N__23633\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_6\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_5_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23597\,
            in2 => \_gnd_net_\,
            in3 => \N__23612\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_8\,
            ltout => OPEN,
            carryin => \bfn_5_26_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_5_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23576\,
            in2 => \_gnd_net_\,
            in3 => \N__23591\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_8\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_5_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23570\,
            in2 => \_gnd_net_\,
            in3 => \N__23537\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_9\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_5_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__24031\,
            in1 => \N__23534\,
            in2 => \_gnd_net_\,
            in3 => \N__23513\,
            lcout => \pwm_generator_inst.un19_threshold_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_10\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_5_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23505\,
            in2 => \_gnd_net_\,
            in3 => \N__23480\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_11\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_5_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23817\,
            in2 => \_gnd_net_\,
            in3 => \N__23795\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_12\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_5_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23791\,
            in2 => \_gnd_net_\,
            in3 => \N__23762\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_13\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_5_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23757\,
            in2 => \_gnd_net_\,
            in3 => \N__23735\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_14\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_5_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23731\,
            in2 => \_gnd_net_\,
            in3 => \N__23714\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_5_27_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_5_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23709\,
            in2 => \_gnd_net_\,
            in3 => \N__23684\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_16\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_5_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24099\,
            in2 => \_gnd_net_\,
            in3 => \N__23681\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_17\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_5_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23678\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27207\,
            in1 => \N__29008\,
            in2 => \_gnd_net_\,
            in3 => \N__31993\,
            lcout => \elapsed_time_ns_1_RNI36DN9_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__26980\,
            in1 => \N__31989\,
            in2 => \_gnd_net_\,
            in3 => \N__26960\,
            lcout => \elapsed_time_ns_1_RNIDV2T9_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31992\,
            in1 => \N__26100\,
            in2 => \_gnd_net_\,
            in3 => \N__26077\,
            lcout => \elapsed_time_ns_1_RNIE03T9_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26041\,
            in1 => \N__27751\,
            in2 => \_gnd_net_\,
            in3 => \N__31991\,
            lcout => \elapsed_time_ns_1_RNIF13T9_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31990\,
            in1 => \N__26184\,
            in2 => \_gnd_net_\,
            in3 => \N__27683\,
            lcout => \elapsed_time_ns_1_RNIG23T9_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_25_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27208\,
            in1 => \N__29007\,
            in2 => \_gnd_net_\,
            in3 => \N__31995\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47686\,
            ce => \N__32574\,
            sr => \N__46859\
        );

    \phase_controller_inst1.stoper_hc.target_time_1_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26958\,
            in1 => \N__26976\,
            in2 => \_gnd_net_\,
            in3 => \N__31994\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47686\,
            ce => \N__32574\,
            sr => \N__46859\
        );

    \phase_controller_inst1.stoper_hc.target_time_3_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26037\,
            in1 => \N__27752\,
            in2 => \_gnd_net_\,
            in3 => \N__31996\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47686\,
            ce => \N__32574\,
            sr => \N__46859\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011100110001"
        )
    port map (
            in0 => \N__24346\,
            in1 => \N__24315\,
            in2 => \N__25019\,
            in3 => \N__23953\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__27607\,
            in1 => \N__31939\,
            in2 => \_gnd_net_\,
            in3 => \N__26014\,
            lcout => \elapsed_time_ns_1_RNIH33T9_0_5\,
            ltout => \elapsed_time_ns_1_RNIH33T9_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_5_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__31940\,
            in1 => \_gnd_net_\,
            in2 => \N__23822\,
            in3 => \N__27608\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47675\,
            ce => \N__32654\,
            sr => \N__46864\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001100010000"
        )
    port map (
            in0 => \N__24403\,
            in1 => \N__24379\,
            in2 => \N__25034\,
            in3 => \N__23837\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100101011"
        )
    port map (
            in0 => \N__23836\,
            in1 => \N__24404\,
            in2 => \N__24383\,
            in3 => \N__25030\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_21_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31941\,
            in1 => \N__31453\,
            in2 => \_gnd_net_\,
            in3 => \N__31420\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47666\,
            ce => \N__32655\,
            sr => \N__46869\
        );

    \phase_controller_inst1.stoper_hc.target_time_2_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31942\,
            in1 => \N__26102\,
            in2 => \_gnd_net_\,
            in3 => \N__26073\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47666\,
            ce => \N__32655\,
            sr => \N__46869\
        );

    \phase_controller_inst1.stoper_hc.target_time_RNIO0241_0_30_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010001110"
        )
    port map (
            in0 => \N__26331\,
            in1 => \N__24513\,
            in2 => \N__23940\,
            in3 => \N__24540\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3_28_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32373\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32395\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_RNIO0241_30_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__26332\,
            in1 => \N__24514\,
            in2 => \N__23941\,
            in3 => \N__24541\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un4_running_df30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI4E6P2_28_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110101011101"
        )
    port map (
            in0 => \N__23903\,
            in1 => \N__24937\,
            in2 => \N__23828\,
            in3 => \N__24926\,
            lcout => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23825\,
            in3 => \N__32372\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011001111"
        )
    port map (
            in0 => \N__26333\,
            in1 => \N__24515\,
            in2 => \N__23942\,
            in3 => \N__24542\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26945\,
            in1 => \N__27735\,
            in2 => \N__27677\,
            in3 => \N__26060\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111100000100"
        )
    port map (
            in0 => \N__24350\,
            in1 => \N__25012\,
            in2 => \N__24323\,
            in3 => \N__23957\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_31_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28718\,
            in1 => \N__27817\,
            in2 => \_gnd_net_\,
            in3 => \N__31959\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47630\,
            ce => \N__32653\,
            sr => \N__46884\
        );

    \phase_controller_inst1.state_4_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30811\,
            in2 => \_gnd_net_\,
            in3 => \N__34661\,
            lcout => phase_controller_inst1_state_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47609\,
            ce => 'H',
            sr => \N__46894\
        );

    \phase_controller_inst1.stoper_hc.start_latched_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33762\,
            lcout => \phase_controller_inst1.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47590\,
            ce => 'H',
            sr => \N__46904\
        );

    \delay_measurement_inst.delay_hc_timer.running_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__29277\,
            in1 => \N__32963\,
            in2 => \_gnd_net_\,
            in3 => \N__30920\,
            lcout => \delay_measurement_inst.delay_hc_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47590\,
            ce => 'H',
            sr => \N__46904\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_7_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23879\,
            in2 => \N__24054\,
            in3 => \N__24053\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93\,
            ltout => OPEN,
            carryin => \bfn_7_23_0_\,
            carryout => \pwm_generator_inst.un19_threshold_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_7_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23867\,
            in2 => \_gnd_net_\,
            in3 => \N__23855\,
            lcout => \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_0\,
            carryout => \pwm_generator_inst.un19_threshold_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_7_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23852\,
            in2 => \_gnd_net_\,
            in3 => \N__23840\,
            lcout => \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_1\,
            carryout => \pwm_generator_inst.un19_threshold_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_7_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24209\,
            in2 => \_gnd_net_\,
            in3 => \N__24197\,
            lcout => \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_2\,
            carryout => \pwm_generator_inst.un19_threshold_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_7_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24194\,
            in2 => \_gnd_net_\,
            in3 => \N__24182\,
            lcout => \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_3\,
            carryout => \pwm_generator_inst.un19_threshold_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_7_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24179\,
            in2 => \_gnd_net_\,
            in3 => \N__24167\,
            lcout => \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_4\,
            carryout => \pwm_generator_inst.un19_threshold_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_7_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24164\,
            in2 => \_gnd_net_\,
            in3 => \N__24152\,
            lcout => \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_5\,
            carryout => \pwm_generator_inst.un19_threshold_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_7_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24149\,
            in2 => \_gnd_net_\,
            in3 => \N__24137\,
            lcout => \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_6\,
            carryout => \pwm_generator_inst.un19_threshold_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_7_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23963\,
            in2 => \_gnd_net_\,
            in3 => \N__24134\,
            lcout => \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033\,
            ltout => OPEN,
            carryin => \bfn_7_24_0_\,
            carryout => \pwm_generator_inst.un19_threshold_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_7_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__24131\,
            in1 => \N__24119\,
            in2 => \N__24056\,
            in3 => \N__24107\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_7_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110001011100"
        )
    port map (
            in0 => \N__24104\,
            in1 => \N__24080\,
            in2 => \N__24055\,
            in3 => \N__23975\,
            lcout => \pwm_generator_inst.un19_threshold_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D1_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24266\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_max_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47702\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101000101"
        )
    port map (
            in0 => \N__25954\,
            in1 => \N__25903\,
            in2 => \N__25931\,
            in3 => \N__25888\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24257\,
            in2 => \N__32342\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_5_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32659\,
            in1 => \N__24469\,
            in2 => \_gnd_net_\,
            in3 => \N__24242\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \N__47698\,
            ce => 'H',
            sr => \N__46835\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__32598\,
            in1 => \N__24439\,
            in2 => \N__24239\,
            in3 => \N__24224\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \N__47698\,
            ce => 'H',
            sr => \N__46835\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32660\,
            in1 => \N__24724\,
            in2 => \_gnd_net_\,
            in3 => \N__24221\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \N__47698\,
            ce => 'H',
            sr => \N__46835\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32599\,
            in1 => \N__24700\,
            in2 => \_gnd_net_\,
            in3 => \N__24218\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \N__47698\,
            ce => 'H',
            sr => \N__46835\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32661\,
            in1 => \N__24670\,
            in2 => \_gnd_net_\,
            in3 => \N__24215\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \N__47698\,
            ce => 'H',
            sr => \N__46835\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32600\,
            in1 => \N__24649\,
            in2 => \_gnd_net_\,
            in3 => \N__24212\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \N__47698\,
            ce => 'H',
            sr => \N__46835\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32662\,
            in1 => \N__24625\,
            in2 => \_gnd_net_\,
            in3 => \N__24293\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \N__47698\,
            ce => 'H',
            sr => \N__46835\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32670\,
            in1 => \N__24601\,
            in2 => \_gnd_net_\,
            in3 => \N__24290\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_8_6_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \N__47695\,
            ce => 'H',
            sr => \N__46842\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32609\,
            in1 => \N__24577\,
            in2 => \_gnd_net_\,
            in3 => \N__24287\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \N__47695\,
            ce => 'H',
            sr => \N__46842\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32667\,
            in1 => \N__24880\,
            in2 => \_gnd_net_\,
            in3 => \N__24284\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \N__47695\,
            ce => 'H',
            sr => \N__46842\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32610\,
            in1 => \N__24853\,
            in2 => \_gnd_net_\,
            in3 => \N__24281\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \N__47695\,
            ce => 'H',
            sr => \N__46842\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32668\,
            in1 => \N__24829\,
            in2 => \_gnd_net_\,
            in3 => \N__24278\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \N__47695\,
            ce => 'H',
            sr => \N__46842\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32611\,
            in1 => \N__24802\,
            in2 => \_gnd_net_\,
            in3 => \N__24275\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \N__47695\,
            ce => 'H',
            sr => \N__46842\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32669\,
            in1 => \N__24781\,
            in2 => \_gnd_net_\,
            in3 => \N__24272\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \N__47695\,
            ce => 'H',
            sr => \N__46842\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32612\,
            in1 => \N__25927\,
            in2 => \_gnd_net_\,
            in3 => \N__24269\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \N__47695\,
            ce => 'H',
            sr => \N__46842\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32605\,
            in1 => \N__25953\,
            in2 => \_gnd_net_\,
            in3 => \N__24413\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_8_7_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \N__47687\,
            ce => 'H',
            sr => \N__46847\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32663\,
            in1 => \N__25823\,
            in2 => \_gnd_net_\,
            in3 => \N__24410\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \N__47687\,
            ce => 'H',
            sr => \N__46847\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32606\,
            in1 => \N__25838\,
            in2 => \_gnd_net_\,
            in3 => \N__24407\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \N__47687\,
            ce => 'H',
            sr => \N__46847\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32664\,
            in1 => \N__24402\,
            in2 => \_gnd_net_\,
            in3 => \N__24386\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \N__47687\,
            ce => 'H',
            sr => \N__46847\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32607\,
            in1 => \N__24373\,
            in2 => \_gnd_net_\,
            in3 => \N__24359\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\,
            clk => \N__47687\,
            ce => 'H',
            sr => \N__46847\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32665\,
            in1 => \N__25970\,
            in2 => \_gnd_net_\,
            in3 => \N__24356\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\,
            clk => \N__47687\,
            ce => 'H',
            sr => \N__46847\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32608\,
            in1 => \N__25987\,
            in2 => \_gnd_net_\,
            in3 => \N__24353\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\,
            clk => \N__47687\,
            ce => 'H',
            sr => \N__46847\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32666\,
            in1 => \N__24345\,
            in2 => \_gnd_net_\,
            in3 => \N__24326\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\,
            clk => \N__47687\,
            ce => 'H',
            sr => \N__46847\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32552\,
            in1 => \N__24316\,
            in2 => \_gnd_net_\,
            in3 => \N__24296\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\,
            clk => \N__47676\,
            ce => 'H',
            sr => \N__46853\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32571\,
            in1 => \N__25071\,
            in2 => \_gnd_net_\,
            in3 => \N__24554\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\,
            clk => \N__47676\,
            ce => 'H',
            sr => \N__46853\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32553\,
            in1 => \N__25092\,
            in2 => \_gnd_net_\,
            in3 => \N__24551\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\,
            clk => \N__47676\,
            ce => 'H',
            sr => \N__46853\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32572\,
            in1 => \N__30981\,
            in2 => \_gnd_net_\,
            in3 => \N__24548\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\,
            clk => \N__47676\,
            ce => 'H',
            sr => \N__46853\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32554\,
            in1 => \N__30957\,
            in2 => \_gnd_net_\,
            in3 => \N__24545\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\,
            clk => \N__47676\,
            ce => 'H',
            sr => \N__46853\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32573\,
            in1 => \N__24539\,
            in2 => \_gnd_net_\,
            in3 => \N__24521\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\,
            clk => \N__47676\,
            ce => 'H',
            sr => \N__46853\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32555\,
            in1 => \N__24512\,
            in2 => \_gnd_net_\,
            in3 => \N__24518\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47676\,
            ce => 'H',
            sr => \N__46853\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24491\,
            in2 => \N__24485\,
            in3 => \N__32335\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_8_9_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24476\,
            in2 => \N__24455\,
            in3 => \N__24470\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24446\,
            in2 => \N__24425\,
            in3 => \N__24440\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26165\,
            in2 => \N__24710\,
            in3 => \N__24728\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24701\,
            in1 => \N__24677\,
            in2 => \N__24686\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24671\,
            in1 => \N__24656\,
            in2 => \N__26300\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24650\,
            in1 => \N__31532\,
            in2 => \N__24635\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24626\,
            in1 => \N__25046\,
            in2 => \N__24611\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_7\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24602\,
            in1 => \N__26234\,
            in2 => \N__24587\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_8_10_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26249\,
            in2 => \N__24563\,
            in3 => \N__24578\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26339\,
            in2 => \N__24866\,
            in3 => \N__24881\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26285\,
            in2 => \N__24839\,
            in3 => \N__24857\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26315\,
            in2 => \N__24815\,
            in3 => \N__24830\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24803\,
            in1 => \N__24788\,
            in2 => \N__27041\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24782\,
            in1 => \N__25790\,
            in2 => \N__24767\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24755\,
            in2 => \N__25877\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_15\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25862\,
            in2 => \N__25808\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_11_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24743\,
            in2 => \N__24737\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26228\,
            in2 => \N__26003\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24968\,
            in2 => \N__24962\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24887\,
            in2 => \N__25055\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30932\,
            in2 => \N__31064\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24950\,
            in2 => \N__24944\,
            in3 => \N__24920\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24917\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28903\,
            in1 => \N__31764\,
            in2 => \_gnd_net_\,
            in3 => \N__27391\,
            lcout => \elapsed_time_ns_1_RNI58DN9_0_27\,
            ltout => \elapsed_time_ns_1_RNI58DN9_0_27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_27_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__31765\,
            in1 => \_gnd_net_\,
            in2 => \N__24890\,
            in3 => \N__28904\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47631\,
            ce => \N__32647\,
            sr => \N__46873\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__26308\,
            in1 => \N__25093\,
            in2 => \N__25076\,
            in3 => \N__25105\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010001110"
        )
    port map (
            in0 => \N__25106\,
            in1 => \N__26309\,
            in2 => \N__25097\,
            in3 => \N__25075\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_8_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31770\,
            in1 => \N__29424\,
            in2 => \_gnd_net_\,
            in3 => \N__29408\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47620\,
            ce => \N__32652\,
            sr => \N__46879\
        );

    \phase_controller_inst1.stoper_hc.target_time_20_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31565\,
            in1 => \N__32040\,
            in2 => \_gnd_net_\,
            in3 => \N__31771\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47620\,
            ce => \N__32652\,
            sr => \N__46879\
        );

    \phase_controller_inst1.stoper_hc.target_time_24_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31769\,
            in1 => \N__26913\,
            in2 => \_gnd_net_\,
            in3 => \N__29075\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47620\,
            ce => \N__32652\,
            sr => \N__46879\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27772\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47610\,
            ce => \N__28683\,
            sr => \N__46885\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27703\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47599\,
            ce => \N__28671\,
            sr => \N__46890\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29276\,
            in2 => \_gnd_net_\,
            in3 => \N__30919\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_202_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_0_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29126\,
            in2 => \_gnd_net_\,
            in3 => \N__29300\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47584\,
            ce => 'H',
            sr => \N__46901\
        );

    \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26504\,
            in1 => \N__24974\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axb_0\,
            ltout => OPEN,
            carryin => \bfn_8_19_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_1_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26498\,
            in2 => \_gnd_net_\,
            in3 => \N__25358\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            clk => \N__47574\,
            ce => 'H',
            sr => \N__46908\
        );

    \current_shift_inst.PI_CTRL.error_control_2_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26489\,
            in2 => \_gnd_net_\,
            in3 => \N__25328\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            clk => \N__47574\,
            ce => 'H',
            sr => \N__46908\
        );

    \current_shift_inst.PI_CTRL.error_control_3_LC_8_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26594\,
            in2 => \_gnd_net_\,
            in3 => \N__25298\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            clk => \N__47574\,
            ce => 'H',
            sr => \N__46908\
        );

    \current_shift_inst.PI_CTRL.error_control_4_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26585\,
            in2 => \_gnd_net_\,
            in3 => \N__25268\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            clk => \N__47574\,
            ce => 'H',
            sr => \N__46908\
        );

    \current_shift_inst.PI_CTRL.error_control_5_LC_8_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26576\,
            in2 => \_gnd_net_\,
            in3 => \N__25235\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            clk => \N__47574\,
            ce => 'H',
            sr => \N__46908\
        );

    \current_shift_inst.PI_CTRL.error_control_6_LC_8_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26567\,
            in2 => \_gnd_net_\,
            in3 => \N__25202\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            clk => \N__47574\,
            ce => 'H',
            sr => \N__46908\
        );

    \current_shift_inst.PI_CTRL.error_control_7_LC_8_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26558\,
            in2 => \_gnd_net_\,
            in3 => \N__25169\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            clk => \N__47574\,
            ce => 'H',
            sr => \N__46908\
        );

    \current_shift_inst.PI_CTRL.error_control_8_LC_8_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26549\,
            in2 => \_gnd_net_\,
            in3 => \N__25139\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_8\,
            ltout => OPEN,
            carryin => \bfn_8_20_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            clk => \N__47569\,
            ce => 'H',
            sr => \N__46913\
        );

    \current_shift_inst.PI_CTRL.error_control_9_LC_8_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26540\,
            in2 => \_gnd_net_\,
            in3 => \N__25634\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            clk => \N__47569\,
            ce => 'H',
            sr => \N__46913\
        );

    \current_shift_inst.PI_CTRL.error_control_10_LC_8_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26531\,
            in2 => \_gnd_net_\,
            in3 => \N__25601\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            clk => \N__47569\,
            ce => 'H',
            sr => \N__46913\
        );

    \current_shift_inst.PI_CTRL.error_control_11_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26708\,
            in2 => \_gnd_net_\,
            in3 => \N__25571\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            clk => \N__47569\,
            ce => 'H',
            sr => \N__46913\
        );

    \current_shift_inst.PI_CTRL.error_control_12_LC_8_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26699\,
            in2 => \_gnd_net_\,
            in3 => \N__25541\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            clk => \N__47569\,
            ce => 'H',
            sr => \N__46913\
        );

    \current_shift_inst.PI_CTRL.error_control_13_LC_8_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26675\,
            in2 => \_gnd_net_\,
            in3 => \N__25505\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_13\,
            clk => \N__47569\,
            ce => 'H',
            sr => \N__46913\
        );

    \current_shift_inst.PI_CTRL.error_control_14_LC_8_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26687\,
            in2 => \_gnd_net_\,
            in3 => \N__25502\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47569\,
            ce => 'H',
            sr => \N__46913\
        );

    \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_8_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110101"
        )
    port map (
            in0 => \N__25690\,
            in1 => \N__25735\,
            in2 => \N__25412\,
            in3 => \N__46169\,
            lcout => \pwm_generator_inst.un14_counter_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_8_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110011"
        )
    port map (
            in0 => \N__25736\,
            in1 => \N__25691\,
            in2 => \N__25403\,
            in3 => \N__46249\,
            lcout => \pwm_generator_inst.un14_counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_8_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011000000"
        )
    port map (
            in0 => \N__25734\,
            in1 => \N__25689\,
            in2 => \N__25394\,
            in3 => \N__46248\,
            lcout => \pwm_generator_inst.threshold_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_8_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011000000"
        )
    port map (
            in0 => \N__25733\,
            in1 => \N__25688\,
            in2 => \N__25778\,
            in3 => \N__46247\,
            lcout => \pwm_generator_inst.threshold_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_8_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111111101"
        )
    port map (
            in0 => \N__25687\,
            in1 => \N__25769\,
            in2 => \N__46255\,
            in3 => \N__25732\,
            lcout => \pwm_generator_inst.un14_counter_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_8_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010011"
        )
    port map (
            in0 => \N__25719\,
            in1 => \N__25685\,
            in2 => \N__46259\,
            in3 => \N__25763\,
            lcout => \pwm_generator_inst.un14_counter_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_8_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010000000"
        )
    port map (
            in0 => \N__25720\,
            in1 => \N__46243\,
            in2 => \N__25757\,
            in3 => \N__25686\,
            lcout => \pwm_generator_inst.threshold_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_8_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__25684\,
            in1 => \N__25748\,
            in2 => \N__46254\,
            in3 => \N__25718\,
            lcout => \pwm_generator_inst.threshold_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_8_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__25682\,
            in1 => \N__25742\,
            in2 => \N__46253\,
            in3 => \N__25716\,
            lcout => \pwm_generator_inst.threshold_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_8_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011000000"
        )
    port map (
            in0 => \N__25717\,
            in1 => \N__25683\,
            in2 => \N__25643\,
            in3 => \N__46242\,
            lcout => \pwm_generator_inst.threshold_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_16_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29730\,
            in1 => \N__29713\,
            in2 => \_gnd_net_\,
            in3 => \N__31911\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47701\,
            ce => \N__32657\,
            sr => \N__46812\
        );

    \phase_controller_inst1.stoper_hc.target_time_17_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26895\,
            in1 => \N__28571\,
            in2 => \_gnd_net_\,
            in3 => \N__32009\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47699\,
            ce => \N__32658\,
            sr => \N__46821\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100010000"
        )
    port map (
            in0 => \N__25955\,
            in1 => \N__25926\,
            in2 => \N__25907\,
            in3 => \N__25889\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31969\,
            in1 => \N__26897\,
            in2 => \_gnd_net_\,
            in3 => \N__28569\,
            lcout => \elapsed_time_ns_1_RNI46CN9_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26851\,
            in1 => \N__27910\,
            in2 => \_gnd_net_\,
            in3 => \N__31968\,
            lcout => \elapsed_time_ns_1_RNI13CN9_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__25847\,
            in1 => \N__25837\,
            in2 => \N__27059\,
            in3 => \N__25822\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__31965\,
            in1 => \N__28503\,
            in2 => \_gnd_net_\,
            in3 => \N__27004\,
            lcout => \elapsed_time_ns_1_RNI57CN9_0_18\,
            ltout => \elapsed_time_ns_1_RNI57CN9_0_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_18_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011100010111000"
        )
    port map (
            in0 => \N__28504\,
            in1 => \N__31967\,
            in2 => \N__25850\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47688\,
            ce => \N__32671\,
            sr => \N__46836\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__25846\,
            in1 => \N__25836\,
            in2 => \N__27058\,
            in3 => \N__25821\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__31963\,
            in1 => \N__29619\,
            in2 => \_gnd_net_\,
            in3 => \N__29584\,
            lcout => \elapsed_time_ns_1_RNI24CN9_0_15\,
            ltout => \elapsed_time_ns_1_RNI24CN9_0_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_15_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011100010111000"
        )
    port map (
            in0 => \N__29620\,
            in1 => \N__31966\,
            in2 => \N__25793\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47688\,
            ce => \N__32671\,
            sr => \N__46836\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31964\,
            in1 => \N__27079\,
            in2 => \_gnd_net_\,
            in3 => \N__28435\,
            lcout => \elapsed_time_ns_1_RNI68CN9_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__30115\,
            in1 => \N__26993\,
            in2 => \N__26114\,
            in3 => \N__30415\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__26992\,
            in1 => \N__30116\,
            in2 => \N__30419\,
            in3 => \N__26110\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_19_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27075\,
            in1 => \N__31972\,
            in2 => \_gnd_net_\,
            in3 => \N__28433\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47677\,
            ce => \N__31312\,
            sr => \N__46843\
        );

    \phase_controller_inst2.stoper_hc.target_time_2_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31970\,
            in1 => \N__26101\,
            in2 => \_gnd_net_\,
            in3 => \N__26078\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47677\,
            ce => \N__31312\,
            sr => \N__46843\
        );

    \phase_controller_inst2.stoper_hc.target_time_3_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__26042\,
            in1 => \N__31973\,
            in2 => \_gnd_net_\,
            in3 => \N__27750\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47677\,
            ce => \N__31312\,
            sr => \N__46843\
        );

    \phase_controller_inst2.stoper_hc.target_time_4_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31971\,
            in1 => \N__26185\,
            in2 => \_gnd_net_\,
            in3 => \N__27681\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47677\,
            ce => \N__31312\,
            sr => \N__46843\
        );

    \phase_controller_inst2.stoper_hc.target_time_5_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__27606\,
            in1 => \N__31974\,
            in2 => \_gnd_net_\,
            in3 => \N__26021\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47677\,
            ce => \N__31312\,
            sr => \N__46843\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__25969\,
            in1 => \N__26198\,
            in2 => \N__26213\,
            in3 => \N__25986\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011001111"
        )
    port map (
            in0 => \N__26197\,
            in1 => \N__26209\,
            in2 => \N__25988\,
            in3 => \N__25968\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28248\,
            in1 => \N__26137\,
            in2 => \_gnd_net_\,
            in3 => \N__31907\,
            lcout => \elapsed_time_ns_1_RNI14DN9_0_23\,
            ltout => \elapsed_time_ns_1_RNI14DN9_0_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_23_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__31909\,
            in1 => \_gnd_net_\,
            in2 => \N__26216\,
            in3 => \N__28249\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47667\,
            ce => \N__32601\,
            sr => \N__46848\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28305\,
            in1 => \N__31906\,
            in2 => \_gnd_net_\,
            in3 => \N__26158\,
            lcout => \elapsed_time_ns_1_RNI03DN9_0_22\,
            ltout => \elapsed_time_ns_1_RNI03DN9_0_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_22_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__31908\,
            in1 => \_gnd_net_\,
            in2 => \N__26201\,
            in3 => \N__28306\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47667\,
            ce => \N__32601\,
            sr => \N__46848\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31910\,
            in1 => \N__26189\,
            in2 => \_gnd_net_\,
            in3 => \N__27682\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47667\,
            ce => \N__32601\,
            sr => \N__46848\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__30359\,
            in1 => \N__30382\,
            in2 => \N__26126\,
            in3 => \N__26147\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__26146\,
            in1 => \N__30358\,
            in2 => \N__30386\,
            in3 => \N__26122\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_22_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__31901\,
            in1 => \N__28307\,
            in2 => \_gnd_net_\,
            in3 => \N__26159\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47654\,
            ce => \N__31311\,
            sr => \N__46854\
        );

    \phase_controller_inst2.stoper_hc.target_time_23_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26138\,
            in1 => \N__28250\,
            in2 => \_gnd_net_\,
            in3 => \N__31903\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47654\,
            ce => \N__31311\,
            sr => \N__46854\
        );

    \phase_controller_inst2.stoper_hc.target_time_11_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31900\,
            in1 => \N__26363\,
            in2 => \_gnd_net_\,
            in3 => \N__28049\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47654\,
            ce => \N__31311\,
            sr => \N__46854\
        );

    \phase_controller_inst2.stoper_hc.target_time_10_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28112\,
            in1 => \N__31902\,
            in2 => \_gnd_net_\,
            in3 => \N__26264\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47654\,
            ce => \N__31311\,
            sr => \N__46854\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28154\,
            in1 => \N__27981\,
            in2 => \N__28111\,
            in3 => \N__28044\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__27597\,
            in1 => \N__27550\,
            in2 => \N__26267\,
            in3 => \N__26243\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__28106\,
            in1 => \_gnd_net_\,
            in2 => \N__31988\,
            in3 => \N__26263\,
            lcout => \elapsed_time_ns_1_RNITUBN9_0_10\,
            ltout => \elapsed_time_ns_1_RNITUBN9_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_10_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28107\,
            in2 => \N__26252\,
            in3 => \N__31898\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47644\,
            ce => \N__32616\,
            sr => \N__46860\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29400\,
            in2 => \_gnd_net_\,
            in3 => \N__31362\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27019\,
            in1 => \N__31894\,
            in2 => \_gnd_net_\,
            in3 => \N__28155\,
            lcout => \elapsed_time_ns_1_RNIL73T9_0_9\,
            ltout => \elapsed_time_ns_1_RNIL73T9_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_9_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__28156\,
            in1 => \_gnd_net_\,
            in2 => \N__26237\,
            in3 => \N__31912\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47644\,
            ce => \N__32616\,
            sr => \N__46860\
        );

    \phase_controller_inst1.stoper_hc.target_time_11_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28045\,
            in1 => \N__26359\,
            in2 => \_gnd_net_\,
            in3 => \N__31899\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47644\,
            ce => \N__32616\,
            sr => \N__46860\
        );

    \phase_controller_inst1.stoper_hc.target_time_30_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27789\,
            in1 => \N__28760\,
            in2 => \_gnd_net_\,
            in3 => \N__31779\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47632\,
            ce => \N__32590\,
            sr => \N__46865\
        );

    \phase_controller_inst1.stoper_hc.target_time_13_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__30470\,
            in1 => \N__31904\,
            in2 => \_gnd_net_\,
            in3 => \N__30443\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47632\,
            ce => \N__32590\,
            sr => \N__46865\
        );

    \phase_controller_inst1.stoper_hc.target_time_26_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30749\,
            in1 => \N__30779\,
            in2 => \_gnd_net_\,
            in3 => \N__31778\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47632\,
            ce => \N__32590\,
            sr => \N__46865\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27549\,
            in1 => \N__26871\,
            in2 => \_gnd_net_\,
            in3 => \N__31780\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47632\,
            ce => \N__32590\,
            sr => \N__46865\
        );

    \phase_controller_inst1.stoper_hc.target_time_12_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27441\,
            in1 => \N__27983\,
            in2 => \_gnd_net_\,
            in3 => \N__31777\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47632\,
            ce => \N__32590\,
            sr => \N__46865\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__28709\,
            in1 => \N__26279\,
            in2 => \N__26372\,
            in3 => \N__26387\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__31446\,
            in1 => \_gnd_net_\,
            in2 => \N__26270\,
            in3 => \N__31413\,
            lcout => \elapsed_time_ns_1_RNIV1DN9_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__27791\,
            in1 => \_gnd_net_\,
            in2 => \N__28758\,
            in3 => \N__31815\,
            lcout => \elapsed_time_ns_1_RNIV2EN9_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__32039\,
            in1 => \N__28483\,
            in2 => \N__28434\,
            in3 => \N__28546\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28710\,
            in1 => \N__27810\,
            in2 => \_gnd_net_\,
            in3 => \N__31814\,
            lcout => \elapsed_time_ns_1_RNI04EN9_0_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28902\,
            in2 => \N__31128\,
            in3 => \N__26396\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26872\,
            in1 => \N__27548\,
            in2 => \_gnd_net_\,
            in3 => \N__31812\,
            lcout => \elapsed_time_ns_1_RNII43T9_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31813\,
            in1 => \N__27445\,
            in2 => \_gnd_net_\,
            in3 => \N__27980\,
            lcout => \elapsed_time_ns_1_RNIV0CN9_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29604\,
            in1 => \N__27894\,
            in2 => \N__29696\,
            in3 => \N__30464\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26420\,
            in1 => \N__26426\,
            in2 => \N__26381\,
            in3 => \N__26378\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__26917\,
            in1 => \N__31748\,
            in2 => \_gnd_net_\,
            in3 => \N__29056\,
            lcout => \elapsed_time_ns_1_RNI25DN9_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__31746\,
            in1 => \N__31121\,
            in2 => \_gnd_net_\,
            in3 => \N__31086\,
            lcout => \elapsed_time_ns_1_RNI69DN9_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__26358\,
            in1 => \N__31749\,
            in2 => \_gnd_net_\,
            in3 => \N__28043\,
            lcout => \elapsed_time_ns_1_RNIUVBN9_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__29428\,
            in1 => \N__31747\,
            in2 => \_gnd_net_\,
            in3 => \N__29396\,
            lcout => \elapsed_time_ns_1_RNIK63T9_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28233\,
            in1 => \N__31409\,
            in2 => \N__28296\,
            in3 => \N__29055\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28739\,
            in1 => \N__30767\,
            in2 => \N__31011\,
            in3 => \N__28983\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.counter_0_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29252\,
            in1 => \N__27768\,
            in2 => \_gnd_net_\,
            in3 => \N__26414\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_9_15_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            clk => \N__47591\,
            ce => \N__29349\,
            sr => \N__46886\
        );

    \delay_measurement_inst.delay_hc_timer.counter_1_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29235\,
            in1 => \N__27702\,
            in2 => \_gnd_net_\,
            in3 => \N__26411\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            clk => \N__47591\,
            ce => \N__29349\,
            sr => \N__46886\
        );

    \delay_measurement_inst.delay_hc_timer.counter_2_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29253\,
            in1 => \N__27627\,
            in2 => \_gnd_net_\,
            in3 => \N__26408\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            clk => \N__47591\,
            ce => \N__29349\,
            sr => \N__46886\
        );

    \delay_measurement_inst.delay_hc_timer.counter_3_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29236\,
            in1 => \N__27570\,
            in2 => \_gnd_net_\,
            in3 => \N__26405\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            clk => \N__47591\,
            ce => \N__29349\,
            sr => \N__46886\
        );

    \delay_measurement_inst.delay_hc_timer.counter_4_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29254\,
            in1 => \N__27513\,
            in2 => \_gnd_net_\,
            in3 => \N__26402\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            clk => \N__47591\,
            ce => \N__29349\,
            sr => \N__46886\
        );

    \delay_measurement_inst.delay_hc_timer.counter_5_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29237\,
            in1 => \N__28206\,
            in2 => \_gnd_net_\,
            in3 => \N__26399\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            clk => \N__47591\,
            ce => \N__29349\,
            sr => \N__46886\
        );

    \delay_measurement_inst.delay_hc_timer.counter_6_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29255\,
            in1 => \N__28176\,
            in2 => \_gnd_net_\,
            in3 => \N__26453\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            clk => \N__47591\,
            ce => \N__29349\,
            sr => \N__46886\
        );

    \delay_measurement_inst.delay_hc_timer.counter_7_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29238\,
            in1 => \N__28126\,
            in2 => \_gnd_net_\,
            in3 => \N__26450\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            clk => \N__47591\,
            ce => \N__29349\,
            sr => \N__46886\
        );

    \delay_measurement_inst.delay_hc_timer.counter_8_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29224\,
            in1 => \N__28071\,
            in2 => \_gnd_net_\,
            in3 => \N__26447\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_9_16_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            clk => \N__47585\,
            ce => \N__29356\,
            sr => \N__46891\
        );

    \delay_measurement_inst.delay_hc_timer.counter_9_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29228\,
            in1 => \N__28005\,
            in2 => \_gnd_net_\,
            in3 => \N__26444\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            clk => \N__47585\,
            ce => \N__29356\,
            sr => \N__46891\
        );

    \delay_measurement_inst.delay_hc_timer.counter_10_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29221\,
            in1 => \N__27951\,
            in2 => \_gnd_net_\,
            in3 => \N__26441\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            clk => \N__47585\,
            ce => \N__29356\,
            sr => \N__46891\
        );

    \delay_measurement_inst.delay_hc_timer.counter_11_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29225\,
            in1 => \N__27925\,
            in2 => \_gnd_net_\,
            in3 => \N__26438\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            clk => \N__47585\,
            ce => \N__29356\,
            sr => \N__46891\
        );

    \delay_measurement_inst.delay_hc_timer.counter_12_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29222\,
            in1 => \N__27870\,
            in2 => \_gnd_net_\,
            in3 => \N__26435\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            clk => \N__47585\,
            ce => \N__29356\,
            sr => \N__46891\
        );

    \delay_measurement_inst.delay_hc_timer.counter_13_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29226\,
            in1 => \N__28617\,
            in2 => \_gnd_net_\,
            in3 => \N__26432\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            clk => \N__47585\,
            ce => \N__29356\,
            sr => \N__46891\
        );

    \delay_measurement_inst.delay_hc_timer.counter_14_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29223\,
            in1 => \N__28587\,
            in2 => \_gnd_net_\,
            in3 => \N__26429\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            clk => \N__47585\,
            ce => \N__29356\,
            sr => \N__46891\
        );

    \delay_measurement_inst.delay_hc_timer.counter_15_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29227\,
            in1 => \N__28521\,
            in2 => \_gnd_net_\,
            in3 => \N__26480\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            clk => \N__47585\,
            ce => \N__29356\,
            sr => \N__46891\
        );

    \delay_measurement_inst.delay_hc_timer.counter_16_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29217\,
            in1 => \N__28458\,
            in2 => \_gnd_net_\,
            in3 => \N__26477\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_9_17_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            clk => \N__47579\,
            ce => \N__29348\,
            sr => \N__46895\
        );

    \delay_measurement_inst.delay_hc_timer.counter_17_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29248\,
            in1 => \N__28377\,
            in2 => \_gnd_net_\,
            in3 => \N__26474\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            clk => \N__47579\,
            ce => \N__29348\,
            sr => \N__46895\
        );

    \delay_measurement_inst.delay_hc_timer.counter_18_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29218\,
            in1 => \N__28350\,
            in2 => \_gnd_net_\,
            in3 => \N__26471\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            clk => \N__47579\,
            ce => \N__29348\,
            sr => \N__46895\
        );

    \delay_measurement_inst.delay_hc_timer.counter_19_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29249\,
            in1 => \N__28323\,
            in2 => \_gnd_net_\,
            in3 => \N__26468\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            clk => \N__47579\,
            ce => \N__29348\,
            sr => \N__46895\
        );

    \delay_measurement_inst.delay_hc_timer.counter_20_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29219\,
            in1 => \N__28266\,
            in2 => \_gnd_net_\,
            in3 => \N__26465\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            clk => \N__47579\,
            ce => \N__29348\,
            sr => \N__46895\
        );

    \delay_measurement_inst.delay_hc_timer.counter_21_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29250\,
            in1 => \N__29094\,
            in2 => \_gnd_net_\,
            in3 => \N__26462\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            clk => \N__47579\,
            ce => \N__29348\,
            sr => \N__46895\
        );

    \delay_measurement_inst.delay_hc_timer.counter_22_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29220\,
            in1 => \N__29025\,
            in2 => \_gnd_net_\,
            in3 => \N__26459\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            clk => \N__47579\,
            ce => \N__29348\,
            sr => \N__46895\
        );

    \delay_measurement_inst.delay_hc_timer.counter_23_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29251\,
            in1 => \N__28956\,
            in2 => \_gnd_net_\,
            in3 => \N__26456\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            clk => \N__47579\,
            ce => \N__29348\,
            sr => \N__46895\
        );

    \delay_measurement_inst.delay_hc_timer.counter_24_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29229\,
            in1 => \N__28926\,
            in2 => \_gnd_net_\,
            in3 => \N__26522\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_9_18_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            clk => \N__47575\,
            ce => \N__29357\,
            sr => \N__46902\
        );

    \delay_measurement_inst.delay_hc_timer.counter_25_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29233\,
            in1 => \N__28863\,
            in2 => \_gnd_net_\,
            in3 => \N__26519\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            clk => \N__47575\,
            ce => \N__29357\,
            sr => \N__46902\
        );

    \delay_measurement_inst.delay_hc_timer.counter_26_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29230\,
            in1 => \N__28839\,
            in2 => \_gnd_net_\,
            in3 => \N__26516\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            clk => \N__47575\,
            ce => \N__29357\,
            sr => \N__46902\
        );

    \delay_measurement_inst.delay_hc_timer.counter_27_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29234\,
            in1 => \N__28782\,
            in2 => \_gnd_net_\,
            in3 => \N__26513\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            clk => \N__47575\,
            ce => \N__29357\,
            sr => \N__46902\
        );

    \delay_measurement_inst.delay_hc_timer.counter_28_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29231\,
            in1 => \N__28819\,
            in2 => \_gnd_net_\,
            in3 => \N__26510\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_28\,
            clk => \N__47575\,
            ce => \N__29357\,
            sr => \N__46902\
        );

    \delay_measurement_inst.delay_hc_timer.counter_29_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__28798\,
            in1 => \N__29232\,
            in2 => \_gnd_net_\,
            in3 => \N__26507\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47575\,
            ce => \N__29357\,
            sr => \N__46902\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29299\,
            in2 => \N__29122\,
            in3 => \N__29118\,
            lcout => \current_shift_inst.control_input_18\,
            ltout => OPEN,
            carryin => \bfn_9_19_0_\,
            carryout => \current_shift_inst.control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33485\,
            in2 => \_gnd_net_\,
            in3 => \N__26492\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_0\,
            carryout => \current_shift_inst.control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33665\,
            in2 => \_gnd_net_\,
            in3 => \N__26483\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_1\,
            carryout => \current_shift_inst.control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33647\,
            in2 => \_gnd_net_\,
            in3 => \N__26588\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_2\,
            carryout => \current_shift_inst.control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33629\,
            in2 => \_gnd_net_\,
            in3 => \N__26579\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_3\,
            carryout => \current_shift_inst.control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33611\,
            in2 => \_gnd_net_\,
            in3 => \N__26570\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_4\,
            carryout => \current_shift_inst.control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33593\,
            in2 => \_gnd_net_\,
            in3 => \N__26561\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_5\,
            carryout => \current_shift_inst.control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33575\,
            in2 => \_gnd_net_\,
            in3 => \N__26552\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_6\,
            carryout => \current_shift_inst.control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33557\,
            in2 => \_gnd_net_\,
            in3 => \N__26543\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_9_20_0_\,
            carryout => \current_shift_inst.control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33833\,
            in2 => \_gnd_net_\,
            in3 => \N__26534\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_8\,
            carryout => \current_shift_inst.control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33815\,
            in2 => \_gnd_net_\,
            in3 => \N__26525\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_9\,
            carryout => \current_shift_inst.control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34481\,
            in2 => \_gnd_net_\,
            in3 => \N__26702\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_10\,
            carryout => \current_shift_inst.control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29132\,
            in2 => \_gnd_net_\,
            in3 => \N__26693\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_11\,
            carryout => \current_shift_inst.control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37634\,
            in2 => \_gnd_net_\,
            in3 => \N__26690\,
            lcout => \current_shift_inst.control_input_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26686\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26657\,
            in2 => \N__26669\,
            in3 => \N__29557\,
            lcout => \pwm_generator_inst.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_9_24_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26642\,
            in2 => \N__26651\,
            in3 => \N__29535\,
            lcout => \pwm_generator_inst.counter_i_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_0\,
            carryout => \pwm_generator_inst.un14_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29514\,
            in1 => \N__26627\,
            in2 => \N__26636\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_1\,
            carryout => \pwm_generator_inst.un14_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_9_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29493\,
            in1 => \N__26612\,
            in2 => \N__26621\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_2\,
            carryout => \pwm_generator_inst.un14_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_9_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29472\,
            in1 => \N__26831\,
            in2 => \N__26606\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_3\,
            carryout => \pwm_generator_inst.un14_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_9_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26813\,
            in2 => \N__26825\,
            in3 => \N__29451\,
            lcout => \pwm_generator_inst.counter_i_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_4\,
            carryout => \pwm_generator_inst.un14_counter_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_9_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29805\,
            in1 => \N__26792\,
            in2 => \N__26807\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_5\,
            carryout => \pwm_generator_inst.un14_counter_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_9_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26777\,
            in2 => \N__26786\,
            in3 => \N__30623\,
            lcout => \pwm_generator_inst.counter_i_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_6\,
            carryout => \pwm_generator_inst.un14_counter_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_9_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30642\,
            in1 => \N__26759\,
            in2 => \N__26771\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_9_25_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_9_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26744\,
            in2 => \N__26753\,
            in3 => \N__30663\,
            lcout => \pwm_generator_inst.counter_i_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_8\,
            carryout => \pwm_generator_inst.un14_counter_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.pwm_out_LC_9_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26738\,
            lcout => pwm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47556\,
            ce => 'H',
            sr => \N__46930\
        );

    \phase_controller_inst2.S1_LC_9_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31178\,
            lcout => s3_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47549\,
            ce => 'H',
            sr => \N__46938\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_10_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29734\,
            in1 => \N__29706\,
            in2 => \_gnd_net_\,
            in3 => \N__32007\,
            lcout => \elapsed_time_ns_1_RNI35CN9_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_19_LC_10_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27080\,
            in1 => \N__28436\,
            in2 => \_gnd_net_\,
            in3 => \N__32008\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47689\,
            ce => \N__32672\,
            sr => \N__46803\
        );

    \phase_controller_inst1.stoper_hc.target_time_14_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26847\,
            in1 => \N__27909\,
            in2 => \_gnd_net_\,
            in3 => \N__31983\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47678\,
            ce => \N__32648\,
            sr => \N__46813\
        );

    \phase_controller_inst2.stoper_hc.target_time_9_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28160\,
            in1 => \N__31980\,
            in2 => \_gnd_net_\,
            in3 => \N__27023\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47669\,
            ce => \N__31314\,
            sr => \N__46822\
        );

    \phase_controller_inst2.stoper_hc.target_time_18_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__31975\,
            in1 => \N__28505\,
            in2 => \_gnd_net_\,
            in3 => \N__27005\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47669\,
            ce => \N__31314\,
            sr => \N__46822\
        );

    \phase_controller_inst2.stoper_hc.target_time_1_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__26984\,
            in1 => \N__31979\,
            in2 => \_gnd_net_\,
            in3 => \N__26959\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47669\,
            ce => \N__31314\,
            sr => \N__46822\
        );

    \phase_controller_inst2.stoper_hc.target_time_24_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31976\,
            in1 => \N__26921\,
            in2 => \_gnd_net_\,
            in3 => \N__29074\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47669\,
            ce => \N__31314\,
            sr => \N__46822\
        );

    \phase_controller_inst2.stoper_hc.target_time_17_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__26896\,
            in1 => \N__31982\,
            in2 => \_gnd_net_\,
            in3 => \N__28570\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47669\,
            ce => \N__31314\,
            sr => \N__46822\
        );

    \phase_controller_inst2.stoper_hc.target_time_6_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__31978\,
            in1 => \N__27554\,
            in2 => \_gnd_net_\,
            in3 => \N__26879\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47669\,
            ce => \N__31314\,
            sr => \N__46822\
        );

    \phase_controller_inst2.stoper_hc.target_time_14_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26852\,
            in1 => \N__27911\,
            in2 => \_gnd_net_\,
            in3 => \N__31981\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47669\,
            ce => \N__31314\,
            sr => \N__46822\
        );

    \phase_controller_inst2.stoper_hc.target_time_25_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31977\,
            in1 => \N__27209\,
            in2 => \_gnd_net_\,
            in3 => \N__29009\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47669\,
            ce => \N__31314\,
            sr => \N__46822\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27176\,
            in2 => \N__27185\,
            in3 => \N__29838\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_10_7_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29821\,
            in1 => \N__27170\,
            in2 => \N__27164\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27155\,
            in2 => \N__27149\,
            in3 => \N__30082\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27140\,
            in2 => \N__27131\,
            in3 => \N__30067\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27119\,
            in2 => \N__27113\,
            in3 => \N__30052\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27104\,
            in2 => \N__27098\,
            in3 => \N__30037\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30022\,
            in1 => \N__31328\,
            in2 => \N__27089\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30007\,
            in1 => \N__27314\,
            in2 => \N__29372\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_7\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27308\,
            in2 => \N__27299\,
            in3 => \N__29993\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_10_8_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29974\,
            in1 => \N__27290\,
            in2 => \N__27284\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27266\,
            in2 => \N__27275\,
            in3 => \N__30244\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27425\,
            in2 => \N__27260\,
            in3 => \N__30229\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30214\,
            in1 => \N__30482\,
            in2 => \N__27251\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27239\,
            in2 => \N__27230\,
            in3 => \N__30199\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29573\,
            in2 => \N__27218\,
            in3 => \N__30184\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29633\,
            in2 => \N__29669\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_15\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27359\,
            in2 => \N__27350\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_9_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31520\,
            in2 => \N__31475\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27335\,
            in2 => \N__27329\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_20\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27455\,
            in2 => \N__27491\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_22\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27416\,
            in2 => \N__27410\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_24\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27368\,
            in2 => \N__27842\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_26\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29870\,
            in2 => \N__29945\,
            in3 => \N__27317\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_28\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27494\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__30334\,
            in1 => \N__27482\,
            in2 => \N__27470\,
            in3 => \N__30315\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011001111"
        )
    port map (
            in0 => \N__27481\,
            in1 => \N__27469\,
            in2 => \N__30317\,
            in3 => \N__30333\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_12_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27449\,
            in1 => \N__27982\,
            in2 => \_gnd_net_\,
            in3 => \N__31905\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47622\,
            ce => \N__31310\,
            sr => \N__46849\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111010101111"
        )
    port map (
            in0 => \N__27379\,
            in1 => \N__30497\,
            in2 => \N__30274\,
            in3 => \N__30295\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010001110"
        )
    port map (
            in0 => \N__30493\,
            in1 => \N__27380\,
            in2 => \N__30275\,
            in3 => \N__30294\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_27_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28901\,
            in1 => \N__31774\,
            in2 => \_gnd_net_\,
            in3 => \N__27398\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47612\,
            ce => \N__31308\,
            sr => \N__46855\
        );

    \phase_controller_inst2.stoper_hc.target_time_28_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__31772\,
            in1 => \N__31132\,
            in2 => \_gnd_net_\,
            in3 => \N__31096\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47612\,
            ce => \N__31308\,
            sr => \N__46855\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__27850\,
            in1 => \N__30571\,
            in2 => \N__30596\,
            in3 => \N__27826\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__30591\,
            in1 => \N__30570\,
            in2 => \N__27830\,
            in3 => \N__27851\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_29_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31023\,
            in1 => \N__31775\,
            in2 => \_gnd_net_\,
            in3 => \N__31046\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47612\,
            ce => \N__31308\,
            sr => \N__46855\
        );

    \phase_controller_inst2.stoper_hc.target_time_31_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__31773\,
            in1 => \N__28717\,
            in2 => \_gnd_net_\,
            in3 => \N__27818\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47612\,
            ce => \N__31308\,
            sr => \N__46855\
        );

    \phase_controller_inst2.stoper_hc.target_time_30_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28759\,
            in1 => \N__27790\,
            in2 => \_gnd_net_\,
            in3 => \N__31776\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47612\,
            ce => \N__31308\,
            sr => \N__46855\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27773\,
            in2 => \N__27632\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\,
            ltout => OPEN,
            carryin => \bfn_10_12_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__47601\,
            ce => \N__28684\,
            sr => \N__46861\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27571\,
            in2 => \N__27710\,
            in3 => \N__27635\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__47601\,
            ce => \N__28684\,
            sr => \N__46861\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27631\,
            in2 => \N__27520\,
            in3 => \N__27575\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__47601\,
            ce => \N__28684\,
            sr => \N__46861\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27572\,
            in2 => \N__28213\,
            in3 => \N__27524\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__47601\,
            ce => \N__28684\,
            sr => \N__46861\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28183\,
            in2 => \N__27521\,
            in3 => \N__27497\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__47601\,
            ce => \N__28684\,
            sr => \N__46861\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28132\,
            in2 => \N__28214\,
            in3 => \N__28190\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__47601\,
            ce => \N__28684\,
            sr => \N__46861\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28078\,
            in2 => \N__28187\,
            in3 => \N__28136\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__47601\,
            ce => \N__28684\,
            sr => \N__46861\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28133\,
            in2 => \N__28018\,
            in3 => \N__28085\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__47601\,
            ce => \N__28684\,
            sr => \N__46861\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27952\,
            in2 => \N__28082\,
            in3 => \N__28022\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\,
            ltout => OPEN,
            carryin => \bfn_10_13_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__47593\,
            ce => \N__28685\,
            sr => \N__46866\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27931\,
            in2 => \N__28019\,
            in3 => \N__27956\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__47593\,
            ce => \N__28685\,
            sr => \N__46866\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27953\,
            in2 => \N__27877\,
            in3 => \N__27935\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__47593\,
            ce => \N__28685\,
            sr => \N__46866\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27932\,
            in2 => \N__28624\,
            in3 => \N__27881\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__47593\,
            ce => \N__28685\,
            sr => \N__46866\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28594\,
            in2 => \N__27878\,
            in3 => \N__27854\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__47593\,
            ce => \N__28685\,
            sr => \N__46866\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28528\,
            in2 => \N__28625\,
            in3 => \N__28601\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__47593\,
            ce => \N__28685\,
            sr => \N__46866\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28465\,
            in2 => \N__28598\,
            in3 => \N__28535\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__47593\,
            ce => \N__28685\,
            sr => \N__46866\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28384\,
            in2 => \N__28532\,
            in3 => \N__28472\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__47593\,
            ce => \N__28685\,
            sr => \N__46866\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28351\,
            in2 => \N__28469\,
            in3 => \N__28388\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\,
            ltout => OPEN,
            carryin => \bfn_10_14_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__47586\,
            ce => \N__28676\,
            sr => \N__46870\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28385\,
            in2 => \N__28330\,
            in3 => \N__28355\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__47586\,
            ce => \N__28676\,
            sr => \N__46870\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28352\,
            in2 => \N__28273\,
            in3 => \N__28334\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__47586\,
            ce => \N__28676\,
            sr => \N__46870\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29095\,
            in2 => \N__28331\,
            in3 => \N__28277\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__47586\,
            ce => \N__28676\,
            sr => \N__46870\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29032\,
            in2 => \N__28274\,
            in3 => \N__28217\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__47586\,
            ce => \N__28676\,
            sr => \N__46870\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28963\,
            in2 => \N__29099\,
            in3 => \N__29039\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__47586\,
            ce => \N__28676\,
            sr => \N__46870\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28933\,
            in2 => \N__29036\,
            in3 => \N__28970\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__47586\,
            ce => \N__28676\,
            sr => \N__46870\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28871\,
            in2 => \N__28967\,
            in3 => \N__28940\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__47586\,
            ce => \N__28676\,
            sr => \N__46870\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28840\,
            in2 => \N__28937\,
            in3 => \N__28874\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\,
            ltout => OPEN,
            carryin => \bfn_10_15_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__47580\,
            ce => \N__28675\,
            sr => \N__46874\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28870\,
            in2 => \N__28783\,
            in3 => \N__28844\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__47580\,
            ce => \N__28675\,
            sr => \N__46874\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28841\,
            in2 => \N__28823\,
            in3 => \N__28805\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__47580\,
            ce => \N__28675\,
            sr => \N__46874\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28802\,
            in2 => \N__28784\,
            in3 => \N__28724\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__47580\,
            ce => \N__28675\,
            sr => \N__46874\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28721\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47580\,
            ce => \N__28675\,
            sr => \N__46874\
        );

    \phase_controller_inst2.stoper_hc.target_time_8_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29432\,
            in1 => \N__29407\,
            in2 => \_gnd_net_\,
            in3 => \N__32003\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47577\,
            ce => \N__31307\,
            sr => \N__46880\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__30915\,
            in1 => \N__29279\,
            in2 => \_gnd_net_\,
            in3 => \N__32959\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_203_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D2_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29318\,
            lcout => \il_max_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47570\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__34331\,
            in1 => \N__32729\,
            in2 => \_gnd_net_\,
            in3 => \N__37589\,
            lcout => \current_shift_inst.control_input_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29278\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.start_timer_tr_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30719\,
            lcout => \delay_measurement_inst.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30677\,
            ce => 'H',
            sr => \N__46892\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37632\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.control_input_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37631\,
            lcout => \current_shift_inst.N_1304_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNISQD2_0_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29515\,
            in2 => \_gnd_net_\,
            in3 => \N__29556\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIBO26_1_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__29473\,
            in1 => \N__29494\,
            in2 => \N__29564\,
            in3 => \N__29536\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlt9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIFA6C_5_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__30602\,
            in1 => \N__29807\,
            in2 => \N__29561\,
            in3 => \N__29453\,
            lcout => \pwm_generator_inst.un1_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_0_LC_10_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29775\,
            in1 => \N__29558\,
            in2 => \_gnd_net_\,
            in3 => \N__29540\,
            lcout => \pwm_generator_inst.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_10_24_0_\,
            carryout => \pwm_generator_inst.counter_cry_0\,
            clk => \N__47555\,
            ce => 'H',
            sr => \N__46918\
        );

    \pwm_generator_inst.counter_1_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29771\,
            in1 => \N__29537\,
            in2 => \_gnd_net_\,
            in3 => \N__29519\,
            lcout => \pwm_generator_inst.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_0\,
            carryout => \pwm_generator_inst.counter_cry_1\,
            clk => \N__47555\,
            ce => 'H',
            sr => \N__46918\
        );

    \pwm_generator_inst.counter_2_LC_10_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29776\,
            in1 => \N__29516\,
            in2 => \_gnd_net_\,
            in3 => \N__29498\,
            lcout => \pwm_generator_inst.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_1\,
            carryout => \pwm_generator_inst.counter_cry_2\,
            clk => \N__47555\,
            ce => 'H',
            sr => \N__46918\
        );

    \pwm_generator_inst.counter_3_LC_10_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29772\,
            in1 => \N__29495\,
            in2 => \_gnd_net_\,
            in3 => \N__29477\,
            lcout => \pwm_generator_inst.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_2\,
            carryout => \pwm_generator_inst.counter_cry_3\,
            clk => \N__47555\,
            ce => 'H',
            sr => \N__46918\
        );

    \pwm_generator_inst.counter_4_LC_10_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29777\,
            in1 => \N__29474\,
            in2 => \_gnd_net_\,
            in3 => \N__29456\,
            lcout => \pwm_generator_inst.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_3\,
            carryout => \pwm_generator_inst.counter_cry_4\,
            clk => \N__47555\,
            ce => 'H',
            sr => \N__46918\
        );

    \pwm_generator_inst.counter_5_LC_10_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29773\,
            in1 => \N__29452\,
            in2 => \_gnd_net_\,
            in3 => \N__29435\,
            lcout => \pwm_generator_inst.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_4\,
            carryout => \pwm_generator_inst.counter_cry_5\,
            clk => \N__47555\,
            ce => 'H',
            sr => \N__46918\
        );

    \pwm_generator_inst.counter_6_LC_10_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29778\,
            in1 => \N__29806\,
            in2 => \_gnd_net_\,
            in3 => \N__29789\,
            lcout => \pwm_generator_inst.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_5\,
            carryout => \pwm_generator_inst.counter_cry_6\,
            clk => \N__47555\,
            ce => 'H',
            sr => \N__46918\
        );

    \pwm_generator_inst.counter_7_LC_10_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29774\,
            in1 => \N__30622\,
            in2 => \_gnd_net_\,
            in3 => \N__29786\,
            lcout => \pwm_generator_inst.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_6\,
            carryout => \pwm_generator_inst.counter_cry_7\,
            clk => \N__47555\,
            ce => 'H',
            sr => \N__46918\
        );

    \pwm_generator_inst.counter_8_LC_10_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29780\,
            in1 => \N__30643\,
            in2 => \_gnd_net_\,
            in3 => \N__29783\,
            lcout => \pwm_generator_inst.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_10_25_0_\,
            carryout => \pwm_generator_inst.counter_cry_8\,
            clk => \N__47552\,
            ce => 'H',
            sr => \N__46922\
        );

    \pwm_generator_inst.counter_9_LC_10_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__30664\,
            in1 => \N__29779\,
            in2 => \_gnd_net_\,
            in3 => \N__29738\,
            lcout => \pwm_generator_inst.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47552\,
            ce => 'H',
            sr => \N__46922\
        );

    \phase_controller_inst2.start_timer_hc_RNO_0_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__31203\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31173\,
            lcout => \phase_controller_inst2.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_16_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29735\,
            in1 => \N__29714\,
            in2 => \_gnd_net_\,
            in3 => \N__32005\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47670\,
            ce => \N__31316\,
            sr => \N__46804\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110101000100"
        )
    port map (
            in0 => \N__30139\,
            in1 => \N__29645\,
            in2 => \N__30170\,
            in3 => \N__29654\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__29653\,
            in1 => \N__30169\,
            in2 => \N__30143\,
            in3 => \N__29644\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_15_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29624\,
            in1 => \N__29588\,
            in2 => \_gnd_net_\,
            in3 => \N__32004\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47656\,
            ce => \N__31315\,
            sr => \N__46814\
        );

    \phase_controller_inst2.stoper_hc.target_time_RNISIH31_30_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__30550\,
            in1 => \N__30524\,
            in2 => \N__29924\,
            in3 => \N__29889\,
            lcout => OPEN,
            ltout => \phase_controller_inst2.stoper_hc.un4_running_df30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIEABO2_28_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100111011"
        )
    port map (
            in0 => \N__29935\,
            in1 => \N__32230\,
            in2 => \N__29960\,
            in3 => \N__29957\,
            lcout => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29948\,
            in3 => \N__32295\,
            lcout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_RNISIH31_0_30_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010001110"
        )
    port map (
            in0 => \N__29919\,
            in1 => \N__30519\,
            in2 => \N__29893\,
            in3 => \N__30549\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3_28_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32296\,
            in2 => \_gnd_net_\,
            in3 => \N__29860\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011001111"
        )
    port map (
            in0 => \N__29920\,
            in1 => \N__30520\,
            in2 => \N__29894\,
            in3 => \N__30551\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010001010000"
        )
    port map (
            in0 => \N__32172\,
            in1 => \N__29861\,
            in2 => \N__29846\,
            in3 => \N__32297\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47646\,
            ce => 'H',
            sr => \N__46823\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29852\,
            in2 => \N__29845\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_8_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32177\,
            in1 => \N__29822\,
            in2 => \_gnd_net_\,
            in3 => \N__29810\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \N__47634\,
            ce => 'H',
            sr => \N__46829\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__32181\,
            in1 => \N__30083\,
            in2 => \N__30092\,
            in3 => \N__30071\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \N__47634\,
            ce => 'H',
            sr => \N__46829\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32178\,
            in1 => \N__30068\,
            in2 => \_gnd_net_\,
            in3 => \N__30056\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \N__47634\,
            ce => 'H',
            sr => \N__46829\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32182\,
            in1 => \N__30053\,
            in2 => \_gnd_net_\,
            in3 => \N__30041\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \N__47634\,
            ce => 'H',
            sr => \N__46829\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32179\,
            in1 => \N__30038\,
            in2 => \_gnd_net_\,
            in3 => \N__30026\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \N__47634\,
            ce => 'H',
            sr => \N__46829\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32183\,
            in1 => \N__30023\,
            in2 => \_gnd_net_\,
            in3 => \N__30011\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \N__47634\,
            ce => 'H',
            sr => \N__46829\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32180\,
            in1 => \N__30008\,
            in2 => \_gnd_net_\,
            in3 => \N__29996\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \N__47634\,
            ce => 'H',
            sr => \N__46829\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32176\,
            in1 => \N__29992\,
            in2 => \_gnd_net_\,
            in3 => \N__29978\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \N__47623\,
            ce => 'H',
            sr => \N__46837\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32188\,
            in1 => \N__29975\,
            in2 => \_gnd_net_\,
            in3 => \N__29963\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \N__47623\,
            ce => 'H',
            sr => \N__46837\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32173\,
            in1 => \N__30245\,
            in2 => \_gnd_net_\,
            in3 => \N__30233\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \N__47623\,
            ce => 'H',
            sr => \N__46837\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32189\,
            in1 => \N__30230\,
            in2 => \_gnd_net_\,
            in3 => \N__30218\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \N__47623\,
            ce => 'H',
            sr => \N__46837\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32174\,
            in1 => \N__30215\,
            in2 => \_gnd_net_\,
            in3 => \N__30203\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \N__47623\,
            ce => 'H',
            sr => \N__46837\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32190\,
            in1 => \N__30200\,
            in2 => \_gnd_net_\,
            in3 => \N__30188\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \N__47623\,
            ce => 'H',
            sr => \N__46837\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32175\,
            in1 => \N__30185\,
            in2 => \_gnd_net_\,
            in3 => \N__30173\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \N__47623\,
            ce => 'H',
            sr => \N__46837\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32191\,
            in1 => \N__30160\,
            in2 => \_gnd_net_\,
            in3 => \N__30146\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \N__47623\,
            ce => 'H',
            sr => \N__46837\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32184\,
            in1 => \N__30138\,
            in2 => \_gnd_net_\,
            in3 => \N__30119\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_11_10_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \N__47613\,
            ce => 'H',
            sr => \N__46844\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32165\,
            in1 => \N__30109\,
            in2 => \_gnd_net_\,
            in3 => \N__30095\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \N__47613\,
            ce => 'H',
            sr => \N__46844\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32185\,
            in1 => \N__30409\,
            in2 => \_gnd_net_\,
            in3 => \N__30395\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \N__47613\,
            ce => 'H',
            sr => \N__46844\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32166\,
            in1 => \N__31510\,
            in2 => \_gnd_net_\,
            in3 => \N__30392\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \N__47613\,
            ce => 'H',
            sr => \N__46844\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32186\,
            in1 => \N__31492\,
            in2 => \_gnd_net_\,
            in3 => \N__30389\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\,
            clk => \N__47613\,
            ce => 'H',
            sr => \N__46844\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32167\,
            in1 => \N__30376\,
            in2 => \_gnd_net_\,
            in3 => \N__30362\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\,
            clk => \N__47613\,
            ce => 'H',
            sr => \N__46844\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32187\,
            in1 => \N__30352\,
            in2 => \_gnd_net_\,
            in3 => \N__30338\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\,
            clk => \N__47613\,
            ce => 'H',
            sr => \N__46844\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32168\,
            in1 => \N__30335\,
            in2 => \_gnd_net_\,
            in3 => \N__30320\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\,
            clk => \N__47613\,
            ce => 'H',
            sr => \N__46844\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32109\,
            in1 => \N__30316\,
            in2 => \_gnd_net_\,
            in3 => \N__30299\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_11_11_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\,
            clk => \N__47602\,
            ce => 'H',
            sr => \N__46850\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32113\,
            in1 => \N__30296\,
            in2 => \_gnd_net_\,
            in3 => \N__30278\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\,
            clk => \N__47602\,
            ce => 'H',
            sr => \N__46850\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32110\,
            in1 => \N__30270\,
            in2 => \_gnd_net_\,
            in3 => \N__30248\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\,
            clk => \N__47602\,
            ce => 'H',
            sr => \N__46850\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32114\,
            in1 => \N__30595\,
            in2 => \_gnd_net_\,
            in3 => \N__30575\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\,
            clk => \N__47602\,
            ce => 'H',
            sr => \N__46850\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32111\,
            in1 => \N__30572\,
            in2 => \_gnd_net_\,
            in3 => \N__30554\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\,
            clk => \N__47602\,
            ce => 'H',
            sr => \N__46850\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32115\,
            in1 => \N__30548\,
            in2 => \_gnd_net_\,
            in3 => \N__30530\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\,
            clk => \N__47602\,
            ce => 'H',
            sr => \N__46850\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32112\,
            in1 => \N__30518\,
            in2 => \_gnd_net_\,
            in3 => \N__30527\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47602\,
            ce => 'H',
            sr => \N__46850\
        );

    \phase_controller_inst2.stoper_hc.target_time_26_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31833\,
            in1 => \N__30745\,
            in2 => \_gnd_net_\,
            in3 => \N__30775\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47594\,
            ce => \N__31309\,
            sr => \N__46856\
        );

    \phase_controller_inst2.stoper_hc.target_time_13_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30435\,
            in1 => \N__30466\,
            in2 => \_gnd_net_\,
            in3 => \N__31834\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47594\,
            ce => \N__31309\,
            sr => \N__46856\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30439\,
            in1 => \N__30465\,
            in2 => \_gnd_net_\,
            in3 => \N__31943\,
            lcout => \elapsed_time_ns_1_RNI02CN9_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44192\,
            in1 => \N__39281\,
            in2 => \N__45051\,
            in3 => \N__42190\,
            lcout => \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__42799\,
            in1 => \N__45003\,
            in2 => \N__39374\,
            in3 => \N__44193\,
            lcout => \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_ns_i_a2_1_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__30810\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34662\,
            lcout => state_ns_i_a2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33444\,
            in2 => \N__30725\,
            in3 => \N__30694\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_205_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30768\,
            in1 => \N__30744\,
            in2 => \_gnd_net_\,
            in3 => \N__31937\,
            lcout => \elapsed_time_ns_1_RNI47DN9_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33443\,
            in2 => \_gnd_net_\,
            in3 => \N__30693\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_204_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__33445\,
            in1 => \N__30724\,
            in2 => \_gnd_net_\,
            in3 => \N__30695\,
            lcout => \delay_measurement_inst.delay_tr_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47571\,
            ce => 'H',
            sr => \N__46875\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \N__45035\,
            in1 => \N__40022\,
            in2 => \N__44416\,
            in3 => \N__43441\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__44355\,
            in1 => \N__40072\,
            in2 => \N__43309\,
            in3 => \N__45036\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_tr_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30720\,
            lcout => \delay_measurement_inst.stop_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30676\,
            ce => 'H',
            sr => \N__46887\
        );

    \pwm_generator_inst.counter_RNIVDL3_9_LC_11_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__30665\,
            in1 => \N__30644\,
            in2 => \_gnd_net_\,
            in3 => \N__30618\,
            lcout => \pwm_generator_inst.un1_counterlto9_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_hc_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32947\,
            lcout => \delay_measurement_inst.stop_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32926\,
            ce => 'H',
            sr => \N__46914\
        );

    \GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_11_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30887\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_clk_12mhz_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_RNIG7JF_2_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__30862\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31275\,
            lcout => \phase_controller_inst2.state_RNIG7JFZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_tr_RNO_0_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__30861\,
            in1 => \N__31276\,
            in2 => \N__33010\,
            in3 => \N__31238\,
            lcout => \phase_controller_inst2.start_timer_tr_RNO_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_tr_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010111010"
        )
    port map (
            in0 => \N__30869\,
            in1 => \N__32891\,
            in2 => \N__32878\,
            in3 => \N__34689\,
            lcout => \phase_controller_inst2.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47668\,
            ce => 'H',
            sr => \N__46792\
        );

    \phase_controller_inst2.state_2_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000111110001000"
        )
    port map (
            in0 => \N__31204\,
            in1 => \N__31169\,
            in2 => \N__31280\,
            in3 => \N__30863\,
            lcout => \phase_controller_inst2.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47668\,
            ce => 'H',
            sr => \N__46792\
        );

    \phase_controller_inst2.start_timer_hc_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__34688\,
            in1 => \N__30838\,
            in2 => \N__32261\,
            in3 => \N__30848\,
            lcout => \phase_controller_inst2.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47668\,
            ce => 'H',
            sr => \N__46792\
        );

    \phase_controller_inst2.state_1_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__31237\,
            in1 => \N__33003\,
            in2 => \_gnd_net_\,
            in3 => \N__30842\,
            lcout => \phase_controller_inst2.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47655\,
            ce => 'H',
            sr => \N__46797\
        );

    \phase_controller_inst2.stoper_tr.start_latched_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32879\,
            lcout => \phase_controller_inst2.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47655\,
            ce => 'H',
            sr => \N__46797\
        );

    \phase_controller_inst2.state_0_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000111110001000"
        )
    port map (
            in0 => \N__31236\,
            in1 => \N__33002\,
            in2 => \N__32852\,
            in3 => \N__32903\,
            lcout => \phase_controller_inst2.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47655\,
            ce => 'H',
            sr => \N__46797\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__33077\,
            in1 => \N__33050\,
            in2 => \N__34728\,
            in3 => \N__34092\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47645\,
            ce => 'H',
            sr => \N__46805\
        );

    \phase_controller_inst2.state_3_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111011100"
        )
    port map (
            in0 => \N__31208\,
            in1 => \N__32890\,
            in2 => \N__31174\,
            in3 => \N__33791\,
            lcout => \phase_controller_inst2.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47645\,
            ce => 'H',
            sr => \N__46805\
        );

    \phase_controller_inst1.stoper_hc.target_time_28_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31133\,
            in1 => \N__31097\,
            in2 => \_gnd_net_\,
            in3 => \N__32006\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47633\,
            ce => \N__32656\,
            sr => \N__46815\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100000010"
        )
    port map (
            in0 => \N__30992\,
            in1 => \N__30982\,
            in2 => \N__30964\,
            in3 => \N__30941\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31024\,
            in1 => \N__31984\,
            in2 => \_gnd_net_\,
            in3 => \N__31039\,
            lcout => \elapsed_time_ns_1_RNI7ADN9_0_29\,
            ltout => \elapsed_time_ns_1_RNI7ADN9_0_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_29_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__31986\,
            in1 => \_gnd_net_\,
            in2 => \N__31028\,
            in3 => \N__31025\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47621\,
            ce => \N__32594\,
            sr => \N__46824\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__30991\,
            in1 => \N__30983\,
            in2 => \N__30965\,
            in3 => \N__30940\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__31985\,
            in1 => \N__31371\,
            in2 => \_gnd_net_\,
            in3 => \N__31339\,
            lcout => \elapsed_time_ns_1_RNIJ53T9_0_7\,
            ltout => \elapsed_time_ns_1_RNIJ53T9_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__31372\,
            in1 => \_gnd_net_\,
            in2 => \N__31535\,
            in3 => \N__31987\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47621\,
            ce => \N__32594\,
            sr => \N__46824\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101110"
        )
    port map (
            in0 => \N__31382\,
            in1 => \N__31463\,
            in2 => \N__31511\,
            in3 => \N__31491\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__31462\,
            in1 => \N__31509\,
            in2 => \N__31493\,
            in3 => \N__31381\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_20_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32045\,
            in1 => \N__31561\,
            in2 => \_gnd_net_\,
            in3 => \N__31958\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47611\,
            ce => \N__31313\,
            sr => \N__46830\
        );

    \phase_controller_inst2.stoper_hc.target_time_21_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31956\,
            in1 => \N__31454\,
            in2 => \_gnd_net_\,
            in3 => \N__31424\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47611\,
            ce => \N__31313\,
            sr => \N__46830\
        );

    \phase_controller_inst2.stoper_hc.target_time_7_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__31957\,
            in1 => \N__31373\,
            in2 => \_gnd_net_\,
            in3 => \N__31340\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47611\,
            ce => \N__31313\,
            sr => \N__46830\
        );

    \phase_controller_inst2.stoper_hc.time_passed_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110000001100"
        )
    port map (
            in0 => \N__31252\,
            in1 => \N__31274\,
            in2 => \N__32294\,
            in3 => \N__32229\,
            lcout => \phase_controller_inst2.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47600\,
            ce => 'H',
            sr => \N__46838\
        );

    \phase_controller_inst2.stoper_hc.start_latched_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32266\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47600\,
            ce => 'H',
            sr => \N__46838\
        );

    \phase_controller_inst2.stoper_hc.running_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111110000"
        )
    port map (
            in0 => \N__32228\,
            in1 => \N__31253\,
            in2 => \N__32312\,
            in3 => \N__32286\,
            lcout => \phase_controller_inst2.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47600\,
            ce => 'H',
            sr => \N__46838\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__42040\,
            in1 => \N__42062\,
            in2 => \N__38674\,
            in3 => \N__47191\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47592\,
            ce => 'H',
            sr => \N__46845\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__32497\,
            in1 => \N__32399\,
            in2 => \N__32384\,
            in3 => \N__32328\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47592\,
            ce => 'H',
            sr => \N__46845\
        );

    \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__32221\,
            in1 => \N__32308\,
            in2 => \_gnd_net_\,
            in3 => \N__32262\,
            lcout => \phase_controller_inst2.stoper_hc.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__32267\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32231\,
            lcout => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31560\,
            in1 => \N__32041\,
            in2 => \_gnd_net_\,
            in3 => \N__31938\,
            lcout => \elapsed_time_ns_1_RNIU0DN9_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42261\,
            lcout => \current_shift_inst.un4_control_input1_1\,
            ltout => \current_shift_inst.un4_control_input1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44191\,
            in2 => \N__31538\,
            in3 => \N__33199\,
            lcout => \current_shift_inst.un38_control_input_cry_0_s0_sf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42416\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47576\,
            ce => \N__43572\,
            sr => \N__46862\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__44189\,
            in1 => \N__44919\,
            in2 => \N__39326\,
            in3 => \N__42226\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__42227\,
            in1 => \N__39325\,
            in2 => \N__45029\,
            in3 => \N__44190\,
            lcout => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34262\,
            in2 => \N__33464\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_15_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45157\,
            in2 => \N__45131\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44858\,
            in2 => \N__32693\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32684\,
            in2 => \N__45004\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44862\,
            in2 => \N__36359\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36098\,
            in2 => \N__45005\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s1_c_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44866\,
            in2 => \N__39770\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s1_c_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32678\,
            in2 => \N__45006\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s1_c_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44870\,
            in2 => \N__36068\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_16_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s1_c_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33275\,
            in2 => \N__45007\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s1_c_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44874\,
            in2 => \N__33290\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s1_c_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33296\,
            in2 => \N__45008\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s1_c_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44878\,
            in2 => \N__33269\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s1_c_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33545\,
            in2 => \N__45009\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s1_c_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44882\,
            in2 => \N__33539\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s1_c_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33281\,
            in2 => \N__45010\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s1_c_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44886\,
            in2 => \N__33515\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_17_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s1_c_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40205\,
            in2 => \N__45011\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s1_c_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44890\,
            in2 => \N__33530\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33521\,
            in2 => \N__45012\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44894\,
            in2 => \N__33506\,
            in3 => \N__32720\,
            lcout => \current_shift_inst.un38_control_input_0_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40214\,
            in2 => \N__45013\,
            in3 => \N__32717\,
            lcout => \current_shift_inst.un38_control_input_0_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44898\,
            in2 => \N__32714\,
            in3 => \N__32702\,
            lcout => \current_shift_inst.un38_control_input_0_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33497\,
            in2 => \N__45014\,
            in3 => \N__32699\,
            lcout => \current_shift_inst.un38_control_input_0_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45015\,
            in2 => \N__33803\,
            in3 => \N__32696\,
            lcout => \current_shift_inst.un38_control_input_0_s1_24\,
            ltout => OPEN,
            carryin => \bfn_12_18_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32783\,
            in2 => \N__45052\,
            in3 => \N__32777\,
            lcout => \current_shift_inst.un38_control_input_0_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45019\,
            in2 => \N__34439\,
            in3 => \N__32774\,
            lcout => \current_shift_inst.un38_control_input_0_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36470\,
            in2 => \N__45053\,
            in3 => \N__32771\,
            lcout => \current_shift_inst.un38_control_input_0_s1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45023\,
            in2 => \N__40232\,
            in3 => \N__32768\,
            lcout => \current_shift_inst.un38_control_input_0_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33677\,
            in2 => \N__45054\,
            in3 => \N__32765\,
            lcout => \current_shift_inst.un38_control_input_0_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45027\,
            in2 => \N__45113\,
            in3 => \N__32762\,
            lcout => \current_shift_inst.un38_control_input_0_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__45028\,
            in1 => \N__44391\,
            in2 => \_gnd_net_\,
            in3 => \N__32759\,
            lcout => \current_shift_inst.un38_control_input_0_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D2_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32735\,
            lcout => \il_min_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47560\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D1_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32756\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_min_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47560\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.S2_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33011\,
            lcout => s4_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47557\,
            ce => 'H',
            sr => \N__46896\
        );

    \delay_measurement_inst.start_timer_hc_LC_12_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32946\,
            lcout => \delay_measurement_inst.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32927\,
            ce => 'H',
            sr => \N__46909\
        );

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46958\,
            lcout => \pll_inst.red_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_RNI9M3O_0_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32847\,
            in2 => \_gnd_net_\,
            in3 => \N__32902\,
            lcout => \phase_controller_inst2.state_RNI9M3OZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_13_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__32801\,
            in1 => \N__32830\,
            in2 => \_gnd_net_\,
            in3 => \N__32870\,
            lcout => \phase_controller_inst2.stoper_tr.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_13_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__32871\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32802\,
            lcout => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.time_passed_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101000011001100"
        )
    port map (
            in0 => \N__35296\,
            in1 => \N__32851\,
            in2 => \N__32813\,
            in3 => \N__33076\,
            lcout => \phase_controller_inst2.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47657\,
            ce => 'H',
            sr => \N__46798\
        );

    \phase_controller_inst2.stoper_tr.running_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111110000"
        )
    port map (
            in0 => \N__32812\,
            in1 => \N__35297\,
            in2 => \N__32831\,
            in3 => \N__33079\,
            lcout => \phase_controller_inst2.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47647\,
            ce => 'H',
            sr => \N__46806\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNISIOB3_28_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100111011"
        )
    port map (
            in0 => \N__35332\,
            in1 => \N__32811\,
            in2 => \N__33038\,
            in3 => \N__35315\,
            lcout => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33083\,
            in3 => \N__33078\,
            lcout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41524\,
            in1 => \N__41503\,
            in2 => \_gnd_net_\,
            in3 => \N__48116\,
            lcout => \elapsed_time_ns_1_RNI1BOBB_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34_28_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33080\,
            in2 => \_gnd_net_\,
            in3 => \N__33049\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48117\,
            in1 => \N__37216\,
            in2 => \_gnd_net_\,
            in3 => \N__37260\,
            lcout => \elapsed_time_ns_1_RNIGF91B_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_0_30_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001100"
        )
    port map (
            in0 => \N__34206\,
            in1 => \N__34023\,
            in2 => \N__33119\,
            in3 => \N__33025\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_30_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__33024\,
            in1 => \N__34207\,
            in2 => \N__34030\,
            in3 => \N__33114\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_df30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_30_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__41063\,
            in1 => \N__48187\,
            in2 => \_gnd_net_\,
            in3 => \N__34001\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47624\,
            ce => \N__45954\,
            sr => \N__46825\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011111011"
        )
    port map (
            in0 => \N__33026\,
            in1 => \N__34208\,
            in2 => \N__34031\,
            in3 => \N__33118\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__34273\,
            in1 => \N__48186\,
            in2 => \_gnd_net_\,
            in3 => \N__38457\,
            lcout => \elapsed_time_ns_1_RNI0AOBB_0_13\,
            ltout => \elapsed_time_ns_1_RNI0AOBB_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_13_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__48189\,
            in1 => \_gnd_net_\,
            in2 => \N__33014\,
            in3 => \N__38458\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47624\,
            ce => \N__45954\,
            sr => \N__46825\
        );

    \phase_controller_inst2.stoper_tr.target_time_31_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__34295\,
            in1 => \N__48188\,
            in2 => \_gnd_net_\,
            in3 => \N__38356\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47624\,
            ce => \N__45954\,
            sr => \N__46825\
        );

    \phase_controller_inst2.stoper_tr.target_time_14_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__41504\,
            in1 => \N__41520\,
            in2 => \N__48206\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47624\,
            ce => \N__45954\,
            sr => \N__46825\
        );

    \delay_measurement_inst.delay_tr_timer.counter_0_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33405\,
            in1 => \N__35604\,
            in2 => \_gnd_net_\,
            in3 => \N__33104\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_13_10_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            clk => \N__47614\,
            ce => \N__33245\,
            sr => \N__46831\
        );

    \delay_measurement_inst.delay_tr_timer.counter_1_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33397\,
            in1 => \N__35577\,
            in2 => \_gnd_net_\,
            in3 => \N__33101\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            clk => \N__47614\,
            ce => \N__33245\,
            sr => \N__46831\
        );

    \delay_measurement_inst.delay_tr_timer.counter_2_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33406\,
            in1 => \N__35547\,
            in2 => \_gnd_net_\,
            in3 => \N__33098\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            clk => \N__47614\,
            ce => \N__33245\,
            sr => \N__46831\
        );

    \delay_measurement_inst.delay_tr_timer.counter_3_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33398\,
            in1 => \N__35526\,
            in2 => \_gnd_net_\,
            in3 => \N__33095\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            clk => \N__47614\,
            ce => \N__33245\,
            sr => \N__46831\
        );

    \delay_measurement_inst.delay_tr_timer.counter_4_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33407\,
            in1 => \N__35502\,
            in2 => \_gnd_net_\,
            in3 => \N__33092\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            clk => \N__47614\,
            ce => \N__33245\,
            sr => \N__46831\
        );

    \delay_measurement_inst.delay_tr_timer.counter_5_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33399\,
            in1 => \N__35472\,
            in2 => \_gnd_net_\,
            in3 => \N__33089\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            clk => \N__47614\,
            ce => \N__33245\,
            sr => \N__46831\
        );

    \delay_measurement_inst.delay_tr_timer.counter_6_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33408\,
            in1 => \N__35453\,
            in2 => \_gnd_net_\,
            in3 => \N__33086\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            clk => \N__47614\,
            ce => \N__33245\,
            sr => \N__46831\
        );

    \delay_measurement_inst.delay_tr_timer.counter_7_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33400\,
            in1 => \N__35427\,
            in2 => \_gnd_net_\,
            in3 => \N__33146\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            clk => \N__47614\,
            ce => \N__33245\,
            sr => \N__46831\
        );

    \delay_measurement_inst.delay_tr_timer.counter_8_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33396\,
            in1 => \N__35394\,
            in2 => \_gnd_net_\,
            in3 => \N__33143\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_13_11_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            clk => \N__47603\,
            ce => \N__33244\,
            sr => \N__46839\
        );

    \delay_measurement_inst.delay_tr_timer.counter_9_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33404\,
            in1 => \N__35823\,
            in2 => \_gnd_net_\,
            in3 => \N__33140\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            clk => \N__47603\,
            ce => \N__33244\,
            sr => \N__46839\
        );

    \delay_measurement_inst.delay_tr_timer.counter_10_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33393\,
            in1 => \N__35793\,
            in2 => \_gnd_net_\,
            in3 => \N__33137\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            clk => \N__47603\,
            ce => \N__33244\,
            sr => \N__46839\
        );

    \delay_measurement_inst.delay_tr_timer.counter_11_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33401\,
            in1 => \N__35769\,
            in2 => \_gnd_net_\,
            in3 => \N__33134\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            clk => \N__47603\,
            ce => \N__33244\,
            sr => \N__46839\
        );

    \delay_measurement_inst.delay_tr_timer.counter_12_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33394\,
            in1 => \N__35739\,
            in2 => \_gnd_net_\,
            in3 => \N__33131\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            clk => \N__47603\,
            ce => \N__33244\,
            sr => \N__46839\
        );

    \delay_measurement_inst.delay_tr_timer.counter_13_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33402\,
            in1 => \N__35715\,
            in2 => \_gnd_net_\,
            in3 => \N__33128\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            clk => \N__47603\,
            ce => \N__33244\,
            sr => \N__46839\
        );

    \delay_measurement_inst.delay_tr_timer.counter_14_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33395\,
            in1 => \N__35688\,
            in2 => \_gnd_net_\,
            in3 => \N__33125\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            clk => \N__47603\,
            ce => \N__33244\,
            sr => \N__46839\
        );

    \delay_measurement_inst.delay_tr_timer.counter_15_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33403\,
            in1 => \N__35666\,
            in2 => \_gnd_net_\,
            in3 => \N__33122\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            clk => \N__47603\,
            ce => \N__33244\,
            sr => \N__46839\
        );

    \delay_measurement_inst.delay_tr_timer.counter_16_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33415\,
            in1 => \N__35637\,
            in2 => \_gnd_net_\,
            in3 => \N__33173\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_13_12_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            clk => \N__47595\,
            ce => \N__33237\,
            sr => \N__46846\
        );

    \delay_measurement_inst.delay_tr_timer.counter_17_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33419\,
            in1 => \N__36030\,
            in2 => \_gnd_net_\,
            in3 => \N__33170\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            clk => \N__47595\,
            ce => \N__33237\,
            sr => \N__46846\
        );

    \delay_measurement_inst.delay_tr_timer.counter_18_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33416\,
            in1 => \N__36001\,
            in2 => \_gnd_net_\,
            in3 => \N__33167\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            clk => \N__47595\,
            ce => \N__33237\,
            sr => \N__46846\
        );

    \delay_measurement_inst.delay_tr_timer.counter_19_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33420\,
            in1 => \N__35976\,
            in2 => \_gnd_net_\,
            in3 => \N__33164\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            clk => \N__47595\,
            ce => \N__33237\,
            sr => \N__46846\
        );

    \delay_measurement_inst.delay_tr_timer.counter_20_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33417\,
            in1 => \N__35955\,
            in2 => \_gnd_net_\,
            in3 => \N__33161\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            clk => \N__47595\,
            ce => \N__33237\,
            sr => \N__46846\
        );

    \delay_measurement_inst.delay_tr_timer.counter_21_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33421\,
            in1 => \N__35931\,
            in2 => \_gnd_net_\,
            in3 => \N__33158\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            clk => \N__47595\,
            ce => \N__33237\,
            sr => \N__46846\
        );

    \delay_measurement_inst.delay_tr_timer.counter_22_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33418\,
            in1 => \N__35901\,
            in2 => \_gnd_net_\,
            in3 => \N__33155\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            clk => \N__47595\,
            ce => \N__33237\,
            sr => \N__46846\
        );

    \delay_measurement_inst.delay_tr_timer.counter_23_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33422\,
            in1 => \N__35874\,
            in2 => \_gnd_net_\,
            in3 => \N__33152\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            clk => \N__47595\,
            ce => \N__33237\,
            sr => \N__46846\
        );

    \delay_measurement_inst.delay_tr_timer.counter_24_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33409\,
            in1 => \N__35844\,
            in2 => \_gnd_net_\,
            in3 => \N__33149\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_13_13_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            clk => \N__47587\,
            ce => \N__33236\,
            sr => \N__46851\
        );

    \delay_measurement_inst.delay_tr_timer.counter_25_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33413\,
            in1 => \N__36279\,
            in2 => \_gnd_net_\,
            in3 => \N__33260\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            clk => \N__47587\,
            ce => \N__33236\,
            sr => \N__46851\
        );

    \delay_measurement_inst.delay_tr_timer.counter_26_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33410\,
            in1 => \N__36235\,
            in2 => \_gnd_net_\,
            in3 => \N__33257\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            clk => \N__47587\,
            ce => \N__33236\,
            sr => \N__46851\
        );

    \delay_measurement_inst.delay_tr_timer.counter_27_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33414\,
            in1 => \N__36192\,
            in2 => \_gnd_net_\,
            in3 => \N__33254\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            clk => \N__47587\,
            ce => \N__33236\,
            sr => \N__46851\
        );

    \delay_measurement_inst.delay_tr_timer.counter_28_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33411\,
            in1 => \N__36253\,
            in2 => \_gnd_net_\,
            in3 => \N__33251\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_28\,
            clk => \N__47587\,
            ce => \N__33236\,
            sr => \N__46851\
        );

    \delay_measurement_inst.delay_tr_timer.counter_29_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__36211\,
            in1 => \N__33412\,
            in2 => \_gnd_net_\,
            in3 => \N__33248\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47587\,
            ce => \N__33236\,
            sr => \N__46851\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40154\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47581\,
            ce => \N__43571\,
            sr => \N__46857\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33194\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_1\,
            ltout => \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__33195\,
            in1 => \_gnd_net_\,
            in2 => \N__33203\,
            in3 => \N__42383\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42415\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_fast_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47581\,
            ce => \N__43571\,
            sr => \N__46857\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44239\,
            in2 => \N__33200\,
            in3 => \N__33179\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_0_c_inv_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__37501\,
            in1 => \N__37759\,
            in2 => \_gnd_net_\,
            in3 => \N__33473\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_31\,
            ltout => \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \N__37760\,
            in1 => \_gnd_net_\,
            in2 => \N__33467\,
            in3 => \N__33463\,
            lcout => \current_shift_inst.un38_control_input_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__44925\,
            in1 => \N__44200\,
            in2 => \N__39710\,
            in3 => \N__43183\,
            lcout => \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33449\,
            lcout => \delay_measurement_inst.delay_tr_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__44924\,
            in1 => \N__44196\,
            in2 => \N__39620\,
            in3 => \N__42631\,
            lcout => \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__44195\,
            in1 => \N__44923\,
            in2 => \N__42671\,
            in3 => \N__39664\,
            lcout => \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__43070\,
            in1 => \N__44199\,
            in2 => \N__45030\,
            in3 => \N__39571\,
            lcout => \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__44194\,
            in1 => \N__39493\,
            in2 => \N__42719\,
            in3 => \N__44931\,
            lcout => \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__44926\,
            in1 => \N__44197\,
            in2 => \N__39709\,
            in3 => \N__43184\,
            lcout => \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__44198\,
            in1 => \N__44927\,
            in2 => \N__39757\,
            in3 => \N__43147\,
            lcout => \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__44291\,
            in1 => \N__44935\,
            in2 => \N__43121\,
            in3 => \N__44061\,
            lcout => \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110011"
        )
    port map (
            in0 => \N__44932\,
            in1 => \N__40018\,
            in2 => \N__43442\,
            in3 => \N__44297\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110110001101"
        )
    port map (
            in0 => \N__44293\,
            in1 => \N__42956\,
            in2 => \N__39925\,
            in3 => \N__44937\,
            lcout => \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__44938\,
            in1 => \N__44294\,
            in2 => \N__43907\,
            in3 => \N__42931\,
            lcout => \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__44292\,
            in1 => \N__44936\,
            in2 => \N__40121\,
            in3 => \N__43031\,
            lcout => \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__44295\,
            in1 => \N__39878\,
            in2 => \N__43520\,
            in3 => \N__44934\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__44933\,
            in1 => \N__44296\,
            in2 => \N__43397\,
            in3 => \N__39971\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__33491\,
            in1 => \N__34316\,
            in2 => \_gnd_net_\,
            in3 => \N__37593\,
            lcout => \current_shift_inst.control_input_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110011"
        )
    port map (
            in0 => \N__44948\,
            in1 => \N__44012\,
            in2 => \N__43727\,
            in3 => \N__44298\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__33671\,
            in1 => \N__34415\,
            in2 => \_gnd_net_\,
            in3 => \N__37594\,
            lcout => \current_shift_inst.control_input_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001011111"
        )
    port map (
            in0 => \N__34403\,
            in1 => \_gnd_net_\,
            in2 => \N__37621\,
            in3 => \N__33653\,
            lcout => \current_shift_inst.control_input_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__33635\,
            in1 => \N__34391\,
            in2 => \_gnd_net_\,
            in3 => \N__37598\,
            lcout => \current_shift_inst.control_input_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__37599\,
            in1 => \N__33617\,
            in2 => \_gnd_net_\,
            in3 => \N__34382\,
            lcout => \current_shift_inst.control_input_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__33599\,
            in1 => \N__34373\,
            in2 => \_gnd_net_\,
            in3 => \N__37600\,
            lcout => \current_shift_inst.control_input_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__37601\,
            in1 => \N__34364\,
            in2 => \_gnd_net_\,
            in3 => \N__33581\,
            lcout => \current_shift_inst.control_input_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__33563\,
            in1 => \N__34355\,
            in2 => \_gnd_net_\,
            in3 => \N__37622\,
            lcout => \current_shift_inst.control_input_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__34343\,
            in1 => \N__37624\,
            in2 => \_gnd_net_\,
            in3 => \N__33839\,
            lcout => \current_shift_inst.control_input_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__33821\,
            in1 => \N__34508\,
            in2 => \_gnd_net_\,
            in3 => \N__37623\,
            lcout => \current_shift_inst.control_input_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44417\,
            in1 => \N__40348\,
            in2 => \N__45046\,
            in3 => \N__43355\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.time_passed_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101000011001100"
        )
    port map (
            in0 => \N__42145\,
            in1 => \N__38079\,
            in2 => \N__45506\,
            in3 => \N__42044\,
            lcout => \phase_controller_inst1.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47562\,
            ce => 'H',
            sr => \N__46881\
        );

    \phase_controller_inst1.state_3_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__36693\,
            in1 => \N__38020\,
            in2 => \N__33716\,
            in3 => \N__33787\,
            lcout => state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47562\,
            ce => 'H',
            sr => \N__46881\
        );

    \phase_controller_inst1.start_timer_hc_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101110101010"
        )
    port map (
            in0 => \N__33722\,
            in1 => \N__34637\,
            in2 => \N__34691\,
            in3 => \N__33741\,
            lcout => \phase_controller_inst1.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47562\,
            ce => 'H',
            sr => \N__46881\
        );

    \phase_controller_inst1.start_timer_hc_RNO_0_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36678\,
            in2 => \_gnd_net_\,
            in3 => \N__33708\,
            lcout => \phase_controller_inst1.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_2_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001100"
        )
    port map (
            in0 => \N__33715\,
            in1 => \N__36636\,
            in2 => \N__34619\,
            in3 => \N__36696\,
            lcout => \phase_controller_inst1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47558\,
            ce => 'H',
            sr => \N__46897\
        );

    \current_shift_inst.timer_s1.running_RNII51H_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34529\,
            in2 => \_gnd_net_\,
            in3 => \N__34843\,
            lcout => \current_shift_inst.timer_s1.N_162_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_LC_13_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__34895\,
            in1 => \N__34534\,
            in2 => \_gnd_net_\,
            in3 => \N__34842\,
            lcout => \current_shift_inst.timer_s1.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47553\,
            ce => 'H',
            sr => \N__46905\
        );

    \phase_controller_inst1.S1_LC_13_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36695\,
            lcout => s1_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47551\,
            ce => 'H',
            sr => \N__46910\
        );

    \current_shift_inst.start_timer_s1_LC_13_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__34860\,
            in1 => \N__34893\,
            in2 => \_gnd_net_\,
            in3 => \N__36694\,
            lcout => \current_shift_inst.start_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47551\,
            ce => 'H',
            sr => \N__46910\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__38160\,
            in1 => \N__38213\,
            in2 => \N__37262\,
            in3 => \N__37280\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35615\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47671\,
            ce => \N__36167\,
            sr => \N__46793\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35588\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47671\,
            ce => \N__36167\,
            sr => \N__46793\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37309\,
            in1 => \N__37281\,
            in2 => \_gnd_net_\,
            in3 => \N__48144\,
            lcout => \elapsed_time_ns_1_RNIDC91B_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__33979\,
            in1 => \N__33955\,
            in2 => \N__33893\,
            in3 => \N__33848\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__33847\,
            in1 => \N__33980\,
            in2 => \N__33959\,
            in3 => \N__33889\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_18_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__42599\,
            in1 => \N__48184\,
            in2 => \_gnd_net_\,
            in3 => \N__41855\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47658\,
            ce => \N__45952\,
            sr => \N__46799\
        );

    \phase_controller_inst2.stoper_tr.target_time_19_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48181\,
            in1 => \N__41936\,
            in2 => \_gnd_net_\,
            in3 => \N__41904\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47658\,
            ce => \N__45952\,
            sr => \N__46799\
        );

    \phase_controller_inst2.stoper_tr.target_time_4_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37261\,
            in1 => \N__48185\,
            in2 => \_gnd_net_\,
            in3 => \N__37212\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47658\,
            ce => \N__45952\,
            sr => \N__46799\
        );

    \phase_controller_inst2.stoper_tr.target_time_5_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48182\,
            in1 => \N__38265\,
            in2 => \_gnd_net_\,
            in3 => \N__36896\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47658\,
            ce => \N__45952\,
            sr => \N__46799\
        );

    \phase_controller_inst2.stoper_tr.target_time_7_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48183\,
            in1 => \N__38762\,
            in2 => \_gnd_net_\,
            in3 => \N__38798\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47658\,
            ce => \N__45952\,
            sr => \N__46799\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33881\,
            in2 => \N__34733\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_8_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34145\,
            in1 => \N__35072\,
            in2 => \_gnd_net_\,
            in3 => \N__33875\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \N__47648\,
            ce => 'H',
            sr => \N__46807\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__34142\,
            in1 => \N__35045\,
            in2 => \N__33872\,
            in3 => \N__33860\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \N__47648\,
            ce => 'H',
            sr => \N__46807\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34146\,
            in1 => \N__35015\,
            in2 => \_gnd_net_\,
            in3 => \N__33857\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \N__47648\,
            ce => 'H',
            sr => \N__46807\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34143\,
            in1 => \N__34988\,
            in2 => \_gnd_net_\,
            in3 => \N__33854\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \N__47648\,
            ce => 'H',
            sr => \N__46807\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34147\,
            in1 => \N__34964\,
            in2 => \_gnd_net_\,
            in3 => \N__33851\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \N__47648\,
            ce => 'H',
            sr => \N__46807\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34144\,
            in1 => \N__34937\,
            in2 => \_gnd_net_\,
            in3 => \N__33920\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \N__47648\,
            ce => 'H',
            sr => \N__46807\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34148\,
            in1 => \N__34916\,
            in2 => \_gnd_net_\,
            in3 => \N__33917\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \N__47648\,
            ce => 'H',
            sr => \N__46807\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34179\,
            in1 => \N__35273\,
            in2 => \_gnd_net_\,
            in3 => \N__33914\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_14_9_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \N__47635\,
            ce => 'H',
            sr => \N__46816\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34181\,
            in1 => \N__35252\,
            in2 => \_gnd_net_\,
            in3 => \N__33911\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \N__47635\,
            ce => 'H',
            sr => \N__46816\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34176\,
            in1 => \N__35231\,
            in2 => \_gnd_net_\,
            in3 => \N__33908\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \N__47635\,
            ce => 'H',
            sr => \N__46816\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34182\,
            in1 => \N__35213\,
            in2 => \_gnd_net_\,
            in3 => \N__33905\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \N__47635\,
            ce => 'H',
            sr => \N__46816\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34177\,
            in1 => \N__35182\,
            in2 => \_gnd_net_\,
            in3 => \N__33902\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \N__47635\,
            ce => 'H',
            sr => \N__46816\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34183\,
            in1 => \N__35144\,
            in2 => \_gnd_net_\,
            in3 => \N__33899\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \N__47635\,
            ce => 'H',
            sr => \N__46816\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34178\,
            in1 => \N__35114\,
            in2 => \_gnd_net_\,
            in3 => \N__33896\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \N__47635\,
            ce => 'H',
            sr => \N__46816\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34184\,
            in1 => \N__34767\,
            in2 => \_gnd_net_\,
            in3 => \N__33986\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \N__47635\,
            ce => 'H',
            sr => \N__46816\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34161\,
            in1 => \N__34795\,
            in2 => \_gnd_net_\,
            in3 => \N__33983\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_14_10_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \N__47625\,
            ce => 'H',
            sr => \N__46826\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34165\,
            in1 => \N__33978\,
            in2 => \_gnd_net_\,
            in3 => \N__33962\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \N__47625\,
            ce => 'H',
            sr => \N__46826\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34162\,
            in1 => \N__33954\,
            in2 => \_gnd_net_\,
            in3 => \N__33938\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \N__47625\,
            ce => 'H',
            sr => \N__46826\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34166\,
            in1 => \N__36829\,
            in2 => \_gnd_net_\,
            in3 => \N__33935\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \N__47625\,
            ce => 'H',
            sr => \N__46826\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34163\,
            in1 => \N__36801\,
            in2 => \_gnd_net_\,
            in3 => \N__33932\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\,
            clk => \N__47625\,
            ce => 'H',
            sr => \N__46826\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34167\,
            in1 => \N__36946\,
            in2 => \_gnd_net_\,
            in3 => \N__33929\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\,
            clk => \N__47625\,
            ce => 'H',
            sr => \N__46826\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34164\,
            in1 => \N__36970\,
            in2 => \_gnd_net_\,
            in3 => \N__33926\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\,
            clk => \N__47625\,
            ce => 'H',
            sr => \N__46826\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34168\,
            in1 => \N__45406\,
            in2 => \_gnd_net_\,
            in3 => \N__33923\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\,
            clk => \N__47625\,
            ce => 'H',
            sr => \N__46826\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34169\,
            in1 => \N__45436\,
            in2 => \_gnd_net_\,
            in3 => \N__34223\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_14_11_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\,
            clk => \N__47615\,
            ce => 'H',
            sr => \N__46832\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34173\,
            in1 => \N__45361\,
            in2 => \_gnd_net_\,
            in3 => \N__34220\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\,
            clk => \N__47615\,
            ce => 'H',
            sr => \N__46832\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34170\,
            in1 => \N__45337\,
            in2 => \_gnd_net_\,
            in3 => \N__34217\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\,
            clk => \N__47615\,
            ce => 'H',
            sr => \N__46832\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34174\,
            in1 => \N__45243\,
            in2 => \_gnd_net_\,
            in3 => \N__34214\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\,
            clk => \N__47615\,
            ce => 'H',
            sr => \N__46832\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34171\,
            in1 => \N__45276\,
            in2 => \_gnd_net_\,
            in3 => \N__34211\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\,
            clk => \N__47615\,
            ce => 'H',
            sr => \N__46832\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34175\,
            in1 => \N__34205\,
            in2 => \_gnd_net_\,
            in3 => \N__34187\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\,
            clk => \N__47615\,
            ce => 'H',
            sr => \N__46832\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34172\,
            in1 => \N__34015\,
            in2 => \_gnd_net_\,
            in3 => \N__34034\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47615\,
            ce => 'H',
            sr => \N__46832\
        );

    \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_0_30_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101110"
        )
    port map (
            in0 => \N__39525\,
            in1 => \N__38841\,
            in2 => \N__39170\,
            in3 => \N__38817\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41045\,
            in1 => \N__33997\,
            in2 => \_gnd_net_\,
            in3 => \N__48194\,
            lcout => \elapsed_time_ns_1_RNIVAQBB_0_30\,
            ltout => \elapsed_time_ns_1_RNIVAQBB_0_30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_30_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__48195\,
            in1 => \_gnd_net_\,
            in2 => \N__34298\,
            in3 => \N__41046\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47604\,
            ce => \N__47208\,
            sr => \N__46840\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38342\,
            in1 => \N__34291\,
            in2 => \_gnd_net_\,
            in3 => \N__48193\,
            lcout => \elapsed_time_ns_1_RNI0CQBB_0_31\,
            ltout => \elapsed_time_ns_1_RNI0CQBB_0_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_31_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__48196\,
            in1 => \_gnd_net_\,
            in2 => \N__34280\,
            in3 => \N__38343\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47604\,
            ce => \N__47208\,
            sr => \N__46840\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__38842\,
            in1 => \N__39169\,
            in2 => \N__38824\,
            in3 => \N__39526\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_13_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__34277\,
            in1 => \N__48197\,
            in2 => \_gnd_net_\,
            in3 => \N__38444\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47604\,
            ce => \N__47208\,
            sr => \N__46840\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34261\,
            in2 => \N__34250\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_13_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45150\,
            in2 => \N__43610\,
            in3 => \N__45071\,
            lcout => \current_shift_inst.un38_control_input_5_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__45072\,
            in1 => \N__44552\,
            in2 => \N__34238\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un38_control_input_5_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34460\,
            in2 => \N__44775\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44556\,
            in2 => \N__36086\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36074\,
            in2 => \N__44776\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44560\,
            in2 => \N__43628\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36320\,
            in2 => \N__44777\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44564\,
            in2 => \N__36311\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_14_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36344\,
            in2 => \N__44778\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44568\,
            in2 => \N__36437\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36053\,
            in2 => \N__44779\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44572\,
            in2 => \N__34307\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36302\,
            in2 => \N__44780\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44576\,
            in2 => \N__36335\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36326\,
            in2 => \N__44781\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44782\,
            in2 => \N__36296\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_15_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34451\,
            in2 => \N__44969\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44786\,
            in2 => \N__36410\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36428\,
            in2 => \N__44970\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44790\,
            in2 => \N__36422\,
            in3 => \N__34319\,
            lcout => \current_shift_inst.un38_control_input_0_s0_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42428\,
            in2 => \N__44971\,
            in3 => \N__34427\,
            lcout => \current_shift_inst.un38_control_input_0_s0_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44794\,
            in2 => \N__34424\,
            in3 => \N__34406\,
            lcout => \current_shift_inst.un38_control_input_0_s0_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36392\,
            in2 => \N__44972\,
            in3 => \N__34394\,
            lcout => \current_shift_inst.un38_control_input_0_s0_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44798\,
            in2 => \N__36386\,
            in3 => \N__34385\,
            lcout => \current_shift_inst.un38_control_input_0_s0_24\,
            ltout => OPEN,
            carryin => \bfn_14_16_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36458\,
            in2 => \N__44973\,
            in3 => \N__34376\,
            lcout => \current_shift_inst.un38_control_input_0_s0_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44802\,
            in2 => \N__36401\,
            in3 => \N__34367\,
            lcout => \current_shift_inst.un38_control_input_0_s0_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36365\,
            in2 => \N__44974\,
            in3 => \N__34358\,
            lcout => \current_shift_inst.un38_control_input_0_s0_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44806\,
            in2 => \N__36374\,
            in3 => \N__34346\,
            lcout => \current_shift_inst.un38_control_input_0_s0_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34466\,
            in2 => \N__44975\,
            in3 => \N__34334\,
            lcout => \current_shift_inst.un38_control_input_0_s0_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44810\,
            in2 => \N__44078\,
            in3 => \N__34499\,
            lcout => \current_shift_inst.un38_control_input_0_s0_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001101010011"
        )
    port map (
            in0 => \N__42479\,
            in1 => \N__34496\,
            in2 => \N__37633\,
            in3 => \N__34484\,
            lcout => \current_shift_inst.control_input_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39434\,
            lcout => \current_shift_inst.un4_control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39474\,
            lcout => \current_shift_inst.un4_control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44400\,
            in1 => \N__44008\,
            in2 => \N__45043\,
            in3 => \N__43726\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44398\,
            in1 => \N__39273\,
            in2 => \N__45044\,
            in3 => \N__42191\,
            lcout => \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__42998\,
            in1 => \N__44979\,
            in2 => \N__43967\,
            in3 => \N__44399\,
            lcout => \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__40191\,
            in1 => \N__44407\,
            in2 => \N__45045\,
            in3 => \N__43262\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39596\,
            lcout => \current_shift_inst.un4_control_input_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40052\,
            lcout => \current_shift_inst.un4_control_input_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39642\,
            lcout => \current_shift_inst.un4_control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_tr_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__34690\,
            in1 => \N__34544\,
            in2 => \N__45539\,
            in3 => \N__38024\,
            lcout => \phase_controller_inst1.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47563\,
            ce => 'H',
            sr => \N__46882\
        );

    \phase_controller_inst1.state_0_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001000100010"
        )
    port map (
            in0 => \N__38046\,
            in1 => \N__38080\,
            in2 => \N__34574\,
            in3 => \N__36576\,
            lcout => \phase_controller_inst1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47563\,
            ce => 'H',
            sr => \N__46882\
        );

    \phase_controller_inst1.state_1_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__36577\,
            in1 => \N__34572\,
            in2 => \_gnd_net_\,
            in3 => \N__34633\,
            lcout => \phase_controller_inst1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47563\,
            ce => 'H',
            sr => \N__46882\
        );

    \phase_controller_inst1.stoper_hc.time_passed_RNIE87F_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36634\,
            in2 => \_gnd_net_\,
            in3 => \N__34614\,
            lcout => \phase_controller_inst1.time_passed_RNIE87F\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIUKI8_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34535\,
            lcout => \current_shift_inst.timer_s1.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_tr_RNO_0_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__36635\,
            in1 => \N__34615\,
            in2 => \N__34573\,
            in3 => \N__36578\,
            lcout => \phase_controller_inst1.start_timer_tr_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIEOIK_LC_14_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__34892\,
            in1 => \N__34533\,
            in2 => \_gnd_net_\,
            in3 => \N__34838\,
            lcout => \current_shift_inst.timer_s1.N_163_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.stop_timer_s1_LC_14_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__34894\,
            in1 => \N__36703\,
            in2 => \N__34844\,
            in3 => \N__34861\,
            lcout => \current_shift_inst.stop_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47554\,
            ce => 'H',
            sr => \N__46906\
        );

    \phase_controller_inst1.S2_LC_14_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__36587\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => s2_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47550\,
            ce => 'H',
            sr => \N__46915\
        );

    \phase_controller_inst1.stoper_tr.target_time_3_LC_15_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__38120\,
            in1 => \N__38159\,
            in2 => \_gnd_net_\,
            in3 => \N__48180\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47690\,
            ce => \N__47219\,
            sr => \N__46785\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100011001110"
        )
    port map (
            in0 => \N__34750\,
            in1 => \N__36863\,
            in2 => \N__34780\,
            in3 => \N__34802\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101000101"
        )
    port map (
            in0 => \N__34801\,
            in1 => \N__34751\,
            in2 => \N__34781\,
            in3 => \N__36862\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_16_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41454\,
            in1 => \N__41420\,
            in2 => \_gnd_net_\,
            in3 => \N__48147\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47679\,
            ce => \N__45953\,
            sr => \N__46788\
        );

    \phase_controller_inst2.stoper_tr.target_time_15_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42518\,
            in1 => \N__42545\,
            in2 => \_gnd_net_\,
            in3 => \N__48146\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47679\,
            ce => \N__45953\,
            sr => \N__46788\
        );

    \phase_controller_inst2.stoper_tr.target_time_1_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48145\,
            in1 => \N__37305\,
            in2 => \_gnd_net_\,
            in3 => \N__37282\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47679\,
            ce => \N__45953\,
            sr => \N__46788\
        );

    \phase_controller_inst2.stoper_tr.target_time_2_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__38191\,
            in1 => \N__38217\,
            in2 => \_gnd_net_\,
            in3 => \N__48148\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47679\,
            ce => \N__45953\,
            sr => \N__46788\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34742\,
            in2 => \N__34700\,
            in3 => \N__34729\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_15_7_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35071\,
            in1 => \N__35060\,
            in2 => \N__35054\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36875\,
            in2 => \N__35033\,
            in3 => \N__35044\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35024\,
            in2 => \N__35003\,
            in3 => \N__35014\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34994\,
            in2 => \N__34976\,
            in3 => \N__34987\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36869\,
            in2 => \N__34952\,
            in3 => \N__34963\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34943\,
            in2 => \N__34925\,
            in3 => \N__34936\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37007\,
            in2 => \N__34904\,
            in3 => \N__34915\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_7\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35261\,
            in2 => \N__37001\,
            in3 => \N__35272\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_15_8_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36992\,
            in2 => \N__35240\,
            in3 => \N__35251\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35219\,
            in2 => \N__36905\,
            in3 => \N__35230\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35201\,
            in2 => \N__37106\,
            in3 => \N__35212\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35195\,
            in2 => \N__35168\,
            in3 => \N__35183\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35159\,
            in2 => \N__35132\,
            in3 => \N__35143\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35123\,
            in2 => \N__35102\,
            in3 => \N__35113\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35093\,
            in2 => \N__35084\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_15\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35369\,
            in2 => \N__35360\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_9_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36773\,
            in2 => \N__36851\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36932\,
            in2 => \N__36986\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_20\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45392\,
            in2 => \N__43781\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_22\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45380\,
            in2 => \N__45323\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_24\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45302\,
            in2 => \N__45731\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_26\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35345\,
            in2 => \N__35336\,
            in3 => \N__35303\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_28\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35300\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35611\,
            in2 => \N__35554\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\,
            ltout => OPEN,
            carryin => \bfn_15_10_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__47636\,
            ce => \N__36166\,
            sr => \N__46817\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35527\,
            in2 => \N__35587\,
            in3 => \N__35558\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__47636\,
            ce => \N__36166\,
            sr => \N__46817\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35503\,
            in2 => \N__35555\,
            in3 => \N__35531\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__47636\,
            ce => \N__36166\,
            sr => \N__46817\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35528\,
            in2 => \N__35479\,
            in3 => \N__35510\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__47636\,
            ce => \N__36166\,
            sr => \N__46817\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35451\,
            in2 => \N__35507\,
            in3 => \N__35483\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__47636\,
            ce => \N__36166\,
            sr => \N__46817\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35428\,
            in2 => \N__35480\,
            in3 => \N__35456\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__47636\,
            ce => \N__36166\,
            sr => \N__46817\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35452\,
            in2 => \N__35405\,
            in3 => \N__35435\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__47636\,
            ce => \N__36166\,
            sr => \N__46817\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35824\,
            in2 => \N__35432\,
            in3 => \N__35408\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__47636\,
            ce => \N__36166\,
            sr => \N__46817\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35794\,
            in2 => \N__35404\,
            in3 => \N__35372\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\,
            ltout => OPEN,
            carryin => \bfn_15_11_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__47626\,
            ce => \N__36158\,
            sr => \N__46827\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35770\,
            in2 => \N__35825\,
            in3 => \N__35798\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__47626\,
            ce => \N__36158\,
            sr => \N__46827\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35795\,
            in2 => \N__35746\,
            in3 => \N__35777\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__47626\,
            ce => \N__36158\,
            sr => \N__46827\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35716\,
            in2 => \N__35774\,
            in3 => \N__35750\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__47626\,
            ce => \N__36158\,
            sr => \N__46827\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35689\,
            in2 => \N__35747\,
            in3 => \N__35723\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__47626\,
            ce => \N__36158\,
            sr => \N__46827\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35664\,
            in2 => \N__35720\,
            in3 => \N__35696\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__47626\,
            ce => \N__36158\,
            sr => \N__46827\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35644\,
            in2 => \N__35693\,
            in3 => \N__35669\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__47626\,
            ce => \N__36158\,
            sr => \N__46827\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35665\,
            in2 => \N__36041\,
            in3 => \N__35648\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__47626\,
            ce => \N__36158\,
            sr => \N__46827\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36000\,
            in2 => \N__35645\,
            in3 => \N__35618\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\,
            ltout => OPEN,
            carryin => \bfn_15_12_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__47616\,
            ce => \N__36159\,
            sr => \N__46833\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35977\,
            in2 => \N__36040\,
            in3 => \N__36008\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__47616\,
            ce => \N__36159\,
            sr => \N__46833\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35956\,
            in2 => \N__36005\,
            in3 => \N__35981\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__47616\,
            ce => \N__36159\,
            sr => \N__46833\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35978\,
            in2 => \N__35936\,
            in3 => \N__35960\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__47616\,
            ce => \N__36159\,
            sr => \N__46833\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35957\,
            in2 => \N__35908\,
            in3 => \N__35939\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__47616\,
            ce => \N__36159\,
            sr => \N__46833\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35935\,
            in2 => \N__35881\,
            in3 => \N__35912\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__47616\,
            ce => \N__36159\,
            sr => \N__46833\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35851\,
            in2 => \N__35909\,
            in3 => \N__35885\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__47616\,
            ce => \N__36159\,
            sr => \N__46833\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36286\,
            in2 => \N__35882\,
            in3 => \N__35858\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__47616\,
            ce => \N__36159\,
            sr => \N__46833\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36234\,
            in2 => \N__35855\,
            in3 => \N__35828\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\,
            ltout => OPEN,
            carryin => \bfn_15_13_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__47605\,
            ce => \N__36157\,
            sr => \N__46841\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36193\,
            in2 => \N__36287\,
            in3 => \N__36257\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__47605\,
            ce => \N__36157\,
            sr => \N__46841\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36254\,
            in2 => \N__36239\,
            in3 => \N__36215\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__47605\,
            ce => \N__36157\,
            sr => \N__46841\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36212\,
            in2 => \N__36197\,
            in3 => \N__36173\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__47605\,
            ce => \N__36157\,
            sr => \N__46841\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36170\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47605\,
            ce => \N__36157\,
            sr => \N__46841\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__44625\,
            in1 => \N__44278\,
            in2 => \N__39823\,
            in3 => \N__42845\,
            lcout => \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__44280\,
            in1 => \N__39407\,
            in2 => \N__42890\,
            in3 => \N__44623\,
            lcout => \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__44624\,
            in1 => \N__44281\,
            in2 => \N__39824\,
            in3 => \N__42844\,
            lcout => \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__44279\,
            in1 => \N__44626\,
            in2 => \N__42760\,
            in3 => \N__39447\,
            lcout => \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__44622\,
            in1 => \N__44282\,
            in2 => \N__39619\,
            in3 => \N__42632\,
            lcout => \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__39406\,
            in1 => \N__44277\,
            in2 => \N__42889\,
            in3 => \N__44627\,
            lcout => \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__45194\,
            in1 => \N__45211\,
            in2 => \_gnd_net_\,
            in3 => \N__42380\,
            lcout => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44361\,
            in1 => \N__39489\,
            in2 => \N__44996\,
            in3 => \N__42715\,
            lcout => \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__44063\,
            in1 => \N__44364\,
            in2 => \N__43117\,
            in3 => \N__44829\,
            lcout => \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__44365\,
            in1 => \N__43069\,
            in2 => \N__44994\,
            in3 => \N__39567\,
            lcout => \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__42803\,
            in1 => \N__44834\,
            in2 => \N__39373\,
            in3 => \N__44359\,
            lcout => \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44360\,
            in1 => \N__39448\,
            in2 => \N__44995\,
            in3 => \N__42761\,
            lcout => \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__43151\,
            in1 => \N__44828\,
            in2 => \N__39758\,
            in3 => \N__44363\,
            lcout => \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001111"
        )
    port map (
            in0 => \N__44833\,
            in1 => \N__43027\,
            in2 => \N__44419\,
            in3 => \N__40120\,
            lcout => \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__42670\,
            in1 => \N__44827\,
            in2 => \N__39665\,
            in3 => \N__44362\,
            lcout => \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110011"
        )
    port map (
            in0 => \N__44852\,
            in1 => \N__43900\,
            in2 => \N__42932\,
            in3 => \N__44402\,
            lcout => \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44403\,
            in1 => \N__39876\,
            in2 => \N__44998\,
            in3 => \N__43516\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__44851\,
            in1 => \N__44401\,
            in2 => \N__39926\,
            in3 => \N__42955\,
            lcout => \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44406\,
            in1 => \N__40192\,
            in2 => \N__44999\,
            in3 => \N__43261\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__42381\,
            in1 => \N__42927\,
            in2 => \_gnd_net_\,
            in3 => \N__43899\,
            lcout => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44404\,
            in1 => \N__39970\,
            in2 => \N__44997\,
            in3 => \N__43396\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__44850\,
            in1 => \N__44405\,
            in2 => \N__40352\,
            in3 => \N__43348\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__44389\,
            in1 => \N__45033\,
            in2 => \N__43754\,
            in3 => \N__40260\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \N__45031\,
            in1 => \N__40303\,
            in2 => \N__44429\,
            in3 => \N__43216\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \N__45032\,
            in1 => \N__40304\,
            in2 => \N__44428\,
            in3 => \N__43217\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39350\,
            lcout => \current_shift_inst.un4_control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__44388\,
            in1 => \N__40065\,
            in2 => \N__43310\,
            in3 => \N__45034\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40567\,
            in2 => \N__40153\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_3\,
            ltout => OPEN,
            carryin => \bfn_15_18_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            clk => \N__47572\,
            ce => \N__43570\,
            sr => \N__46867\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43595\,
            in2 => \N__40547\,
            in3 => \N__36452\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            clk => \N__47572\,
            ce => \N__43570\,
            sr => \N__46867\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40568\,
            in2 => \N__40516\,
            in3 => \N__36449\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            clk => \N__47572\,
            ce => \N__43570\,
            sr => \N__46867\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40546\,
            in2 => \N__40489\,
            in3 => \N__36446\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            clk => \N__47572\,
            ce => \N__43570\,
            sr => \N__46867\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40462\,
            in2 => \N__40517\,
            in3 => \N__36443\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            clk => \N__47572\,
            ce => \N__43570\,
            sr => \N__46867\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40441\,
            in2 => \N__40490\,
            in3 => \N__36440\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            clk => \N__47572\,
            ce => \N__43570\,
            sr => \N__46867\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40463\,
            in2 => \N__40420\,
            in3 => \N__36497\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            clk => \N__47572\,
            ce => \N__43570\,
            sr => \N__46867\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40442\,
            in2 => \N__40387\,
            in3 => \N__36494\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            clk => \N__47572\,
            ce => \N__43570\,
            sr => \N__46867\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40783\,
            in2 => \N__40421\,
            in3 => \N__36491\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_11\,
            ltout => OPEN,
            carryin => \bfn_15_19_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            clk => \N__47567\,
            ce => \N__43569\,
            sr => \N__46871\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40762\,
            in2 => \N__40388\,
            in3 => \N__36488\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            clk => \N__47567\,
            ce => \N__43569\,
            sr => \N__46871\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40784\,
            in2 => \N__40742\,
            in3 => \N__36485\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            clk => \N__47567\,
            ce => \N__43569\,
            sr => \N__46871\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40763\,
            in2 => \N__40715\,
            in3 => \N__36482\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            clk => \N__47567\,
            ce => \N__43569\,
            sr => \N__46871\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40741\,
            in2 => \N__40687\,
            in3 => \N__36479\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            clk => \N__47567\,
            ce => \N__43569\,
            sr => \N__46871\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40714\,
            in2 => \N__40660\,
            in3 => \N__36476\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            clk => \N__47567\,
            ce => \N__43569\,
            sr => \N__46871\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40633\,
            in2 => \N__40688\,
            in3 => \N__36473\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            clk => \N__47567\,
            ce => \N__43569\,
            sr => \N__46871\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40600\,
            in2 => \N__40661\,
            in3 => \N__36524\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            clk => \N__47567\,
            ce => \N__43569\,
            sr => \N__46871\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41017\,
            in2 => \N__40634\,
            in3 => \N__36521\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_19\,
            ltout => OPEN,
            carryin => \bfn_15_20_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            clk => \N__47565\,
            ce => \N__43568\,
            sr => \N__46876\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40993\,
            in2 => \N__40601\,
            in3 => \N__36518\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            clk => \N__47565\,
            ce => \N__43568\,
            sr => \N__46876\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41018\,
            in2 => \N__40969\,
            in3 => \N__36515\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            clk => \N__47565\,
            ce => \N__43568\,
            sr => \N__46876\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40942\,
            in2 => \N__40997\,
            in3 => \N__36512\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            clk => \N__47565\,
            ce => \N__43568\,
            sr => \N__46876\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40921\,
            in2 => \N__40970\,
            in3 => \N__36509\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            clk => \N__47565\,
            ce => \N__43568\,
            sr => \N__46876\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40943\,
            in2 => \N__40900\,
            in3 => \N__36506\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            clk => \N__47565\,
            ce => \N__43568\,
            sr => \N__46876\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40922\,
            in2 => \N__40874\,
            in3 => \N__36503\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            clk => \N__47565\,
            ce => \N__43568\,
            sr => \N__46876\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40837\,
            in2 => \N__40901\,
            in3 => \N__36500\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            clk => \N__47565\,
            ce => \N__43568\,
            sr => \N__46876\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40804\,
            in2 => \N__40873\,
            in3 => \N__36764\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_27\,
            ltout => OPEN,
            carryin => \bfn_15_21_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            clk => \N__47564\,
            ce => \N__43567\,
            sr => \N__46883\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41395\,
            in2 => \N__40838\,
            in3 => \N__36761\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            clk => \N__47564\,
            ce => \N__43567\,
            sr => \N__46883\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40805\,
            in2 => \N__41375\,
            in3 => \N__36758\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            clk => \N__47564\,
            ce => \N__43567\,
            sr => \N__46883\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41396\,
            in2 => \N__41216\,
            in3 => \N__36755\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\,
            clk => \N__47564\,
            ce => \N__43567\,
            sr => \N__46883\
        );

    \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36752\,
            lcout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.T12_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__36739\,
            in1 => \N__36579\,
            in2 => \_gnd_net_\,
            in3 => \N__36650\,
            lcout => \T12_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47561\,
            ce => 'H',
            sr => \N__46893\
        );

    \phase_controller_inst1.T45_LC_15_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__36710\,
            in1 => \N__38056\,
            in2 => \_gnd_net_\,
            in3 => \N__36721\,
            lcout => \T45_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47559\,
            ce => 'H',
            sr => \N__46898\
        );

    \phase_controller_inst1.T01_LC_15_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__36598\,
            in1 => \N__36709\,
            in2 => \_gnd_net_\,
            in3 => \N__36649\,
            lcout => \T01_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47559\,
            ce => 'H',
            sr => \N__46898\
        );

    \phase_controller_inst1.T23_LC_15_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100001010"
        )
    port map (
            in0 => \N__36535\,
            in1 => \_gnd_net_\,
            in2 => \N__38060\,
            in3 => \N__36586\,
            lcout => \T23_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47559\,
            ce => 'H',
            sr => \N__46898\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_16_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38266\,
            in1 => \N__36889\,
            in2 => \_gnd_net_\,
            in3 => \N__48022\,
            lcout => \elapsed_time_ns_1_RNIHG91B_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_5_LC_16_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38267\,
            in1 => \N__36888\,
            in2 => \_gnd_net_\,
            in3 => \N__48023\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47696\,
            ce => \N__47209\,
            sr => \N__46783\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_LC_16_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38309\,
            in1 => \N__38097\,
            in2 => \_gnd_net_\,
            in3 => \N__48024\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47696\,
            ce => \N__47209\,
            sr => \N__46783\
        );

    \phase_controller_inst2.stoper_tr.target_time_3_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48006\,
            in1 => \N__38118\,
            in2 => \_gnd_net_\,
            in3 => \N__38161\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47691\,
            ce => \N__45955\,
            sr => \N__46786\
        );

    \phase_controller_inst2.stoper_tr.target_time_21_LC_16_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41111\,
            in1 => \N__38414\,
            in2 => \_gnd_net_\,
            in3 => \N__48009\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47691\,
            ce => \N__45955\,
            sr => \N__46786\
        );

    \phase_controller_inst2.stoper_tr.target_time_6_LC_16_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48007\,
            in1 => \N__38301\,
            in2 => \_gnd_net_\,
            in3 => \N__38098\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47691\,
            ce => \N__45955\,
            sr => \N__46786\
        );

    \phase_controller_inst2.stoper_tr.target_time_17_LC_16_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41765\,
            in1 => \N__41738\,
            in2 => \_gnd_net_\,
            in3 => \N__48008\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47691\,
            ce => \N__45955\,
            sr => \N__46786\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001100"
        )
    port map (
            in0 => \N__36835\,
            in1 => \N__36785\,
            in2 => \N__36814\,
            in3 => \N__37016\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__37015\,
            in1 => \N__36836\,
            in2 => \N__36815\,
            in3 => \N__36784\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_20_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47995\,
            in1 => \N__38866\,
            in2 => \_gnd_net_\,
            in3 => \N__38911\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47680\,
            ce => \N__45956\,
            sr => \N__46789\
        );

    \phase_controller_inst2.stoper_tr.target_time_8_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47996\,
            in1 => \N__38520\,
            in2 => \_gnd_net_\,
            in3 => \N__38498\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47680\,
            ce => \N__45956\,
            sr => \N__46789\
        );

    \phase_controller_inst2.stoper_tr.target_time_9_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47997\,
            in1 => \N__41834\,
            in2 => \_gnd_net_\,
            in3 => \N__41809\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47680\,
            ce => \N__45956\,
            sr => \N__46789\
        );

    \phase_controller_inst2.stoper_tr.target_time_10_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__37040\,
            in1 => \N__37082\,
            in2 => \_gnd_net_\,
            in3 => \N__47998\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47680\,
            ce => \N__45956\,
            sr => \N__46789\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__36976\,
            in1 => \N__36952\,
            in2 => \N__36917\,
            in3 => \N__36926\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__36925\,
            in1 => \N__36977\,
            in2 => \N__36956\,
            in3 => \N__36913\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_22_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48010\,
            in1 => \N__38558\,
            in2 => \_gnd_net_\,
            in3 => \N__41149\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47672\,
            ce => \N__45957\,
            sr => \N__46794\
        );

    \phase_controller_inst2.stoper_tr.target_time_23_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48004\,
            in1 => \N__41692\,
            in2 => \_gnd_net_\,
            in3 => \N__41674\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47672\,
            ce => \N__45957\,
            sr => \N__46794\
        );

    \phase_controller_inst2.stoper_tr.target_time_11_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__37064\,
            in1 => \N__37097\,
            in2 => \_gnd_net_\,
            in3 => \N__48005\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47672\,
            ce => \N__45957\,
            sr => \N__46794\
        );

    \phase_controller_inst2.stoper_tr.target_time_12_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48003\,
            in1 => \N__38698\,
            in2 => \_gnd_net_\,
            in3 => \N__38735\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47672\,
            ce => \N__45957\,
            sr => \N__46794\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__37059\,
            in1 => \_gnd_net_\,
            in2 => \N__48179\,
            in3 => \N__37096\,
            lcout => \elapsed_time_ns_1_RNIU7OBB_0_11\,
            ltout => \elapsed_time_ns_1_RNIU7OBB_0_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_11_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37060\,
            in2 => \N__37085\,
            in3 => \N__48096\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47659\,
            ce => \N__47203\,
            sr => \N__46800\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48091\,
            in1 => \N__37032\,
            in2 => \_gnd_net_\,
            in3 => \N__37078\,
            lcout => \elapsed_time_ns_1_RNIT6OBB_0_10\,
            ltout => \elapsed_time_ns_1_RNIT6OBB_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_10_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__37033\,
            in1 => \_gnd_net_\,
            in2 => \N__37067\,
            in3 => \N__48095\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47659\,
            ce => \N__47203\,
            sr => \N__46800\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__37058\,
            in1 => \N__37031\,
            in2 => \N__38736\,
            in3 => \N__41791\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_12_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38738\,
            in1 => \N__38697\,
            in2 => \_gnd_net_\,
            in3 => \N__48097\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47659\,
            ce => \N__47203\,
            sr => \N__46800\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110101000100"
        )
    port map (
            in0 => \N__39053\,
            in1 => \N__38395\,
            in2 => \N__39077\,
            in3 => \N__37322\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_20_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48099\,
            in1 => \N__38867\,
            in2 => \_gnd_net_\,
            in3 => \N__38903\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47649\,
            ce => \N__47171\,
            sr => \N__46808\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__37321\,
            in1 => \N__39052\,
            in2 => \N__38399\,
            in3 => \N__39076\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_1_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48098\,
            in1 => \N__37313\,
            in2 => \_gnd_net_\,
            in3 => \N__37289\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47649\,
            ce => \N__47171\,
            sr => \N__46808\
        );

    \phase_controller_inst1.stoper_tr.target_time_2_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38228\,
            in1 => \N__38192\,
            in2 => \_gnd_net_\,
            in3 => \N__48100\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47649\,
            ce => \N__47171\,
            sr => \N__46808\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__37247\,
            in1 => \N__37220\,
            in2 => \_gnd_net_\,
            in3 => \N__48101\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47649\,
            ce => \N__47171\,
            sr => \N__46808\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37184\,
            in2 => \N__37193\,
            in3 => \N__38670\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_16_11_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37178\,
            in2 => \N__37172\,
            in3 => \N__38647\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38632\,
            in1 => \N__37163\,
            in2 => \N__37151\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38617\,
            in1 => \N__37133\,
            in2 => \N__37142\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37127\,
            in2 => \N__37115\,
            in3 => \N__39031\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__39016\,
            in1 => \N__37433\,
            in2 => \N__37424\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__39001\,
            in1 => \N__38534\,
            in2 => \N__37415\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37406\,
            in2 => \N__38471\,
            in3 => \N__38986\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_7\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37400\,
            in2 => \N__41780\,
            in3 => \N__38971\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_16_12_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37382\,
            in2 => \N__37394\,
            in3 => \N__38956\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37376\,
            in2 => \N__37367\,
            in3 => \N__38941\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37358\,
            in2 => \N__37349\,
            in3 => \N__38926\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__39133\,
            in1 => \N__37328\,
            in2 => \N__37340\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__39118\,
            in1 => \N__41471\,
            in2 => \N__37478\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42488\,
            in2 => \N__37466\,
            in3 => \N__39103\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41540\,
            in2 => \N__41618\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_15\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41996\,
            in2 => \N__41951\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_13_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37457\,
            in2 => \N__37448\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38588\,
            in2 => \N__38573\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46379\,
            in2 => \N__46460\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45566\,
            in2 => \N__46295\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45647\,
            in2 => \N__45578\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42110\,
            in2 => \N__37526\,
            in3 => \N__37511\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37508\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_0_c_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45079\,
            in2 => \N__37505\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_14_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37947\,
            in2 => \N__37487\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_0\,
            carryout => \current_shift_inst.un10_control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39293\,
            in2 => \N__37994\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_1\,
            carryout => \current_shift_inst.un10_control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37951\,
            in2 => \N__39248\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_2\,
            carryout => \current_shift_inst.un10_control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39380\,
            in2 => \N__37995\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_3\,
            carryout => \current_shift_inst.un10_control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37955\,
            in2 => \N__39788\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_4\,
            carryout => \current_shift_inst.un10_control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39287\,
            in2 => \N__37996\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_5\,
            carryout => \current_shift_inst.un10_control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37959\,
            in2 => \N__39335\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_6\,
            carryout => \current_shift_inst.un10_control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37943\,
            in2 => \N__39416\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_15_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39458\,
            in2 => \N__37993\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_8\,
            carryout => \current_shift_inst.un10_control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37931\,
            in2 => \N__39629\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_9\,
            carryout => \current_shift_inst.un10_control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39578\,
            in2 => \N__37990\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_10\,
            carryout => \current_shift_inst.un10_control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37935\,
            in2 => \N__39674\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_11\,
            carryout => \current_shift_inst.un10_control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39716\,
            in2 => \N__37991\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_12\,
            carryout => \current_shift_inst.un10_control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37939\,
            in2 => \N__39779\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_13\,
            carryout => \current_shift_inst.un10_control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39536\,
            in2 => \N__37992\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_14\,
            carryout => \current_shift_inst.un10_control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37761\,
            in2 => \N__40082\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_16_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39977\,
            in2 => \N__37843\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_16\,
            carryout => \current_shift_inst.un10_control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37765\,
            in2 => \N__39887\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_17\,
            carryout => \current_shift_inst.un10_control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37532\,
            in2 => \N__37844\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_18\,
            carryout => \current_shift_inst.un10_control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37769\,
            in2 => \N__39842\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_19\,
            carryout => \current_shift_inst.un10_control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39932\,
            in2 => \N__37845\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_20\,
            carryout => \current_shift_inst.un10_control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37773\,
            in2 => \N__39986\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_21\,
            carryout => \current_shift_inst.un10_control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39938\,
            in2 => \N__37846\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_22\,
            carryout => \current_shift_inst.un10_control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40310\,
            in2 => \N__37997\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_17_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37963\,
            in2 => \N__40031\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_24\,
            carryout => \current_shift_inst.un10_control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40160\,
            in2 => \N__37998\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_25\,
            carryout => \current_shift_inst.un10_control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37967\,
            in2 => \N__40277\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_26\,
            carryout => \current_shift_inst.un10_control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40268\,
            in2 => \N__37999\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_27\,
            carryout => \current_shift_inst.un10_control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37971\,
            in2 => \N__39833\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_28\,
            carryout => \current_shift_inst.un10_control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43694\,
            in2 => \N__38000\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_29\,
            carryout => \current_shift_inst.un10_control_input_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44390\,
            in2 => \_gnd_net_\,
            in3 => \N__37637\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39266\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39391\,
            lcout => \current_shift_inst.un4_control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39804\,
            lcout => \current_shift_inst.un4_control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39306\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39687\,
            lcout => \current_shift_inst.un4_control_input_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40095\,
            lcout => \current_shift_inst.un4_control_input_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39552\,
            lcout => \current_shift_inst.un4_control_input_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39999\,
            lcout => \current_shift_inst.un4_control_input_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.time_passed_RNI7NN7_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__38081\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38055\,
            lcout => \phase_controller_inst1.time_passed_RNI7NN7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42444\,
            lcout => \current_shift_inst.un4_control_input_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39727\,
            lcout => \current_shift_inst.un4_control_input_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39951\,
            lcout => \current_shift_inst.un4_control_input_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40288\,
            lcout => \current_shift_inst.un4_control_input_1_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39900\,
            lcout => \current_shift_inst.un4_control_input_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39860\,
            lcout => \current_shift_inst.un4_control_input_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40328\,
            lcout => \current_shift_inst.un4_control_input_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40178\,
            lcout => \current_shift_inst.un4_control_input_1_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40248\,
            lcout => \current_shift_inst.un4_control_input_1_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_17_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__38184\,
            in1 => \N__38227\,
            in2 => \_gnd_net_\,
            in3 => \N__48019\,
            lcout => \elapsed_time_ns_1_RNIED91B_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_17_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48020\,
            in1 => \N__38119\,
            in2 => \_gnd_net_\,
            in3 => \N__38165\,
            lcout => \elapsed_time_ns_1_RNIFE91B_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_17_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__38099\,
            in1 => \N__38308\,
            in2 => \_gnd_net_\,
            in3 => \N__48021\,
            lcout => \elapsed_time_ns_1_RNIIH91B_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_17_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41906\,
            in1 => \N__42596\,
            in2 => \N__41741\,
            in3 => \N__38912\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_17_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41113\,
            in1 => \N__38413\,
            in2 => \_gnd_net_\,
            in3 => \N__47986\,
            lcout => \elapsed_time_ns_1_RNIV9PBB_0_21\,
            ltout => \elapsed_time_ns_1_RNIV9PBB_0_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_21_LC_17_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__47987\,
            in1 => \_gnd_net_\,
            in2 => \N__38402\,
            in3 => \N__41114\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47697\,
            ce => \N__47229\,
            sr => \N__46784\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__41069\,
            in1 => \N__41024\,
            in2 => \N__38381\,
            in3 => \N__38423\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_17_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__45704\,
            in1 => \N__48284\,
            in2 => \_gnd_net_\,
            in3 => \N__38369\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__38357\,
            in1 => \N__38594\,
            in2 => \N__38321\,
            in3 => \N__38318\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3\,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38500\,
            in2 => \N__38312\,
            in3 => \N__38521\,
            lcout => \elapsed_time_ns_1_RNIKJ91B_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__38499\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38795\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_17_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__38300\,
            in1 => \N__38264\,
            in2 => \N__38231\,
            in3 => \N__38603\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41693\,
            in1 => \N__41673\,
            in2 => \_gnd_net_\,
            in3 => \N__47988\,
            lcout => \elapsed_time_ns_1_RNI1CPBB_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001100"
        )
    port map (
            in0 => \N__39235\,
            in1 => \N__41630\,
            in2 => \N__39212\,
            in3 => \N__38543\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__38542\,
            in1 => \N__39208\,
            in2 => \N__39239\,
            in3 => \N__41629\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41147\,
            in1 => \N__38557\,
            in2 => \_gnd_net_\,
            in3 => \N__47982\,
            lcout => \elapsed_time_ns_1_RNI0BPBB_0_22\,
            ltout => \elapsed_time_ns_1_RNI0BPBB_0_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_22_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__47983\,
            in1 => \_gnd_net_\,
            in2 => \N__38546\,
            in3 => \N__41148\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47681\,
            ce => \N__47220\,
            sr => \N__46790\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__38754\,
            in1 => \N__38797\,
            in2 => \_gnd_net_\,
            in3 => \N__47985\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47681\,
            ce => \N__47220\,
            sr => \N__46790\
        );

    \phase_controller_inst1.stoper_tr.target_time_8_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__47984\,
            in1 => \_gnd_net_\,
            in2 => \N__38522\,
            in3 => \N__38501\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47681\,
            ce => \N__47220\,
            sr => \N__46790\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__42546\,
            in1 => \N__41501\,
            in2 => \N__38459\,
            in3 => \N__41447\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42510\,
            in1 => \N__42547\,
            in2 => \_gnd_net_\,
            in3 => \N__48087\,
            lcout => \elapsed_time_ns_1_RNI2COBB_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48089\,
            in1 => \N__38865\,
            in2 => \_gnd_net_\,
            in3 => \N__38910\,
            lcout => \elapsed_time_ns_1_RNIU8PBB_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_30_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__39165\,
            in1 => \N__38846\,
            in2 => \N__39527\,
            in3 => \N__38825\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_df30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48088\,
            in1 => \N__38758\,
            in2 => \_gnd_net_\,
            in3 => \N__38796\,
            lcout => \elapsed_time_ns_1_RNIJI91B_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__38699\,
            in1 => \N__38737\,
            in2 => \_gnd_net_\,
            in3 => \N__48090\,
            lcout => \elapsed_time_ns_1_RNIV8OBB_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42002\,
            in2 => \N__38681\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_10_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47113\,
            in1 => \N__38648\,
            in2 => \_gnd_net_\,
            in3 => \N__38636\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \N__47660\,
            ce => 'H',
            sr => \N__46801\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__47117\,
            in1 => \N__38633\,
            in2 => \N__42158\,
            in3 => \N__38621\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \N__47660\,
            ce => 'H',
            sr => \N__46801\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47114\,
            in1 => \N__38618\,
            in2 => \_gnd_net_\,
            in3 => \N__38606\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \N__47660\,
            ce => 'H',
            sr => \N__46801\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47118\,
            in1 => \N__39032\,
            in2 => \_gnd_net_\,
            in3 => \N__39020\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \N__47660\,
            ce => 'H',
            sr => \N__46801\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47115\,
            in1 => \N__39017\,
            in2 => \_gnd_net_\,
            in3 => \N__39005\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \N__47660\,
            ce => 'H',
            sr => \N__46801\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47119\,
            in1 => \N__39002\,
            in2 => \_gnd_net_\,
            in3 => \N__38990\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \N__47660\,
            ce => 'H',
            sr => \N__46801\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47116\,
            in1 => \N__38987\,
            in2 => \_gnd_net_\,
            in3 => \N__38975\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \N__47660\,
            ce => 'H',
            sr => \N__46801\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47157\,
            in1 => \N__38972\,
            in2 => \_gnd_net_\,
            in3 => \N__38960\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_17_11_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \N__47650\,
            ce => 'H',
            sr => \N__46809\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47150\,
            in1 => \N__38957\,
            in2 => \_gnd_net_\,
            in3 => \N__38945\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \N__47650\,
            ce => 'H',
            sr => \N__46809\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47154\,
            in1 => \N__38942\,
            in2 => \_gnd_net_\,
            in3 => \N__38930\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \N__47650\,
            ce => 'H',
            sr => \N__46809\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47151\,
            in1 => \N__38927\,
            in2 => \_gnd_net_\,
            in3 => \N__38915\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \N__47650\,
            ce => 'H',
            sr => \N__46809\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47155\,
            in1 => \N__39134\,
            in2 => \_gnd_net_\,
            in3 => \N__39122\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \N__47650\,
            ce => 'H',
            sr => \N__46809\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47152\,
            in1 => \N__39119\,
            in2 => \_gnd_net_\,
            in3 => \N__39107\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \N__47650\,
            ce => 'H',
            sr => \N__46809\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47156\,
            in1 => \N__39104\,
            in2 => \_gnd_net_\,
            in3 => \N__39092\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \N__47650\,
            ce => 'H',
            sr => \N__46809\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47153\,
            in1 => \N__41587\,
            in2 => \_gnd_net_\,
            in3 => \N__39089\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \N__47650\,
            ce => 'H',
            sr => \N__46809\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47158\,
            in1 => \N__41568\,
            in2 => \_gnd_net_\,
            in3 => \N__39086\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_17_12_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \N__47637\,
            ce => 'H',
            sr => \N__46818\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47162\,
            in1 => \N__41968\,
            in2 => \_gnd_net_\,
            in3 => \N__39083\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \N__47637\,
            ce => 'H',
            sr => \N__46818\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47159\,
            in1 => \N__41984\,
            in2 => \_gnd_net_\,
            in3 => \N__39080\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \N__47637\,
            ce => 'H',
            sr => \N__46818\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47163\,
            in1 => \N__39072\,
            in2 => \_gnd_net_\,
            in3 => \N__39056\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \N__47637\,
            ce => 'H',
            sr => \N__46818\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47160\,
            in1 => \N__39051\,
            in2 => \_gnd_net_\,
            in3 => \N__39035\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\,
            clk => \N__47637\,
            ce => 'H',
            sr => \N__46818\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47164\,
            in1 => \N__39234\,
            in2 => \_gnd_net_\,
            in3 => \N__39215\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\,
            clk => \N__47637\,
            ce => 'H',
            sr => \N__46818\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47161\,
            in1 => \N__39207\,
            in2 => \_gnd_net_\,
            in3 => \N__39191\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\,
            clk => \N__47637\,
            ce => 'H',
            sr => \N__46818\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47165\,
            in1 => \N__46402\,
            in2 => \_gnd_net_\,
            in3 => \N__39188\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\,
            clk => \N__47637\,
            ce => 'H',
            sr => \N__46818\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47067\,
            in1 => \N__46434\,
            in2 => \_gnd_net_\,
            in3 => \N__39185\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_17_13_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\,
            clk => \N__47627\,
            ce => 'H',
            sr => \N__46828\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47188\,
            in1 => \N__46365\,
            in2 => \_gnd_net_\,
            in3 => \N__39182\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\,
            clk => \N__47627\,
            ce => 'H',
            sr => \N__46828\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47068\,
            in1 => \N__46329\,
            in2 => \_gnd_net_\,
            in3 => \N__39179\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\,
            clk => \N__47627\,
            ce => 'H',
            sr => \N__46828\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47189\,
            in1 => \N__45615\,
            in2 => \_gnd_net_\,
            in3 => \N__39176\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\,
            clk => \N__47627\,
            ce => 'H',
            sr => \N__46828\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47069\,
            in1 => \N__45594\,
            in2 => \_gnd_net_\,
            in3 => \N__39173\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\,
            clk => \N__47627\,
            ce => 'H',
            sr => \N__46828\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47190\,
            in1 => \N__39159\,
            in2 => \_gnd_net_\,
            in3 => \N__39137\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\,
            clk => \N__47627\,
            ce => 'H',
            sr => \N__46828\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47070\,
            in1 => \N__39516\,
            in2 => \_gnd_net_\,
            in3 => \N__39530\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47627\,
            ce => 'H',
            sr => \N__46828\
        );

    \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__42313\,
            in1 => \N__39494\,
            in2 => \_gnd_net_\,
            in3 => \N__42702\,
            lcout => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__42317\,
            in1 => \N__39452\,
            in2 => \_gnd_net_\,
            in3 => \N__42747\,
            lcout => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__42312\,
            in1 => \N__39405\,
            in2 => \_gnd_net_\,
            in3 => \N__42876\,
            lcout => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__42316\,
            in1 => \N__39369\,
            in2 => \_gnd_net_\,
            in3 => \N__42792\,
            lcout => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__42310\,
            in1 => \N__39321\,
            in2 => \_gnd_net_\,
            in3 => \N__42217\,
            lcout => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__42315\,
            in1 => \N__43685\,
            in2 => \_gnd_net_\,
            in3 => \N__43644\,
            lcout => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__42311\,
            in1 => \N__39280\,
            in2 => \_gnd_net_\,
            in3 => \N__42177\,
            lcout => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__42314\,
            in1 => \N__39822\,
            in2 => \_gnd_net_\,
            in3 => \N__42838\,
            lcout => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__44062\,
            in1 => \N__42362\,
            in2 => \_gnd_net_\,
            in3 => \N__43101\,
            lcout => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__43680\,
            in1 => \N__44418\,
            in2 => \N__45038\,
            in3 => \N__43645\,
            lcout => \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__39750\,
            in1 => \N__42361\,
            in2 => \_gnd_net_\,
            in3 => \N__43140\,
            lcout => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__42360\,
            in1 => \N__39702\,
            in2 => \_gnd_net_\,
            in3 => \N__43177\,
            lcout => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43679\,
            lcout => \current_shift_inst.un4_control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__42358\,
            in1 => \N__39660\,
            in2 => \_gnd_net_\,
            in3 => \N__42660\,
            lcout => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__39615\,
            in1 => \N__42359\,
            in2 => \_gnd_net_\,
            in3 => \N__42621\,
            lcout => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__42363\,
            in1 => \N__39572\,
            in2 => \_gnd_net_\,
            in3 => \N__43062\,
            lcout => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__40113\,
            in1 => \N__42364\,
            in2 => \_gnd_net_\,
            in3 => \N__43017\,
            lcout => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44426\,
            in1 => \N__40073\,
            in2 => \_gnd_net_\,
            in3 => \N__43290\,
            lcout => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__40017\,
            in1 => \N__42369\,
            in2 => \_gnd_net_\,
            in3 => \N__43423\,
            lcout => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__42365\,
            in1 => \_gnd_net_\,
            in2 => \N__42994\,
            in3 => \N__43959\,
            lcout => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__43392\,
            in1 => \N__39969\,
            in2 => \_gnd_net_\,
            in3 => \N__42370\,
            lcout => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__42368\,
            in1 => \N__42462\,
            in2 => \_gnd_net_\,
            in3 => \N__43473\,
            lcout => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__39918\,
            in1 => \N__42366\,
            in2 => \_gnd_net_\,
            in3 => \N__42948\,
            lcout => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__42367\,
            in1 => \N__39877\,
            in2 => \_gnd_net_\,
            in3 => \N__43506\,
            lcout => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__44007\,
            in1 => \N__44424\,
            in2 => \_gnd_net_\,
            in3 => \N__43716\,
            lcout => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__42382\,
            in1 => \N__40347\,
            in2 => \_gnd_net_\,
            in3 => \N__43341\,
            lcout => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44427\,
            in1 => \N__40302\,
            in2 => \_gnd_net_\,
            in3 => \N__43210\,
            lcout => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44423\,
            in1 => \N__40261\,
            in2 => \_gnd_net_\,
            in3 => \N__43743\,
            lcout => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__40262\,
            in1 => \N__44425\,
            in2 => \N__43750\,
            in3 => \N__44961\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44421\,
            in1 => \N__42466\,
            in2 => \N__45039\,
            in3 => \N__43474\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__44965\,
            in1 => \N__44420\,
            in2 => \N__43966\,
            in3 => \N__42993\,
            lcout => \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44422\,
            in1 => \N__40193\,
            in2 => \_gnd_net_\,
            in3 => \N__43248\,
            lcout => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.counter_0_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41325\,
            in1 => \N__40146\,
            in2 => \_gnd_net_\,
            in3 => \N__40127\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_17_18_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_0\,
            clk => \N__47582\,
            ce => \N__41197\,
            sr => \N__46858\
        );

    \current_shift_inst.timer_s1.counter_1_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41351\,
            in1 => \N__43593\,
            in2 => \_gnd_net_\,
            in3 => \N__40124\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_0\,
            carryout => \current_shift_inst.timer_s1.counter_cry_1\,
            clk => \N__47582\,
            ce => \N__41197\,
            sr => \N__46858\
        );

    \current_shift_inst.timer_s1.counter_2_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41326\,
            in1 => \N__40566\,
            in2 => \_gnd_net_\,
            in3 => \N__40550\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_1\,
            carryout => \current_shift_inst.timer_s1.counter_cry_2\,
            clk => \N__47582\,
            ce => \N__41197\,
            sr => \N__46858\
        );

    \current_shift_inst.timer_s1.counter_3_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41352\,
            in1 => \N__40536\,
            in2 => \_gnd_net_\,
            in3 => \N__40520\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_2\,
            carryout => \current_shift_inst.timer_s1.counter_cry_3\,
            clk => \N__47582\,
            ce => \N__41197\,
            sr => \N__46858\
        );

    \current_shift_inst.timer_s1.counter_4_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41327\,
            in1 => \N__40509\,
            in2 => \_gnd_net_\,
            in3 => \N__40493\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_3\,
            carryout => \current_shift_inst.timer_s1.counter_cry_4\,
            clk => \N__47582\,
            ce => \N__41197\,
            sr => \N__46858\
        );

    \current_shift_inst.timer_s1.counter_5_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41353\,
            in1 => \N__40482\,
            in2 => \_gnd_net_\,
            in3 => \N__40466\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_4\,
            carryout => \current_shift_inst.timer_s1.counter_cry_5\,
            clk => \N__47582\,
            ce => \N__41197\,
            sr => \N__46858\
        );

    \current_shift_inst.timer_s1.counter_6_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41328\,
            in1 => \N__40461\,
            in2 => \_gnd_net_\,
            in3 => \N__40445\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_5\,
            carryout => \current_shift_inst.timer_s1.counter_cry_6\,
            clk => \N__47582\,
            ce => \N__41197\,
            sr => \N__46858\
        );

    \current_shift_inst.timer_s1.counter_7_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41354\,
            in1 => \N__40440\,
            in2 => \_gnd_net_\,
            in3 => \N__40424\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_6\,
            carryout => \current_shift_inst.timer_s1.counter_cry_7\,
            clk => \N__47582\,
            ce => \N__41197\,
            sr => \N__46858\
        );

    \current_shift_inst.timer_s1.counter_8_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41344\,
            in1 => \N__40413\,
            in2 => \_gnd_net_\,
            in3 => \N__40391\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_17_19_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_8\,
            clk => \N__47578\,
            ce => \N__41198\,
            sr => \N__46863\
        );

    \current_shift_inst.timer_s1.counter_9_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41340\,
            in1 => \N__40374\,
            in2 => \_gnd_net_\,
            in3 => \N__40355\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_8\,
            carryout => \current_shift_inst.timer_s1.counter_cry_9\,
            clk => \N__47578\,
            ce => \N__41198\,
            sr => \N__46863\
        );

    \current_shift_inst.timer_s1.counter_10_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41341\,
            in1 => \N__40782\,
            in2 => \_gnd_net_\,
            in3 => \N__40766\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_9\,
            carryout => \current_shift_inst.timer_s1.counter_cry_10\,
            clk => \N__47578\,
            ce => \N__41198\,
            sr => \N__46863\
        );

    \current_shift_inst.timer_s1.counter_11_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41337\,
            in1 => \N__40761\,
            in2 => \_gnd_net_\,
            in3 => \N__40745\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_10\,
            carryout => \current_shift_inst.timer_s1.counter_cry_11\,
            clk => \N__47578\,
            ce => \N__41198\,
            sr => \N__46863\
        );

    \current_shift_inst.timer_s1.counter_12_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41342\,
            in1 => \N__40737\,
            in2 => \_gnd_net_\,
            in3 => \N__40718\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_11\,
            carryout => \current_shift_inst.timer_s1.counter_cry_12\,
            clk => \N__47578\,
            ce => \N__41198\,
            sr => \N__46863\
        );

    \current_shift_inst.timer_s1.counter_13_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41338\,
            in1 => \N__40710\,
            in2 => \_gnd_net_\,
            in3 => \N__40691\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_12\,
            carryout => \current_shift_inst.timer_s1.counter_cry_13\,
            clk => \N__47578\,
            ce => \N__41198\,
            sr => \N__46863\
        );

    \current_shift_inst.timer_s1.counter_14_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41343\,
            in1 => \N__40680\,
            in2 => \_gnd_net_\,
            in3 => \N__40664\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_13\,
            carryout => \current_shift_inst.timer_s1.counter_cry_14\,
            clk => \N__47578\,
            ce => \N__41198\,
            sr => \N__46863\
        );

    \current_shift_inst.timer_s1.counter_15_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41339\,
            in1 => \N__40653\,
            in2 => \_gnd_net_\,
            in3 => \N__40637\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_14\,
            carryout => \current_shift_inst.timer_s1.counter_cry_15\,
            clk => \N__47578\,
            ce => \N__41198\,
            sr => \N__46863\
        );

    \current_shift_inst.timer_s1.counter_16_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41347\,
            in1 => \N__40626\,
            in2 => \_gnd_net_\,
            in3 => \N__40604\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_17_20_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_16\,
            clk => \N__47573\,
            ce => \N__41193\,
            sr => \N__46868\
        );

    \current_shift_inst.timer_s1.counter_17_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41333\,
            in1 => \N__40587\,
            in2 => \_gnd_net_\,
            in3 => \N__40571\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_16\,
            carryout => \current_shift_inst.timer_s1.counter_cry_17\,
            clk => \N__47573\,
            ce => \N__41193\,
            sr => \N__46868\
        );

    \current_shift_inst.timer_s1.counter_18_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41348\,
            in1 => \N__41016\,
            in2 => \_gnd_net_\,
            in3 => \N__41000\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_17\,
            carryout => \current_shift_inst.timer_s1.counter_cry_18\,
            clk => \N__47573\,
            ce => \N__41193\,
            sr => \N__46868\
        );

    \current_shift_inst.timer_s1.counter_19_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41334\,
            in1 => \N__40992\,
            in2 => \_gnd_net_\,
            in3 => \N__40973\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_18\,
            carryout => \current_shift_inst.timer_s1.counter_cry_19\,
            clk => \N__47573\,
            ce => \N__41193\,
            sr => \N__46868\
        );

    \current_shift_inst.timer_s1.counter_20_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41349\,
            in1 => \N__40962\,
            in2 => \_gnd_net_\,
            in3 => \N__40946\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_19\,
            carryout => \current_shift_inst.timer_s1.counter_cry_20\,
            clk => \N__47573\,
            ce => \N__41193\,
            sr => \N__46868\
        );

    \current_shift_inst.timer_s1.counter_21_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41335\,
            in1 => \N__40941\,
            in2 => \_gnd_net_\,
            in3 => \N__40925\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_20\,
            carryout => \current_shift_inst.timer_s1.counter_cry_21\,
            clk => \N__47573\,
            ce => \N__41193\,
            sr => \N__46868\
        );

    \current_shift_inst.timer_s1.counter_22_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41350\,
            in1 => \N__40920\,
            in2 => \_gnd_net_\,
            in3 => \N__40904\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_21\,
            carryout => \current_shift_inst.timer_s1.counter_cry_22\,
            clk => \N__47573\,
            ce => \N__41193\,
            sr => \N__46868\
        );

    \current_shift_inst.timer_s1.counter_23_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41336\,
            in1 => \N__40893\,
            in2 => \_gnd_net_\,
            in3 => \N__40877\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_22\,
            carryout => \current_shift_inst.timer_s1.counter_cry_23\,
            clk => \N__47573\,
            ce => \N__41193\,
            sr => \N__46868\
        );

    \current_shift_inst.timer_s1.counter_24_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41329\,
            in1 => \N__40863\,
            in2 => \_gnd_net_\,
            in3 => \N__40841\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_17_21_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_24\,
            clk => \N__47568\,
            ce => \N__41186\,
            sr => \N__46872\
        );

    \current_shift_inst.timer_s1.counter_25_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41345\,
            in1 => \N__40830\,
            in2 => \_gnd_net_\,
            in3 => \N__40808\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_24\,
            carryout => \current_shift_inst.timer_s1.counter_cry_25\,
            clk => \N__47568\,
            ce => \N__41186\,
            sr => \N__46872\
        );

    \current_shift_inst.timer_s1.counter_26_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41330\,
            in1 => \N__40803\,
            in2 => \_gnd_net_\,
            in3 => \N__40787\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_25\,
            carryout => \current_shift_inst.timer_s1.counter_cry_26\,
            clk => \N__47568\,
            ce => \N__41186\,
            sr => \N__46872\
        );

    \current_shift_inst.timer_s1.counter_27_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41346\,
            in1 => \N__41394\,
            in2 => \_gnd_net_\,
            in3 => \N__41378\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_26\,
            carryout => \current_shift_inst.timer_s1.counter_cry_27\,
            clk => \N__47568\,
            ce => \N__41186\,
            sr => \N__46872\
        );

    \current_shift_inst.timer_s1.counter_28_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41331\,
            in1 => \N__41371\,
            in2 => \_gnd_net_\,
            in3 => \N__41357\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_27\,
            carryout => \current_shift_inst.timer_s1.counter_cry_28\,
            clk => \N__47568\,
            ce => \N__41186\,
            sr => \N__46872\
        );

    \current_shift_inst.timer_s1.counter_29_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__41212\,
            in1 => \N__41332\,
            in2 => \_gnd_net_\,
            in3 => \N__41219\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47568\,
            ce => \N__41186\,
            sr => \N__46872\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_18_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41672\,
            in1 => \N__41150\,
            in2 => \N__45840\,
            in3 => \N__41112\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_18_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41764\,
            in1 => \N__41739\,
            in2 => \_gnd_net_\,
            in3 => \N__47980\,
            lcout => \elapsed_time_ns_1_RNI4EOBB_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_18_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__45926\,
            in1 => \N__45757\,
            in2 => \N__47777\,
            in3 => \N__41062\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_18_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41833\,
            in1 => \N__41808\,
            in2 => \_gnd_net_\,
            in3 => \N__47981\,
            lcout => \elapsed_time_ns_1_RNILK91B_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_16_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41459\,
            in1 => \N__41416\,
            in2 => \_gnd_net_\,
            in3 => \N__48001\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47692\,
            ce => \N__47204\,
            sr => \N__46787\
        );

    \phase_controller_inst1.stoper_tr.target_time_9_LC_18_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48000\,
            in1 => \N__41829\,
            in2 => \_gnd_net_\,
            in3 => \N__41813\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47692\,
            ce => \N__47204\,
            sr => \N__46787\
        );

    \phase_controller_inst1.stoper_tr.target_time_17_LC_18_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__41754\,
            in1 => \_gnd_net_\,
            in2 => \N__41740\,
            in3 => \N__48002\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47692\,
            ce => \N__47204\,
            sr => \N__46787\
        );

    \phase_controller_inst1.stoper_tr.target_time_23_LC_18_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47999\,
            in1 => \N__41691\,
            in2 => \_gnd_net_\,
            in3 => \N__41675\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47692\,
            ce => \N__47204\,
            sr => \N__46787\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__41593\,
            in1 => \N__41603\,
            in2 => \N__41552\,
            in3 => \N__41572\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__41602\,
            in1 => \N__41594\,
            in2 => \N__41573\,
            in3 => \N__41551\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_14_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41528\,
            in1 => \N__41502\,
            in2 => \_gnd_net_\,
            in3 => \N__48051\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47682\,
            ce => \N__47202\,
            sr => \N__46791\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41415\,
            in1 => \N__41455\,
            in2 => \_gnd_net_\,
            in3 => \N__48026\,
            lcout => \elapsed_time_ns_1_RNI3DOBB_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48025\,
            in1 => \N__41925\,
            in2 => \_gnd_net_\,
            in3 => \N__41905\,
            lcout => \elapsed_time_ns_1_RNI6GOBB_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__45497\,
            in1 => \N__42121\,
            in2 => \_gnd_net_\,
            in3 => \N__45556\,
            lcout => \phase_controller_inst1.stoper_tr.un2_start_0\,
            ltout => \phase_controller_inst1.stoper_tr.un2_start_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4_28_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42161\,
            in3 => \N__42058\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.running_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111001100"
        )
    port map (
            in0 => \N__45499\,
            in1 => \N__42122\,
            in2 => \N__42149\,
            in3 => \N__42021\,
            lcout => \phase_controller_inst1.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47661\,
            ce => 'H',
            sr => \N__46802\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIIMJC3_28_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100111011"
        )
    port map (
            in0 => \N__42109\,
            in1 => \N__45498\,
            in2 => \N__42086\,
            in3 => \N__42074\,
            lcout => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42047\,
            in3 => \N__42020\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__41982\,
            in1 => \N__41964\,
            in2 => \N__41867\,
            in3 => \N__42560\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__42559\,
            in1 => \N__41983\,
            in2 => \N__41969\,
            in3 => \N__41863\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_19_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__48131\,
            in1 => \_gnd_net_\,
            in2 => \N__41935\,
            in3 => \N__41900\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47651\,
            ce => \N__47172\,
            sr => \N__46810\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42597\,
            in1 => \N__41845\,
            in2 => \_gnd_net_\,
            in3 => \N__48129\,
            lcout => \elapsed_time_ns_1_RNI5FOBB_0_18\,
            ltout => \elapsed_time_ns_1_RNI5FOBB_0_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_18_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__48130\,
            in1 => \_gnd_net_\,
            in2 => \N__42602\,
            in3 => \N__42598\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47651\,
            ce => \N__47172\,
            sr => \N__46810\
        );

    \phase_controller_inst1.stoper_tr.target_time_15_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42551\,
            in1 => \N__42517\,
            in2 => \_gnd_net_\,
            in3 => \N__48132\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47651\,
            ce => \N__47172\,
            sr => \N__46810\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__44415\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44954\,
            lcout => \current_shift_inst.un38_control_input_axb_31_s0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__42467\,
            in1 => \N__44414\,
            in2 => \N__45037\,
            in3 => \N__43478\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42414\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47638\,
            ce => \N__43574\,
            sr => \N__46819\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43544\,
            in2 => \N__42266\,
            in3 => \N__42265\,
            lcout => \current_shift_inst.un4_control_input1_2\,
            ltout => OPEN,
            carryin => \bfn_18_14_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42242\,
            in2 => \_gnd_net_\,
            in3 => \N__42206\,
            lcout => \current_shift_inst.un4_control_input1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_1\,
            carryout => \current_shift_inst.un4_control_input_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42203\,
            in2 => \_gnd_net_\,
            in3 => \N__42164\,
            lcout => \current_shift_inst.un4_control_input1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_2\,
            carryout => \current_shift_inst.un4_control_input_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42902\,
            in2 => \_gnd_net_\,
            in3 => \N__42863\,
            lcout => \current_shift_inst.un4_control_input1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_3\,
            carryout => \current_shift_inst.un4_control_input_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42860\,
            in2 => \_gnd_net_\,
            in3 => \N__42827\,
            lcout => \current_shift_inst.un4_control_input1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_4\,
            carryout => \current_shift_inst.un4_control_input_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42824\,
            in2 => \_gnd_net_\,
            in3 => \N__42818\,
            lcout => \current_shift_inst.un4_control_input1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_5\,
            carryout => \current_shift_inst.un4_control_input_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42815\,
            in2 => \_gnd_net_\,
            in3 => \N__42776\,
            lcout => \current_shift_inst.un4_control_input1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_6\,
            carryout => \current_shift_inst.un4_control_input_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42773\,
            in2 => \_gnd_net_\,
            in3 => \N__42734\,
            lcout => \current_shift_inst.un4_control_input1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_7\,
            carryout => \current_shift_inst.un4_control_input_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42731\,
            in2 => \_gnd_net_\,
            in3 => \N__42689\,
            lcout => \current_shift_inst.un4_control_input1_10\,
            ltout => OPEN,
            carryin => \bfn_18_15_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42686\,
            in2 => \_gnd_net_\,
            in3 => \N__42647\,
            lcout => \current_shift_inst.un4_control_input1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_9\,
            carryout => \current_shift_inst.un4_control_input_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42644\,
            in2 => \_gnd_net_\,
            in3 => \N__42605\,
            lcout => \current_shift_inst.un4_control_input1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_10\,
            carryout => \current_shift_inst.un4_control_input_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43196\,
            in2 => \_gnd_net_\,
            in3 => \N__43166\,
            lcout => \current_shift_inst.un4_control_input1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_11\,
            carryout => \current_shift_inst.un4_control_input_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43163\,
            in2 => \_gnd_net_\,
            in3 => \N__43124\,
            lcout => \current_shift_inst.un4_control_input1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_12\,
            carryout => \current_shift_inst.un4_control_input_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44024\,
            in2 => \_gnd_net_\,
            in3 => \N__43085\,
            lcout => \current_shift_inst.un4_control_input1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_13\,
            carryout => \current_shift_inst.un4_control_input_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43082\,
            in2 => \_gnd_net_\,
            in3 => \N__43046\,
            lcout => \current_shift_inst.un4_control_input1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_14\,
            carryout => \current_shift_inst.un4_control_input_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43043\,
            in2 => \_gnd_net_\,
            in3 => \N__43001\,
            lcout => \current_shift_inst.un4_control_input1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_15\,
            carryout => \current_shift_inst.un4_control_input_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43916\,
            in2 => \_gnd_net_\,
            in3 => \N__42971\,
            lcout => \current_shift_inst.un4_control_input1_18\,
            ltout => OPEN,
            carryin => \bfn_18_16_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42968\,
            in2 => \_gnd_net_\,
            in3 => \N__42935\,
            lcout => \current_shift_inst.un4_control_input1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_17\,
            carryout => \current_shift_inst.un4_control_input_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43871\,
            in2 => \_gnd_net_\,
            in3 => \N__42905\,
            lcout => \current_shift_inst.un4_control_input1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_18\,
            carryout => \current_shift_inst.un4_control_input_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43532\,
            in2 => \_gnd_net_\,
            in3 => \N__43493\,
            lcout => \current_shift_inst.un4_control_input1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_19\,
            carryout => \current_shift_inst.un4_control_input_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43490\,
            in2 => \_gnd_net_\,
            in3 => \N__43457\,
            lcout => \current_shift_inst.un4_control_input1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_20\,
            carryout => \current_shift_inst.un4_control_input_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43454\,
            in2 => \_gnd_net_\,
            in3 => \N__43412\,
            lcout => \current_shift_inst.un4_control_input1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_21\,
            carryout => \current_shift_inst.un4_control_input_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43409\,
            in2 => \_gnd_net_\,
            in3 => \N__43370\,
            lcout => \current_shift_inst.un4_control_input1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_22\,
            carryout => \current_shift_inst.un4_control_input_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_18_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43367\,
            in2 => \_gnd_net_\,
            in3 => \N__43325\,
            lcout => \current_shift_inst.un4_control_input1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_23\,
            carryout => \current_shift_inst.un4_control_input_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43322\,
            in2 => \_gnd_net_\,
            in3 => \N__43277\,
            lcout => \current_shift_inst.un4_control_input1_26\,
            ltout => OPEN,
            carryin => \bfn_18_17_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43274\,
            in2 => \_gnd_net_\,
            in3 => \N__43232\,
            lcout => \current_shift_inst.un4_control_input1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_25\,
            carryout => \current_shift_inst.un4_control_input_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43229\,
            in2 => \_gnd_net_\,
            in3 => \N__43199\,
            lcout => \current_shift_inst.un4_control_input1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_26\,
            carryout => \current_shift_inst.un4_control_input_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43766\,
            in2 => \_gnd_net_\,
            in3 => \N__43730\,
            lcout => \current_shift_inst.un4_control_input1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_27\,
            carryout => \current_shift_inst.un4_control_input_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43976\,
            in2 => \_gnd_net_\,
            in3 => \N__43703\,
            lcout => \current_shift_inst.un4_control_input1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_28\,
            carryout => \current_shift_inst.un4_control_input1_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43700\,
            lcout => \current_shift_inst.un4_control_input1_31_THRU_CO\,
            ltout => \current_shift_inst.un4_control_input1_31_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43697\,
            in3 => \N__44397\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44396\,
            in1 => \N__43684\,
            in2 => \N__45055\,
            in3 => \N__43649\,
            lcout => \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__44393\,
            in1 => \N__45218\,
            in2 => \N__45167\,
            in3 => \N__45186\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43594\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47588\,
            ce => \N__43573\,
            sr => \N__46852\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45182\,
            lcout => \current_shift_inst.un4_control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__45217\,
            in1 => \N__44392\,
            in2 => \N__45190\,
            in3 => \N__45166\,
            lcout => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__44394\,
            in1 => \N__45050\,
            in2 => \N__45092\,
            in3 => \N__45100\,
            lcout => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__45101\,
            in1 => \N__45088\,
            in2 => \N__45056\,
            in3 => \N__44395\,
            lcout => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44046\,
            lcout => \current_shift_inst.un4_control_input_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43997\,
            lcout => \current_shift_inst.un4_control_input_1_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43949\,
            lcout => \current_shift_inst.un4_control_input_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43890\,
            lcout => \current_shift_inst.un4_control_input_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_10_LC_18_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43862\,
            lcout => \N_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47566\,
            ce => 'H',
            sr => \N__46877\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_20_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001100"
        )
    port map (
            in0 => \N__45418\,
            in1 => \N__45971\,
            in2 => \N__45449\,
            in3 => \N__45992\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_20_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__45991\,
            in1 => \N__45448\,
            in2 => \N__45422\,
            in3 => \N__45970\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_20_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__45310\,
            in1 => \N__45371\,
            in2 => \N__45347\,
            in3 => \N__45979\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_20_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__45370\,
            in1 => \N__45311\,
            in2 => \N__45983\,
            in3 => \N__45346\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_20_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45705\,
            in1 => \N__45667\,
            in2 => \_gnd_net_\,
            in3 => \N__48152\,
            lcout => \elapsed_time_ns_1_RNI6HPBB_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_26_LC_20_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45787\,
            in1 => \N__45770\,
            in2 => \_gnd_net_\,
            in3 => \N__48178\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47693\,
            ce => \N__45958\,
            sr => \N__46795\
        );

    \phase_controller_inst2.stoper_tr.target_time_29_LC_20_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48177\,
            in1 => \N__45884\,
            in2 => \_gnd_net_\,
            in3 => \N__45928\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47693\,
            ce => \N__45958\,
            sr => \N__46795\
        );

    \phase_controller_inst2.stoper_tr.target_time_28_LC_20_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48176\,
            in1 => \N__45713\,
            in2 => \_gnd_net_\,
            in3 => \N__45663\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47693\,
            ce => \N__45958\,
            sr => \N__46795\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_20_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101110"
        )
    port map (
            in0 => \N__45227\,
            in1 => \N__45287\,
            in2 => \N__45256\,
            in3 => \N__45278\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_20_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__45286\,
            in1 => \N__45277\,
            in2 => \N__45257\,
            in3 => \N__45226\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_20_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__47722\,
            in1 => \N__48151\,
            in2 => \_gnd_net_\,
            in3 => \N__47775\,
            lcout => \elapsed_time_ns_1_RNI3EPBB_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_28_LC_20_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45712\,
            in1 => \N__45668\,
            in2 => \_gnd_net_\,
            in3 => \N__48199\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47674\,
            ce => \N__47237\,
            sr => \N__46811\
        );

    \phase_controller_inst1.stoper_tr.target_time_29_LC_20_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48198\,
            in1 => \N__45883\,
            in2 => \_gnd_net_\,
            in3 => \N__45929\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47674\,
            ce => \N__47237\,
            sr => \N__46811\
        );

    \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_20_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45488\,
            in2 => \_gnd_net_\,
            in3 => \N__45557\,
            lcout => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_20_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__45628\,
            in1 => \N__45619\,
            in2 => \N__45599\,
            in3 => \N__45637\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_20_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101110"
        )
    port map (
            in0 => \N__45638\,
            in1 => \N__45629\,
            in2 => \N__45620\,
            in3 => \N__45598\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_20_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__46346\,
            in1 => \N__46330\,
            in2 => \N__46370\,
            in3 => \N__46307\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.start_latched_LC_20_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45555\,
            lcout => \phase_controller_inst1.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47640\,
            ce => 'H',
            sr => \N__46834\
        );

    \phase_controller_inst2.stoper_tr.target_time_24_LC_21_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__45863\,
            in1 => \_gnd_net_\,
            in2 => \N__48204\,
            in3 => \N__45842\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47700\,
            ce => \N__45959\,
            sr => \N__46796\
        );

    \phase_controller_inst2.stoper_tr.target_time_27_LC_21_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__48286\,
            in1 => \N__48169\,
            in2 => \_gnd_net_\,
            in3 => \N__48222\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47700\,
            ce => \N__45959\,
            sr => \N__46796\
        );

    \phase_controller_inst2.stoper_tr.target_time_25_LC_21_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__47723\,
            in1 => \_gnd_net_\,
            in2 => \N__48205\,
            in3 => \N__47776\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47700\,
            ce => \N__45959\,
            sr => \N__46796\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_21_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__48285\,
            in1 => \N__48226\,
            in2 => \_gnd_net_\,
            in3 => \N__48153\,
            lcout => \elapsed_time_ns_1_RNI5GPBB_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_21_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48154\,
            in1 => \N__45882\,
            in2 => \_gnd_net_\,
            in3 => \N__45927\,
            lcout => \elapsed_time_ns_1_RNI7IPBB_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_21_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45862\,
            in1 => \N__45841\,
            in2 => \_gnd_net_\,
            in3 => \N__48149\,
            lcout => \elapsed_time_ns_1_RNI2DPBB_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_21_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48150\,
            in1 => \N__45788\,
            in2 => \_gnd_net_\,
            in3 => \N__45769\,
            lcout => \elapsed_time_ns_1_RNI4FPBB_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_24_LC_21_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45858\,
            in1 => \N__45830\,
            in2 => \_gnd_net_\,
            in3 => \N__48202\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47683\,
            ce => \N__47236\,
            sr => \N__46820\
        );

    \phase_controller_inst1.stoper_tr.target_time_26_LC_21_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48201\,
            in1 => \N__45786\,
            in2 => \_gnd_net_\,
            in3 => \N__45756\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47683\,
            ce => \N__47236\,
            sr => \N__46820\
        );

    \phase_controller_inst1.stoper_tr.target_time_27_LC_21_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__48287\,
            in1 => \N__48227\,
            in2 => \_gnd_net_\,
            in3 => \N__48203\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47683\,
            ce => \N__47236\,
            sr => \N__46820\
        );

    \phase_controller_inst1.stoper_tr.target_time_25_LC_21_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48200\,
            in1 => \N__47762\,
            in2 => \_gnd_net_\,
            in3 => \N__47718\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47683\,
            ce => \N__47236\,
            sr => \N__46820\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_21_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__46445\,
            in1 => \N__46435\,
            in2 => \N__46414\,
            in3 => \N__46388\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_21_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__46444\,
            in1 => \N__46436\,
            in2 => \N__46415\,
            in3 => \N__46387\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_21_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111100001101"
        )
    port map (
            in0 => \N__46366\,
            in1 => \N__46345\,
            in2 => \N__46334\,
            in3 => \N__46306\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_24_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__46270\,
            in1 => \N__46209\,
            in2 => \_gnd_net_\,
            in3 => \N__46079\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
